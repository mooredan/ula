magic
tech amic5n
timestamp 1624387645
<< nwell >>
rect -130 550 1930 1495
<< ntransistor >>
rect 175 115 235 400
rect 365 115 425 400
rect 555 115 615 400
rect 745 115 805 400
rect 935 115 995 400
rect 1125 115 1185 400
rect 1315 115 1375 400
rect 1505 115 1565 400
<< ptransistor >>
rect 175 705 235 1300
rect 365 705 425 1300
rect 555 705 615 1300
rect 745 705 805 1300
rect 935 705 995 1300
rect 1125 705 1185 1300
rect 1315 705 1375 1300
rect 1505 705 1565 1300
<< nselect >>
rect -10 0 1810 430
<< pselect >>
rect -10 670 1810 1440
<< ndiffusion >>
rect 55 370 175 400
rect 55 320 85 370
rect 135 320 175 370
rect 55 205 175 320
rect 55 155 85 205
rect 135 155 175 205
rect 55 115 175 155
rect 235 370 365 400
rect 235 320 275 370
rect 325 320 365 370
rect 235 205 365 320
rect 235 155 275 205
rect 325 155 365 205
rect 235 115 365 155
rect 425 345 555 400
rect 425 295 465 345
rect 515 295 555 345
rect 425 205 555 295
rect 425 155 465 205
rect 515 155 555 205
rect 425 115 555 155
rect 615 370 745 400
rect 615 320 655 370
rect 705 320 745 370
rect 615 205 745 320
rect 615 155 655 205
rect 705 155 745 205
rect 615 115 745 155
rect 805 345 935 400
rect 805 295 845 345
rect 895 295 935 345
rect 805 205 935 295
rect 805 155 845 205
rect 895 155 935 205
rect 805 115 935 155
rect 995 370 1125 400
rect 995 320 1035 370
rect 1085 320 1125 370
rect 995 205 1125 320
rect 995 155 1035 205
rect 1085 155 1125 205
rect 995 115 1125 155
rect 1185 355 1315 400
rect 1185 305 1225 355
rect 1275 305 1315 355
rect 1185 205 1315 305
rect 1185 155 1225 205
rect 1275 155 1315 205
rect 1185 115 1315 155
rect 1375 370 1505 400
rect 1375 320 1415 370
rect 1465 320 1505 370
rect 1375 205 1505 320
rect 1375 155 1415 205
rect 1465 155 1505 205
rect 1375 115 1505 155
rect 1565 345 1695 400
rect 1565 295 1605 345
rect 1655 295 1695 345
rect 1565 205 1695 295
rect 1565 155 1605 205
rect 1655 155 1695 205
rect 1565 115 1695 155
<< pdiffusion >>
rect 55 1260 175 1300
rect 55 1210 85 1260
rect 135 1210 175 1260
rect 55 1115 175 1210
rect 55 1065 85 1115
rect 135 1065 175 1115
rect 55 1015 175 1065
rect 55 965 85 1015
rect 135 965 175 1015
rect 55 915 175 965
rect 55 865 85 915
rect 135 865 175 915
rect 55 815 175 865
rect 55 765 85 815
rect 135 765 175 815
rect 55 705 175 765
rect 235 1260 365 1300
rect 235 1210 275 1260
rect 325 1210 365 1260
rect 235 1080 365 1210
rect 235 1030 275 1080
rect 325 1030 365 1080
rect 235 980 365 1030
rect 235 930 275 980
rect 325 930 365 980
rect 235 825 365 930
rect 235 775 275 825
rect 325 775 365 825
rect 235 705 365 775
rect 425 1260 555 1300
rect 425 1210 465 1260
rect 515 1210 555 1260
rect 425 1115 555 1210
rect 425 1065 465 1115
rect 515 1065 555 1115
rect 425 975 555 1065
rect 425 925 465 975
rect 515 925 555 975
rect 425 705 555 925
rect 615 1260 745 1300
rect 615 1210 655 1260
rect 705 1210 745 1260
rect 615 1080 745 1210
rect 615 1030 655 1080
rect 705 1030 745 1080
rect 615 980 745 1030
rect 615 930 655 980
rect 705 930 745 980
rect 615 825 745 930
rect 615 775 655 825
rect 705 775 745 825
rect 615 705 745 775
rect 805 1260 935 1300
rect 805 1210 845 1260
rect 895 1210 935 1260
rect 805 1115 935 1210
rect 805 1065 845 1115
rect 895 1065 935 1115
rect 805 975 935 1065
rect 805 925 845 975
rect 895 925 935 975
rect 805 705 935 925
rect 995 1260 1125 1300
rect 995 1210 1035 1260
rect 1085 1210 1125 1260
rect 995 1080 1125 1210
rect 995 1030 1035 1080
rect 1085 1030 1125 1080
rect 995 980 1125 1030
rect 995 930 1035 980
rect 1085 930 1125 980
rect 995 825 1125 930
rect 995 775 1035 825
rect 1085 775 1125 825
rect 995 705 1125 775
rect 1185 1260 1315 1300
rect 1185 1210 1225 1260
rect 1275 1210 1315 1260
rect 1185 1115 1315 1210
rect 1185 1065 1225 1115
rect 1275 1065 1315 1115
rect 1185 975 1315 1065
rect 1185 925 1225 975
rect 1275 925 1315 975
rect 1185 705 1315 925
rect 1375 1260 1505 1300
rect 1375 1210 1415 1260
rect 1465 1210 1505 1260
rect 1375 1080 1505 1210
rect 1375 1030 1415 1080
rect 1465 1030 1505 1080
rect 1375 980 1505 1030
rect 1375 930 1415 980
rect 1465 930 1505 980
rect 1375 825 1505 930
rect 1375 775 1415 825
rect 1465 775 1505 825
rect 1375 705 1505 775
rect 1565 1260 1695 1300
rect 1565 1210 1605 1260
rect 1655 1210 1695 1260
rect 1565 1115 1695 1210
rect 1565 1065 1605 1115
rect 1655 1065 1695 1115
rect 1565 975 1695 1065
rect 1565 925 1605 975
rect 1655 925 1695 975
rect 1565 705 1695 925
<< ndcontact >>
rect 85 320 135 370
rect 85 155 135 205
rect 275 320 325 370
rect 275 155 325 205
rect 465 295 515 345
rect 465 155 515 205
rect 655 320 705 370
rect 655 155 705 205
rect 845 295 895 345
rect 845 155 895 205
rect 1035 320 1085 370
rect 1035 155 1085 205
rect 1225 305 1275 355
rect 1225 155 1275 205
rect 1415 320 1465 370
rect 1415 155 1465 205
rect 1605 295 1655 345
rect 1605 155 1655 205
<< pdcontact >>
rect 85 1210 135 1260
rect 85 1065 135 1115
rect 85 965 135 1015
rect 85 865 135 915
rect 85 765 135 815
rect 275 1210 325 1260
rect 275 1030 325 1080
rect 275 930 325 980
rect 275 775 325 825
rect 465 1210 515 1260
rect 465 1065 515 1115
rect 465 925 515 975
rect 655 1210 705 1260
rect 655 1030 705 1080
rect 655 930 705 980
rect 655 775 705 825
rect 845 1210 895 1260
rect 845 1065 895 1115
rect 845 925 895 975
rect 1035 1210 1085 1260
rect 1035 1030 1085 1080
rect 1035 930 1085 980
rect 1035 775 1085 825
rect 1225 1210 1275 1260
rect 1225 1065 1275 1115
rect 1225 925 1275 975
rect 1415 1210 1465 1260
rect 1415 1030 1465 1080
rect 1415 930 1465 980
rect 1415 775 1465 825
rect 1605 1210 1655 1260
rect 1605 1065 1655 1115
rect 1605 925 1655 975
<< polysilicon >>
rect 175 1300 235 1365
rect 365 1300 425 1365
rect 555 1300 615 1365
rect 745 1300 805 1365
rect 935 1300 995 1365
rect 1125 1300 1185 1365
rect 1315 1300 1375 1365
rect 1505 1300 1565 1365
rect 175 685 235 705
rect 365 685 425 705
rect 555 685 615 705
rect 745 685 805 705
rect 935 685 995 705
rect 1125 685 1185 705
rect 1315 685 1375 705
rect 1505 685 1565 705
rect 65 665 1565 685
rect 65 615 85 665
rect 135 615 185 665
rect 235 615 285 665
rect 335 615 385 665
rect 435 615 485 665
rect 535 615 585 665
rect 635 615 685 665
rect 735 615 825 665
rect 875 615 925 665
rect 975 615 1025 665
rect 1075 615 1125 665
rect 1175 615 1225 665
rect 1275 615 1325 665
rect 1375 615 1425 665
rect 1475 615 1565 665
rect 65 595 1565 615
rect 175 400 235 595
rect 365 400 425 595
rect 555 400 615 595
rect 745 400 805 595
rect 935 400 995 595
rect 1125 400 1185 595
rect 1315 400 1375 595
rect 1505 400 1565 595
rect 175 50 235 115
rect 365 50 425 115
rect 555 50 615 115
rect 745 50 805 115
rect 935 50 995 115
rect 1125 50 1185 115
rect 1315 50 1375 115
rect 1505 50 1565 115
<< polycontact >>
rect 85 615 135 665
rect 185 615 235 665
rect 285 615 335 665
rect 385 615 435 665
rect 485 615 535 665
rect 585 615 635 665
rect 685 615 735 665
rect 825 615 875 665
rect 925 615 975 665
rect 1025 615 1075 665
rect 1125 615 1175 665
rect 1225 615 1275 665
rect 1325 615 1375 665
rect 1425 615 1475 665
<< metal1 >>
rect 0 1395 1800 1485
rect 65 1260 155 1395
rect 65 1210 85 1260
rect 135 1210 155 1260
rect 65 1115 155 1210
rect 65 1065 85 1115
rect 135 1065 155 1115
rect 65 1015 155 1065
rect 65 965 85 1015
rect 135 965 155 1015
rect 65 915 155 965
rect 65 865 85 915
rect 135 865 155 915
rect 65 815 155 865
rect 65 765 85 815
rect 135 765 155 815
rect 65 745 155 765
rect 255 1260 345 1290
rect 255 1210 275 1260
rect 325 1210 345 1260
rect 255 1080 345 1210
rect 255 1030 275 1080
rect 325 1030 345 1080
rect 255 980 345 1030
rect 255 930 275 980
rect 325 930 345 980
rect 255 845 345 930
rect 445 1260 535 1395
rect 445 1210 465 1260
rect 515 1210 535 1260
rect 445 1115 535 1210
rect 445 1065 465 1115
rect 515 1065 535 1115
rect 445 975 535 1065
rect 445 925 465 975
rect 515 925 535 975
rect 445 905 535 925
rect 635 1260 725 1290
rect 635 1210 655 1260
rect 705 1210 725 1260
rect 635 1080 725 1210
rect 635 1030 655 1080
rect 705 1030 725 1080
rect 635 980 725 1030
rect 635 930 655 980
rect 705 930 725 980
rect 635 845 725 930
rect 825 1260 915 1395
rect 825 1210 845 1260
rect 895 1210 915 1260
rect 825 1115 915 1210
rect 825 1065 845 1115
rect 895 1065 915 1115
rect 825 975 915 1065
rect 825 925 845 975
rect 895 925 915 975
rect 825 905 915 925
rect 1015 1260 1105 1290
rect 1015 1210 1035 1260
rect 1085 1210 1105 1260
rect 1015 1080 1105 1210
rect 1015 1030 1035 1080
rect 1085 1030 1105 1080
rect 1015 980 1105 1030
rect 1015 930 1035 980
rect 1085 930 1105 980
rect 1015 845 1105 930
rect 1205 1260 1295 1395
rect 1205 1210 1225 1260
rect 1275 1210 1295 1260
rect 1205 1115 1295 1210
rect 1205 1065 1225 1115
rect 1275 1065 1295 1115
rect 1205 975 1295 1065
rect 1205 925 1225 975
rect 1275 925 1295 975
rect 1205 905 1295 925
rect 1395 1260 1485 1290
rect 1395 1210 1415 1260
rect 1465 1210 1485 1260
rect 1395 1080 1485 1210
rect 1395 1030 1415 1080
rect 1465 1030 1485 1080
rect 1395 980 1485 1030
rect 1395 930 1415 980
rect 1465 930 1485 980
rect 1395 845 1485 930
rect 1585 1260 1675 1395
rect 1585 1210 1605 1260
rect 1655 1210 1675 1260
rect 1585 1115 1675 1210
rect 1585 1065 1605 1115
rect 1655 1065 1675 1115
rect 1585 975 1675 1065
rect 1585 925 1605 975
rect 1655 925 1675 975
rect 1585 905 1675 925
rect 255 825 1675 845
rect 255 775 275 825
rect 325 775 655 825
rect 705 775 1035 825
rect 1085 775 1415 825
rect 1465 775 1675 825
rect 255 755 1675 775
rect 65 665 1505 685
rect 65 615 85 665
rect 135 615 185 665
rect 235 615 285 665
rect 335 615 385 665
rect 435 615 485 665
rect 535 615 585 665
rect 635 615 685 665
rect 735 615 825 665
rect 875 615 925 665
rect 975 615 1025 665
rect 1075 615 1125 665
rect 1175 615 1225 665
rect 1275 615 1325 665
rect 1375 615 1425 665
rect 1475 615 1505 665
rect 65 595 1505 615
rect 1585 525 1675 755
rect 255 435 1675 525
rect 65 370 155 390
rect 65 320 85 370
rect 135 320 155 370
rect 65 205 155 320
rect 65 155 85 205
rect 135 155 155 205
rect 65 45 155 155
rect 255 370 345 435
rect 255 320 275 370
rect 325 320 345 370
rect 635 370 725 435
rect 255 205 345 320
rect 255 155 275 205
rect 325 155 345 205
rect 255 125 345 155
rect 445 345 535 365
rect 445 295 465 345
rect 515 295 535 345
rect 445 205 535 295
rect 445 155 465 205
rect 515 155 535 205
rect 445 45 535 155
rect 635 320 655 370
rect 705 320 725 370
rect 1015 370 1105 435
rect 635 205 725 320
rect 635 155 655 205
rect 705 155 725 205
rect 635 125 725 155
rect 825 345 915 365
rect 825 295 845 345
rect 895 295 915 345
rect 825 205 915 295
rect 825 155 845 205
rect 895 155 915 205
rect 825 45 915 155
rect 1015 320 1035 370
rect 1085 320 1105 370
rect 1015 205 1105 320
rect 1015 155 1035 205
rect 1085 155 1105 205
rect 1015 125 1105 155
rect 1205 355 1295 375
rect 1205 305 1225 355
rect 1275 305 1295 355
rect 1205 205 1295 305
rect 1205 155 1225 205
rect 1275 155 1295 205
rect 1205 45 1295 155
rect 1395 370 1485 435
rect 1395 320 1415 370
rect 1465 320 1485 370
rect 1395 205 1485 320
rect 1395 155 1415 205
rect 1465 155 1485 205
rect 1395 125 1485 155
rect 1585 345 1675 365
rect 1585 295 1605 345
rect 1655 295 1675 345
rect 1585 205 1675 295
rect 1585 155 1605 205
rect 1655 155 1675 205
rect 1585 45 1675 155
rect 0 -45 1800 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 3 ne
flabel metal1 s 20 1430 20 1430 2 FreeSans 400 0 0 0 vdd
port 2 ne
flabel metal1 s 285 470 285 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 85 605 85 605 2 FreeSans 400 0 0 0 a
port 1 ne
flabel nwell 50 555 50 555 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
