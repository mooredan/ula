`celldefine
module decap3 ();
endmodule
`endcelldefine
