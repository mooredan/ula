* Transient simulation of pad_x0_top and pad_in_top
*
* CMOS inverter for the crystal pad

.include pad_xtal.cir
.include mag/pad_in_top.cir
.include mag/pad_x0_top.cir
.include mag/schmitt.cir

.lib device_models/AMI_C5N.lib TT
.lib device_models/AMI_C5N_rmodels.lib NOM 

.param VDD_VAL=5
+      FREQ=6.5Meg
+      PER={1 / FREQ}
+      PH={PER / 2.0}
+      TRF={PER * 0.1}
+      VO=0
+      VA=0.100

.csparam tgt_freq={FREQ}


* power supply
Vvdd vdd 0 DC VDD_VAL
Vvss vss 0 DC 0

Vsrc src 0 DC 0 AC {VA}
Rsrc src 0 50

Cin src srcx 1.0e-6
vin srcx xin DC 0

xdut xout xin ckout vdd vss pad_xtal

Cckout ckout 0 0.1e-12

Rf xout xin 2.2Meg

RL xout 0 1.0k
CL xout 0 30.0e-12

.save all

.ac lin 20001 0.01Meg 20.01Meg

.control
destroy all
run

setplot ac1 
* plot mag(v(a)) mag(v(pad))

let gaindb = 20 * log10(mag(v(xout))/mag(v(xin)))
let f = re(frequency)
let v_xin = v(xin)
let i_xin = i(vin)
let z_xin = v_xin / i_xin
let xc = -im(z_xin)
let c_xin = 1 / (2 * pi * f * xc)

* locate index of frequency in question
let idx = 0
let len = length(frequency)

dowhile idx < len
   if frequency[idx] >= 6.5e6
      break
   end
   let idx = idx + 1
end
   
print idx
print frequency[idx]
print z_xin[idx]
print mag(z_xin[idx])
print ph(z_xin[idx])
print ph(z_xin[idx]) * 180 / pi
print c_xin[idx]

.endc

.end
