magic
tech scmos
timestamp 1591540907
<< nwell >>
rect -1 29 22 81
<< metal1 >>
rect 5 76 16 79
rect 6 69 9 73
rect 12 69 15 73
rect 6 62 9 66
rect 12 62 15 66
rect 6 55 9 59
rect 12 55 15 59
rect 6 48 9 52
rect 12 48 15 52
rect 6 41 9 45
rect 12 41 15 45
rect 6 34 9 38
rect 12 34 15 38
rect 6 27 9 31
rect 12 27 15 31
rect 6 20 9 24
rect 12 20 15 24
rect 6 13 9 17
rect 12 13 15 17
rect 6 6 9 10
rect 12 6 15 10
rect 5 0 16 3
rect -2 -10 2 -3
rect 5 -10 9 -3
rect 12 -10 16 -3
rect 19 -10 23 -3
<< bb >>
rect 0 0 21 79
<< labels >>
rlabel metal1 5 0 5 0 2 Gnd
port 3 ne
rlabel nwell 5 30 5 30 2 Vdd
rlabel metal1 5 76 5 76 2 Vdd
port 2 ne
<< end >>
