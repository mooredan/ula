magic
tech scmos
timestamp 1511725328
<< nwell >>
rect 42 123 43 129
rect 97 125 112 127
<< metal1 >>
rect 5 187 9 191
rect 19 186 35 192
rect 45 189 60 192
rect 72 189 87 192
rect 97 187 112 192
rect 123 187 127 191
rect 38 166 50 170
rect 82 166 87 170
rect 5 124 9 128
rect 19 126 34 128
rect 38 120 42 166
rect 101 159 105 170
rect 109 165 113 170
rect 47 126 59 127
rect 73 126 85 127
rect 34 116 42 120
rect 90 93 94 142
rect 97 125 112 127
rect 123 124 127 128
rect 49 86 53 93
rect 90 89 105 93
rect 101 86 105 89
rect 12 82 24 86
rect 5 61 9 65
rect 12 40 16 82
rect 21 63 33 64
rect 38 44 42 86
rect 47 63 59 64
rect 64 57 68 86
rect 82 82 87 86
rect 73 63 85 64
rect 64 53 72 57
rect 90 44 94 86
rect 97 61 113 65
rect 123 61 127 65
rect 38 40 50 44
rect 90 40 102 44
rect 23 33 27 40
rect 79 37 83 40
rect 79 33 109 37
rect 5 -2 9 2
rect 32 1 34 3
rect 21 0 33 1
rect 47 0 59 1
rect 73 0 85 1
rect 19 -3 34 0
rect 45 -3 60 0
rect 72 -3 87 0
rect 97 -3 113 3
rect 123 -2 127 2
<< metal2 >>
rect 5 187 127 191
rect 56 166 87 170
rect 72 159 105 163
rect 90 138 112 142
rect 5 124 127 128
rect 49 89 76 93
rect 38 82 60 86
rect 64 82 87 86
rect 90 82 112 86
rect 5 61 127 65
rect 12 40 34 44
rect 23 33 60 37
rect 5 -2 127 2
<< gv1 >>
rect 6 188 8 190
rect 21 188 23 190
rect 26 188 28 190
rect 31 188 33 190
rect 47 188 49 190
rect 52 188 54 190
rect 57 188 59 190
rect 73 188 75 190
rect 78 188 80 190
rect 83 188 85 190
rect 99 188 101 190
rect 104 188 106 190
rect 109 188 111 190
rect 124 188 126 190
rect 57 167 59 169
rect 84 167 86 169
rect 73 160 75 162
rect 102 160 104 162
rect 91 139 93 141
rect 109 139 111 141
rect 6 125 8 127
rect 21 125 23 127
rect 26 125 28 127
rect 31 125 33 127
rect 47 125 49 127
rect 52 125 54 127
rect 57 125 59 127
rect 73 125 75 127
rect 78 125 80 127
rect 83 125 85 127
rect 99 125 101 127
rect 104 125 106 127
rect 109 125 111 127
rect 124 125 126 127
rect 50 90 52 92
rect 73 90 75 92
rect 39 83 41 85
rect 57 83 59 85
rect 65 83 67 85
rect 84 83 86 85
rect 91 83 93 85
rect 109 83 111 85
rect 6 62 8 64
rect 21 62 23 64
rect 26 62 28 64
rect 31 62 33 64
rect 47 62 49 64
rect 52 62 54 64
rect 57 62 59 64
rect 73 62 75 64
rect 78 62 80 64
rect 83 62 85 64
rect 99 62 101 64
rect 104 62 106 64
rect 109 62 111 64
rect 124 62 126 64
rect 13 41 15 43
rect 31 41 33 43
rect 24 34 26 36
rect 57 34 59 36
rect 6 -1 8 1
rect 21 -1 23 1
rect 26 -1 28 1
rect 31 -1 33 1
rect 47 -1 49 1
rect 52 -1 54 1
rect 57 -1 59 1
rect 73 -1 75 1
rect 78 -1 80 1
rect 83 -1 85 1
rect 99 -1 101 1
rect 104 -1 106 1
rect 109 -1 111 1
rect 124 -1 126 1
use SUBC_1  SUBC_1_1
timestamp 1511591118
transform 1 0 0 0 -1 189
box -1 0 15 65
use INV_B  INV_B_7
timestamp 1511685112
transform 1 0 14 0 -1 189
box -1 0 26 65
use INV_B  INV_B_6
timestamp 1511685112
transform 1 0 40 0 -1 189
box -1 0 26 65
use INV_B  INV_B_8
timestamp 1511685112
transform -1 0 92 0 -1 189
box -1 0 26 65
use INV_B  INV_B_9
timestamp 1511685112
transform 1 0 92 0 -1 189
box -1 0 26 65
use SUBC_1  SUBC_1_3
timestamp 1511591118
transform -1 0 132 0 -1 189
box -1 0 15 65
use SUBC_1  SUBC_1_0
timestamp 1511591118
transform 1 0 0 0 1 63
box -1 0 15 65
use INV_B  INV_B_1
timestamp 1511685112
transform 1 0 14 0 1 63
box -1 0 26 65
use INV_B  INV_B_0
timestamp 1511685112
transform 1 0 40 0 1 63
box -1 0 26 65
use INV_B  INV_B_2
timestamp 1511685112
transform -1 0 92 0 1 63
box -1 0 26 65
use INV_B  INV_B_10
timestamp 1511685112
transform 1 0 92 0 1 63
box -1 0 26 65
use SUBC_1  SUBC_1_4
timestamp 1511591118
transform -1 0 132 0 1 63
box -1 0 15 65
use SUBC_1  SUBC_1_2
timestamp 1511591118
transform 1 0 0 0 -1 63
box -1 0 15 65
use INV_B  INV_B_4
timestamp 1511685112
transform 1 0 14 0 -1 63
box -1 0 26 65
use INV_B  INV_B_3
timestamp 1511685112
transform 1 0 40 0 -1 63
box -1 0 26 65
use INV_B  INV_B_5
timestamp 1511685112
transform -1 0 92 0 -1 63
box -1 0 26 65
use INV_B  INV_B_11
timestamp 1511685112
transform 1 0 92 0 -1 63
box -1 0 26 65
use SUBC_1  SUBC_1_5
timestamp 1511591118
transform -1 0 132 0 -1 63
box -1 0 15 65
<< labels >>
rlabel metal1 111 63 111 63 6 Gnd
port 3 ne
rlabel metal1 111 189 111 189 6 Gnd
port 3 ne
rlabel metal2 10 190 10 190 2 Gnd
port 3 ne
rlabel metal2 10 127 10 127 2 Vdd
rlabel metal2 10 64 10 64 2 Gnd
rlabel metal2 10 1 10 1 2 Vdd
port 4 ne
rlabel metal1 110 167 110 167 2 Out
port 5 ne
rlabel metal1 65 66 65 66 2 n101
<< end >>
