`celldefine
module buf_d (z, a);
  output z;
  input  a;

  buf G1 (z, a);
endmodule
`endcelldefine
