magic
tech amic5n
timestamp 1624630388
<< nwell >>
rect -130 550 580 1495
<< ntransistor >>
rect 225 95 285 400
<< ptransistor >>
rect 225 700 285 1345
<< nselect >>
rect -10 0 460 430
<< pselect >>
rect -10 670 460 1440
<< ndiffusion >>
rect 105 370 225 400
rect 105 320 135 370
rect 185 320 225 370
rect 105 175 225 320
rect 105 125 135 175
rect 185 125 225 175
rect 105 95 225 125
rect 285 370 405 400
rect 285 320 325 370
rect 375 320 405 370
rect 285 175 405 320
rect 285 125 325 175
rect 375 125 405 175
rect 285 95 405 125
<< pdiffusion >>
rect 105 1315 225 1345
rect 105 1265 135 1315
rect 185 1265 225 1315
rect 105 1215 225 1265
rect 105 1165 135 1215
rect 185 1165 225 1215
rect 105 1115 225 1165
rect 105 1065 135 1115
rect 185 1065 225 1115
rect 105 1015 225 1065
rect 105 965 135 1015
rect 185 965 225 1015
rect 105 915 225 965
rect 105 865 135 915
rect 185 865 225 915
rect 105 815 225 865
rect 105 765 135 815
rect 185 765 225 815
rect 105 700 225 765
rect 285 1315 405 1345
rect 285 1265 325 1315
rect 375 1265 405 1315
rect 285 1180 405 1265
rect 285 1130 325 1180
rect 375 1130 405 1180
rect 285 1080 405 1130
rect 285 1030 325 1080
rect 375 1030 405 1080
rect 285 980 405 1030
rect 285 930 325 980
rect 375 930 405 980
rect 285 880 405 930
rect 285 830 325 880
rect 375 830 405 880
rect 285 780 405 830
rect 285 730 325 780
rect 375 730 405 780
rect 285 700 405 730
<< ndcontact >>
rect 135 320 185 370
rect 135 125 185 175
rect 325 320 375 370
rect 325 125 375 175
<< pdcontact >>
rect 135 1265 185 1315
rect 135 1165 185 1215
rect 135 1065 185 1115
rect 135 965 185 1015
rect 135 865 185 915
rect 135 765 185 815
rect 325 1265 375 1315
rect 325 1130 375 1180
rect 325 1030 375 1080
rect 325 930 375 980
rect 325 830 375 880
rect 325 730 375 780
<< polysilicon >>
rect 225 1345 285 1410
rect 225 630 285 700
rect 115 610 285 630
rect 115 560 135 610
rect 185 560 285 610
rect 115 540 285 560
rect 225 400 285 540
rect 225 30 285 95
<< polycontact >>
rect 135 560 185 610
<< metal1 >>
rect 0 1395 450 1485
rect 115 1315 205 1395
rect 115 1265 135 1315
rect 185 1265 205 1315
rect 115 1215 205 1265
rect 115 1165 135 1215
rect 185 1165 205 1215
rect 115 1115 205 1165
rect 115 1065 135 1115
rect 185 1065 205 1115
rect 115 1015 205 1065
rect 115 965 135 1015
rect 185 965 205 1015
rect 115 915 205 965
rect 115 865 135 915
rect 185 865 205 915
rect 115 815 205 865
rect 115 765 135 815
rect 185 765 205 815
rect 115 745 205 765
rect 305 1315 420 1335
rect 305 1265 325 1315
rect 375 1265 420 1315
rect 305 1180 420 1265
rect 305 1130 325 1180
rect 375 1130 420 1180
rect 305 1080 420 1130
rect 305 1030 325 1080
rect 375 1030 420 1080
rect 305 980 420 1030
rect 305 930 325 980
rect 375 930 420 980
rect 305 880 420 930
rect 305 830 325 880
rect 375 830 420 880
rect 305 780 420 830
rect 305 730 325 780
rect 375 730 420 780
rect 30 610 205 685
rect 30 595 135 610
rect 115 560 135 595
rect 185 560 205 610
rect 115 540 205 560
rect 115 370 205 390
rect 115 320 135 370
rect 185 320 205 370
rect 115 175 205 320
rect 115 125 135 175
rect 185 125 205 175
rect 115 45 205 125
rect 305 370 420 730
rect 305 320 325 370
rect 375 320 420 370
rect 305 175 420 320
rect 305 125 325 175
rect 375 125 420 175
rect 305 105 420 125
rect 0 -45 450 45
<< labels >>
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 2 ne
flabel nwell 395 600 395 600 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 335 470 335 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 135 550 135 550 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 3 ne
<< properties >>
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
string FIXED_BBOX 0 0 450 1440
<< end >>
