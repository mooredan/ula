magic
tech amic5n
timestamp 1623521091
<< nwell >>
rect -130 550 1630 1495
<< ntransistor >>
rect 175 250 235 375
rect 385 95 445 400
rect 625 95 685 400
rect 815 95 875 400
rect 1055 95 1115 400
rect 1265 220 1325 345
<< ptransistor >>
rect 175 955 235 1140
rect 385 865 445 1345
rect 625 865 685 1345
rect 815 865 875 1345
rect 1055 865 1115 1345
rect 1265 915 1325 1100
<< nselect >>
rect -10 0 1510 430
<< pselect >>
rect -10 670 1510 1440
<< ndiffusion >>
rect 265 375 385 400
rect 55 345 175 375
rect 55 295 85 345
rect 135 295 175 345
rect 55 250 175 295
rect 235 345 385 375
rect 235 295 295 345
rect 345 295 385 345
rect 235 250 385 295
rect 265 175 385 250
rect 265 125 295 175
rect 345 125 385 175
rect 265 95 385 125
rect 445 95 625 400
rect 685 345 815 400
rect 685 295 725 345
rect 775 295 815 345
rect 685 95 815 295
rect 875 95 1055 400
rect 1115 345 1235 400
rect 1115 295 1155 345
rect 1205 295 1265 345
rect 1115 220 1265 295
rect 1325 315 1445 345
rect 1325 265 1365 315
rect 1415 265 1445 315
rect 1325 220 1445 265
rect 1115 175 1235 220
rect 1115 125 1155 175
rect 1205 125 1235 175
rect 1115 95 1235 125
<< pdiffusion >>
rect 265 1315 385 1345
rect 265 1265 295 1315
rect 345 1265 385 1315
rect 265 1215 385 1265
rect 265 1165 295 1215
rect 345 1165 385 1215
rect 265 1140 385 1165
rect 55 1070 175 1140
rect 55 1020 85 1070
rect 135 1020 175 1070
rect 55 955 175 1020
rect 235 1115 385 1140
rect 235 1065 295 1115
rect 345 1065 385 1115
rect 235 985 385 1065
rect 235 955 295 985
rect 265 935 295 955
rect 345 935 385 985
rect 265 865 385 935
rect 445 865 625 1345
rect 685 1315 815 1345
rect 685 1265 725 1315
rect 775 1265 815 1315
rect 685 1215 815 1265
rect 685 1165 725 1215
rect 775 1165 815 1215
rect 685 1115 815 1165
rect 685 1065 725 1115
rect 775 1065 815 1115
rect 685 865 815 1065
rect 875 865 1055 1345
rect 1115 1315 1235 1345
rect 1115 1265 1155 1315
rect 1205 1265 1235 1315
rect 1115 1215 1235 1265
rect 1115 1165 1155 1215
rect 1205 1165 1235 1215
rect 1115 1115 1235 1165
rect 1115 1065 1155 1115
rect 1205 1100 1235 1115
rect 1205 1065 1265 1100
rect 1115 985 1265 1065
rect 1115 935 1155 985
rect 1205 935 1265 985
rect 1115 915 1265 935
rect 1325 1030 1445 1100
rect 1325 980 1365 1030
rect 1415 980 1445 1030
rect 1325 915 1445 980
rect 1115 865 1235 915
<< ndcontact >>
rect 85 295 135 345
rect 295 295 345 345
rect 295 125 345 175
rect 725 295 775 345
rect 1155 295 1205 345
rect 1365 265 1415 315
rect 1155 125 1205 175
<< pdcontact >>
rect 295 1265 345 1315
rect 295 1165 345 1215
rect 85 1020 135 1070
rect 295 1065 345 1115
rect 295 935 345 985
rect 725 1265 775 1315
rect 725 1165 775 1215
rect 725 1065 775 1115
rect 1155 1265 1205 1315
rect 1155 1165 1205 1215
rect 1155 1065 1205 1115
rect 1155 935 1205 985
rect 1365 980 1415 1030
<< polysilicon >>
rect 385 1345 445 1410
rect 625 1345 685 1410
rect 815 1345 875 1410
rect 1055 1345 1115 1410
rect 175 1140 235 1205
rect 175 525 235 955
rect 1265 1100 1325 1165
rect 385 525 445 865
rect 625 685 685 865
rect 535 665 685 685
rect 535 615 555 665
rect 605 615 685 665
rect 535 595 685 615
rect 815 845 875 865
rect 815 825 965 845
rect 815 775 895 825
rect 945 775 965 825
rect 815 755 965 775
rect 175 505 445 525
rect 175 455 275 505
rect 325 455 445 505
rect 175 435 445 455
rect 535 505 685 525
rect 535 455 555 505
rect 605 455 685 505
rect 535 435 685 455
rect 175 375 235 435
rect 385 400 445 435
rect 625 400 685 435
rect 815 400 875 755
rect 1055 685 1115 865
rect 1265 685 1325 915
rect 965 665 1325 685
rect 965 615 985 665
rect 1035 615 1175 665
rect 1225 615 1325 665
rect 965 595 1325 615
rect 1055 505 1205 525
rect 1055 455 1135 505
rect 1185 455 1205 505
rect 1055 435 1205 455
rect 1055 400 1115 435
rect 175 185 235 250
rect 1265 345 1325 595
rect 1265 155 1325 220
rect 385 30 445 95
rect 625 30 685 95
rect 815 30 875 95
rect 1055 30 1115 95
<< polycontact >>
rect 555 615 605 665
rect 895 775 945 825
rect 275 455 325 505
rect 555 455 605 505
rect 985 615 1035 665
rect 1175 615 1225 665
rect 1135 455 1185 505
<< metal1 >>
rect 0 1395 1500 1485
rect 275 1315 365 1395
rect 275 1265 295 1315
rect 345 1265 365 1315
rect 275 1215 365 1265
rect 275 1165 295 1215
rect 345 1165 365 1215
rect 275 1115 365 1165
rect 65 1070 155 1100
rect 65 1020 85 1070
rect 135 1020 155 1070
rect 65 825 155 1020
rect 275 1065 295 1115
rect 345 1065 365 1115
rect 275 985 365 1065
rect 275 935 295 985
rect 345 935 365 985
rect 275 915 365 935
rect 705 1315 795 1335
rect 705 1265 725 1315
rect 775 1265 795 1315
rect 705 1215 795 1265
rect 705 1165 725 1215
rect 775 1165 795 1215
rect 705 1115 795 1165
rect 705 1065 725 1115
rect 775 1065 795 1115
rect 65 775 85 825
rect 135 775 155 825
rect 65 345 155 775
rect 535 665 625 685
rect 535 615 555 665
rect 605 615 625 665
rect 535 595 625 615
rect 255 505 430 525
rect 255 455 275 505
rect 325 455 430 505
rect 255 435 430 455
rect 535 505 625 525
rect 535 455 555 505
rect 605 455 625 505
rect 65 295 85 345
rect 135 295 155 345
rect 65 260 155 295
rect 275 345 365 365
rect 275 295 295 345
rect 345 295 365 345
rect 275 175 365 295
rect 275 125 295 175
rect 345 125 365 175
rect 275 45 365 125
rect 535 205 625 455
rect 705 345 795 1065
rect 1135 1315 1225 1395
rect 1135 1265 1155 1315
rect 1205 1265 1225 1315
rect 1135 1215 1225 1265
rect 1135 1165 1155 1215
rect 1205 1165 1225 1215
rect 1135 1115 1225 1165
rect 1135 1065 1155 1115
rect 1205 1065 1225 1115
rect 1135 985 1225 1065
rect 1135 935 1155 985
rect 1205 935 1225 985
rect 1135 915 1225 935
rect 1345 1030 1435 1060
rect 1345 980 1365 1030
rect 1415 980 1435 1030
rect 875 825 965 845
rect 875 775 895 825
rect 945 775 965 825
rect 875 755 965 775
rect 705 295 725 345
rect 775 295 795 345
rect 705 275 795 295
rect 965 665 1245 685
rect 965 615 985 665
rect 1035 615 1175 665
rect 1225 615 1245 665
rect 965 595 1245 615
rect 965 205 1055 595
rect 1345 525 1435 980
rect 1115 505 1435 525
rect 1115 455 1135 505
rect 1185 455 1435 505
rect 1115 435 1435 455
rect 535 115 1055 205
rect 1135 345 1225 365
rect 1135 295 1155 345
rect 1205 295 1225 345
rect 1135 175 1225 295
rect 1345 315 1435 435
rect 1345 265 1365 315
rect 1415 265 1435 315
rect 1345 230 1435 265
rect 1135 125 1155 175
rect 1205 125 1225 175
rect 1135 45 1225 125
rect 0 -45 1500 45
<< via1 >>
rect 85 775 135 825
rect 555 615 605 665
rect 895 775 945 825
rect 1135 455 1185 505
<< metal2 >>
rect 65 825 965 845
rect 65 775 85 825
rect 135 775 895 825
rect 945 775 965 825
rect 65 755 965 775
rect 535 665 795 685
rect 535 615 555 665
rect 605 615 795 665
rect 535 595 795 615
rect 705 525 795 595
rect 705 505 1205 525
rect 705 455 1135 505
rect 1185 455 1205 505
rect 705 435 1205 455
<< labels >>
flabel polysilicon 645 460 645 460 1 FreeSans 200 0 0 0 b
flabel polysilicon 400 650 400 650 1 FreeSans 200 0 0 0 a
flabel polysilicon 640 650 640 650 1 FreeSans 200 0 0 0 nb
flabel polysilicon 835 465 835 465 1 FreeSans 200 0 0 0 na
flabel polysilicon 1080 460 1080 460 1 FreeSans 200 0 0 0 nb
flabel polysilicon 1080 640 1080 640 1 FreeSans 200 0 0 0 b
flabel metal1 s 310 445 310 445 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 1121 630 1121 630 2 FreeSans 400 0 0 0 b
port 2 ne
flabel metal1 s 730 940 730 940 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 75 -20 75 -20 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 55 1420 55 1420 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel nwell -35 610 -35 610 2 FreeSans 400 0 0 0 vdd
flabel ndiffusion s 465 210 465 210 2 FreeSans 200 0 0 0 n1
flabel ndiffusion s 905 245 905 245 2 FreeSans 200 0 0 0 n2
flabel pdiffusion s 500 1015 500 1015 2 FreeSans 200 0 0 0 p1
flabel pdiffusion s 920 1085 920 1085 2 FreeSans 200 0 0 0 p2
<< end >>
