magic
tech amic5n
timestamp 1622213957
<< nwell >>
rect -105 805 495 2455
rect 1245 760 1845 2295
rect 2595 720 3195 2135
rect 3945 675 4545 1975
rect 5295 635 5895 1815
rect 6645 590 7245 1655
rect 7995 550 8595 1495
rect 9345 505 9945 1335
rect 10695 460 11295 1175
rect 12045 415 12645 1015
rect 13545 370 14145 855
<< ntransistor >>
rect 165 95 225 655
rect 1515 95 1575 610
rect 2865 95 2925 570
rect 4215 95 4275 525
rect 5565 95 5625 485
rect 6915 95 6975 440
rect 8265 95 8325 400
rect 9615 95 9675 355
rect 10965 95 11025 310
rect 12315 95 12375 265
rect 13815 95 13875 220
<< ptransistor >>
rect 165 955 225 2305
rect 1515 910 1575 2145
rect 2865 870 2925 1985
rect 4215 825 4275 1825
rect 5565 785 5625 1665
rect 6915 740 6975 1505
rect 8265 700 8325 1345
rect 9615 655 9675 1185
rect 10965 610 11025 1025
rect 12315 565 12375 865
rect 13815 520 13875 705
<< nselect >>
rect 0 0 390 685
rect 1350 0 1740 640
rect 2700 0 3090 600
rect 4050 0 4440 555
rect 5400 0 5790 515
rect 6750 0 7140 470
rect 8100 0 8490 430
rect 9450 0 9840 385
rect 10800 0 11190 340
rect 12150 0 12540 295
rect 13650 0 14040 250
<< pselect >>
rect 0 925 390 2400
rect 1350 880 1740 2240
rect 2700 840 3090 2080
rect 4050 795 4440 1920
rect 5400 755 5790 1760
rect 6750 710 7140 1600
rect 8100 670 8490 1440
rect 9450 625 9840 1280
rect 10800 580 11190 1120
rect 12150 535 12540 960
rect 13650 490 14040 800
<< ndiffusion >>
rect 45 175 165 655
rect 45 125 75 175
rect 125 125 165 175
rect 45 95 165 125
rect 225 175 345 655
rect 225 125 265 175
rect 315 125 345 175
rect 225 95 345 125
rect 1395 175 1515 610
rect 1395 125 1425 175
rect 1475 125 1515 175
rect 1395 95 1515 125
rect 1575 175 1695 610
rect 1575 125 1615 175
rect 1665 125 1695 175
rect 1575 95 1695 125
rect 2745 175 2865 570
rect 2745 125 2775 175
rect 2825 125 2865 175
rect 2745 95 2865 125
rect 2925 175 3045 570
rect 2925 125 2965 175
rect 3015 125 3045 175
rect 2925 95 3045 125
rect 4095 175 4215 525
rect 4095 125 4125 175
rect 4175 125 4215 175
rect 4095 95 4215 125
rect 4275 175 4395 525
rect 4275 125 4315 175
rect 4365 125 4395 175
rect 4275 95 4395 125
rect 5445 175 5565 485
rect 5445 125 5475 175
rect 5525 125 5565 175
rect 5445 95 5565 125
rect 5625 175 5745 485
rect 5625 125 5665 175
rect 5715 125 5745 175
rect 5625 95 5745 125
rect 6795 175 6915 440
rect 6795 125 6825 175
rect 6875 125 6915 175
rect 6795 95 6915 125
rect 6975 175 7095 440
rect 6975 125 7015 175
rect 7065 125 7095 175
rect 6975 95 7095 125
rect 8145 175 8265 400
rect 8145 125 8175 175
rect 8225 125 8265 175
rect 8145 95 8265 125
rect 8325 175 8445 400
rect 8325 125 8365 175
rect 8415 125 8445 175
rect 8325 95 8445 125
rect 9495 175 9615 355
rect 9495 125 9525 175
rect 9575 125 9615 175
rect 9495 95 9615 125
rect 9675 175 9795 355
rect 9675 125 9715 175
rect 9765 125 9795 175
rect 9675 95 9795 125
rect 10845 175 10965 310
rect 10845 125 10875 175
rect 10925 125 10965 175
rect 10845 95 10965 125
rect 11025 175 11145 310
rect 11025 125 11065 175
rect 11115 125 11145 175
rect 11025 95 11145 125
rect 12195 175 12315 265
rect 12195 125 12225 175
rect 12275 125 12315 175
rect 12195 95 12315 125
rect 12375 175 12495 265
rect 12375 125 12415 175
rect 12465 125 12495 175
rect 12375 95 12495 125
rect 13695 175 13815 220
rect 13695 125 13725 175
rect 13775 125 13815 175
rect 13695 95 13815 125
rect 13875 175 13995 220
rect 13875 125 13915 175
rect 13965 125 13995 175
rect 13875 95 13995 125
<< pdiffusion >>
rect 45 2275 165 2305
rect 45 2225 75 2275
rect 125 2225 165 2275
rect 45 1035 165 2225
rect 45 985 75 1035
rect 125 985 165 1035
rect 45 955 165 985
rect 225 2275 345 2305
rect 225 2225 265 2275
rect 315 2225 345 2275
rect 225 1035 345 2225
rect 225 985 265 1035
rect 315 985 345 1035
rect 225 955 345 985
rect 1395 2115 1515 2145
rect 1395 2065 1425 2115
rect 1475 2065 1515 2115
rect 1395 990 1515 2065
rect 1395 940 1425 990
rect 1475 940 1515 990
rect 1395 910 1515 940
rect 1575 2115 1695 2145
rect 1575 2065 1615 2115
rect 1665 2065 1695 2115
rect 1575 990 1695 2065
rect 1575 940 1615 990
rect 1665 940 1695 990
rect 1575 910 1695 940
rect 2745 1955 2865 1985
rect 2745 1905 2775 1955
rect 2825 1905 2865 1955
rect 2745 950 2865 1905
rect 2745 900 2775 950
rect 2825 900 2865 950
rect 2745 870 2865 900
rect 2925 1955 3045 1985
rect 2925 1905 2965 1955
rect 3015 1905 3045 1955
rect 2925 950 3045 1905
rect 2925 900 2965 950
rect 3015 900 3045 950
rect 2925 870 3045 900
rect 4095 1795 4215 1825
rect 4095 1745 4125 1795
rect 4175 1745 4215 1795
rect 4095 905 4215 1745
rect 4095 855 4125 905
rect 4175 855 4215 905
rect 4095 825 4215 855
rect 4275 1795 4395 1825
rect 4275 1745 4315 1795
rect 4365 1745 4395 1795
rect 4275 905 4395 1745
rect 4275 855 4315 905
rect 4365 855 4395 905
rect 4275 825 4395 855
rect 5445 1635 5565 1665
rect 5445 1585 5475 1635
rect 5525 1585 5565 1635
rect 5445 865 5565 1585
rect 5445 815 5475 865
rect 5525 815 5565 865
rect 5445 785 5565 815
rect 5625 1635 5745 1665
rect 5625 1585 5665 1635
rect 5715 1585 5745 1635
rect 5625 865 5745 1585
rect 5625 815 5665 865
rect 5715 815 5745 865
rect 5625 785 5745 815
rect 6795 1475 6915 1505
rect 6795 1425 6825 1475
rect 6875 1425 6915 1475
rect 6795 820 6915 1425
rect 6795 770 6825 820
rect 6875 770 6915 820
rect 6795 740 6915 770
rect 6975 1475 7095 1505
rect 6975 1425 7015 1475
rect 7065 1425 7095 1475
rect 6975 820 7095 1425
rect 6975 770 7015 820
rect 7065 770 7095 820
rect 6975 740 7095 770
rect 8145 1315 8265 1345
rect 8145 1265 8175 1315
rect 8225 1265 8265 1315
rect 8145 780 8265 1265
rect 8145 730 8175 780
rect 8225 730 8265 780
rect 8145 700 8265 730
rect 8325 1315 8445 1345
rect 8325 1265 8365 1315
rect 8415 1265 8445 1315
rect 8325 780 8445 1265
rect 8325 730 8365 780
rect 8415 730 8445 780
rect 8325 700 8445 730
rect 9495 1155 9615 1185
rect 9495 1105 9525 1155
rect 9575 1105 9615 1155
rect 9495 735 9615 1105
rect 9495 685 9525 735
rect 9575 685 9615 735
rect 9495 655 9615 685
rect 9675 1155 9795 1185
rect 9675 1105 9715 1155
rect 9765 1105 9795 1155
rect 9675 735 9795 1105
rect 9675 685 9715 735
rect 9765 685 9795 735
rect 9675 655 9795 685
rect 10845 995 10965 1025
rect 10845 945 10875 995
rect 10925 945 10965 995
rect 10845 690 10965 945
rect 10845 640 10875 690
rect 10925 640 10965 690
rect 10845 610 10965 640
rect 11025 995 11145 1025
rect 11025 945 11065 995
rect 11115 945 11145 995
rect 11025 690 11145 945
rect 11025 640 11065 690
rect 11115 640 11145 690
rect 11025 610 11145 640
rect 12195 835 12315 865
rect 12195 785 12225 835
rect 12275 785 12315 835
rect 12195 645 12315 785
rect 12195 595 12225 645
rect 12275 595 12315 645
rect 12195 565 12315 595
rect 12375 835 12495 865
rect 12375 785 12415 835
rect 12465 785 12495 835
rect 12375 645 12495 785
rect 12375 595 12415 645
rect 12465 595 12495 645
rect 12375 565 12495 595
rect 13695 600 13815 705
rect 13695 550 13725 600
rect 13775 550 13815 600
rect 13695 520 13815 550
rect 13875 600 13995 705
rect 13875 550 13915 600
rect 13965 550 13995 600
rect 13875 520 13995 550
<< ndcontact >>
rect 75 125 125 175
rect 265 125 315 175
rect 1425 125 1475 175
rect 1615 125 1665 175
rect 2775 125 2825 175
rect 2965 125 3015 175
rect 4125 125 4175 175
rect 4315 125 4365 175
rect 5475 125 5525 175
rect 5665 125 5715 175
rect 6825 125 6875 175
rect 7015 125 7065 175
rect 8175 125 8225 175
rect 8365 125 8415 175
rect 9525 125 9575 175
rect 9715 125 9765 175
rect 10875 125 10925 175
rect 11065 125 11115 175
rect 12225 125 12275 175
rect 12415 125 12465 175
rect 13725 125 13775 175
rect 13915 125 13965 175
<< pdcontact >>
rect 75 2225 125 2275
rect 75 985 125 1035
rect 265 2225 315 2275
rect 265 985 315 1035
rect 1425 2065 1475 2115
rect 1425 940 1475 990
rect 1615 2065 1665 2115
rect 1615 940 1665 990
rect 2775 1905 2825 1955
rect 2775 900 2825 950
rect 2965 1905 3015 1955
rect 2965 900 3015 950
rect 4125 1745 4175 1795
rect 4125 855 4175 905
rect 4315 1745 4365 1795
rect 4315 855 4365 905
rect 5475 1585 5525 1635
rect 5475 815 5525 865
rect 5665 1585 5715 1635
rect 5665 815 5715 865
rect 6825 1425 6875 1475
rect 6825 770 6875 820
rect 7015 1425 7065 1475
rect 7015 770 7065 820
rect 8175 1265 8225 1315
rect 8175 730 8225 780
rect 8365 1265 8415 1315
rect 8365 730 8415 780
rect 9525 1105 9575 1155
rect 9525 685 9575 735
rect 9715 1105 9765 1155
rect 9715 685 9765 735
rect 10875 945 10925 995
rect 10875 640 10925 690
rect 11065 945 11115 995
rect 11065 640 11115 690
rect 12225 785 12275 835
rect 12225 595 12275 645
rect 12415 785 12465 835
rect 12415 595 12465 645
rect 13725 550 13775 600
rect 13915 550 13965 600
<< polysilicon >>
rect 165 2305 225 2370
rect 1515 2145 1575 2210
rect 165 845 225 955
rect 2865 1985 2925 2050
rect 55 825 225 845
rect 55 775 75 825
rect 125 775 225 825
rect 1515 800 1575 910
rect 4215 1825 4275 1890
rect 55 755 225 775
rect 165 655 225 755
rect 1405 780 1575 800
rect 1405 730 1425 780
rect 1475 730 1575 780
rect 2865 760 2925 870
rect 5565 1665 5625 1730
rect 1405 710 1575 730
rect 1515 610 1575 710
rect 2755 740 2925 760
rect 2755 690 2775 740
rect 2825 690 2925 740
rect 4215 715 4275 825
rect 6915 1505 6975 1570
rect 2755 670 2925 690
rect 2865 570 2925 670
rect 4105 695 4275 715
rect 4105 645 4125 695
rect 4175 645 4275 695
rect 5565 675 5625 785
rect 8265 1345 8325 1410
rect 4105 625 4275 645
rect 4215 525 4275 625
rect 5455 655 5625 675
rect 5455 605 5475 655
rect 5525 605 5625 655
rect 6915 630 6975 740
rect 9615 1185 9675 1250
rect 5455 585 5625 605
rect 5565 485 5625 585
rect 6805 610 6975 630
rect 6805 560 6825 610
rect 6875 560 6975 610
rect 8265 590 8325 700
rect 10965 1025 11025 1090
rect 6805 540 6975 560
rect 6915 440 6975 540
rect 8155 570 8325 590
rect 8155 520 8175 570
rect 8225 520 8325 570
rect 9615 545 9675 655
rect 12315 865 12375 930
rect 8155 500 8325 520
rect 8265 400 8325 500
rect 9505 525 9675 545
rect 9505 475 9525 525
rect 9575 475 9675 525
rect 10965 500 11025 610
rect 13815 705 13875 770
rect 9505 455 9675 475
rect 9615 355 9675 455
rect 10855 480 11025 500
rect 10855 430 10875 480
rect 10925 430 11025 480
rect 12315 455 12375 565
rect 10855 410 11025 430
rect 10965 310 11025 410
rect 12205 435 12375 455
rect 12205 385 12225 435
rect 12275 385 12375 435
rect 13815 410 13875 520
rect 12205 365 12375 385
rect 12315 265 12375 365
rect 13705 390 13875 410
rect 13705 340 13725 390
rect 13775 340 13875 390
rect 13705 320 13875 340
rect 13815 220 13875 320
rect 165 30 225 95
rect 1515 30 1575 95
rect 2865 30 2925 95
rect 4215 30 4275 95
rect 5565 30 5625 95
rect 6915 30 6975 95
rect 8265 30 8325 95
rect 9615 30 9675 95
rect 10965 30 11025 95
rect 12315 30 12375 95
rect 13815 30 13875 95
<< polycontact >>
rect 75 775 125 825
rect 1425 730 1475 780
rect 2775 690 2825 740
rect 4125 645 4175 695
rect 5475 605 5525 655
rect 6825 560 6875 610
rect 8175 520 8225 570
rect 9525 475 9575 525
rect 10875 430 10925 480
rect 12225 385 12275 435
rect 13725 340 13775 390
<< metal1 >>
rect 0 2425 390 2445
rect 0 2375 295 2425
rect 345 2375 390 2425
rect 0 2355 390 2375
rect 55 2275 145 2355
rect 55 2225 75 2275
rect 125 2225 145 2275
rect 55 1035 145 2225
rect 55 985 75 1035
rect 125 985 145 1035
rect 55 965 145 985
rect 245 2275 335 2295
rect 245 2225 265 2275
rect 315 2225 335 2275
rect 245 1035 335 2225
rect 1350 2265 1740 2285
rect 1350 2215 1650 2265
rect 1700 2215 1740 2265
rect 1350 2195 1740 2215
rect 245 985 265 1035
rect 315 985 335 1035
rect 55 825 145 845
rect 55 775 75 825
rect 125 775 145 825
rect 55 755 145 775
rect 55 175 145 645
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 245 175 335 985
rect 1405 2115 1495 2195
rect 1405 2065 1425 2115
rect 1475 2065 1495 2115
rect 1405 990 1495 2065
rect 1405 940 1425 990
rect 1475 940 1495 990
rect 1405 920 1495 940
rect 1595 2115 1685 2135
rect 1595 2065 1615 2115
rect 1665 2065 1685 2115
rect 1595 990 1685 2065
rect 2700 2105 3090 2125
rect 2700 2055 2990 2105
rect 3040 2055 3090 2105
rect 2700 2035 3090 2055
rect 1595 940 1615 990
rect 1665 940 1685 990
rect 1405 780 1495 800
rect 1405 730 1425 780
rect 1475 730 1495 780
rect 1405 710 1495 730
rect 245 125 265 175
rect 315 125 335 175
rect 245 105 335 125
rect 1405 175 1495 600
rect 1405 125 1425 175
rect 1475 125 1495 175
rect 1405 45 1495 125
rect 1595 175 1685 940
rect 2755 1955 2845 2035
rect 2755 1905 2775 1955
rect 2825 1905 2845 1955
rect 2755 950 2845 1905
rect 2755 900 2775 950
rect 2825 900 2845 950
rect 2755 880 2845 900
rect 2945 1955 3035 1975
rect 2945 1905 2965 1955
rect 3015 1905 3035 1955
rect 2945 950 3035 1905
rect 4050 1945 4440 1965
rect 4050 1895 4345 1945
rect 4395 1895 4440 1945
rect 4050 1875 4440 1895
rect 2945 900 2965 950
rect 3015 900 3035 950
rect 2755 740 2845 760
rect 2755 690 2775 740
rect 2825 690 2845 740
rect 2755 670 2845 690
rect 1595 125 1615 175
rect 1665 125 1685 175
rect 1595 105 1685 125
rect 2755 175 2845 560
rect 2755 125 2775 175
rect 2825 125 2845 175
rect 2755 45 2845 125
rect 2945 175 3035 900
rect 4105 1795 4195 1875
rect 4105 1745 4125 1795
rect 4175 1745 4195 1795
rect 4105 905 4195 1745
rect 4105 855 4125 905
rect 4175 855 4195 905
rect 4105 835 4195 855
rect 4295 1795 4385 1815
rect 4295 1745 4315 1795
rect 4365 1745 4385 1795
rect 4295 905 4385 1745
rect 5400 1785 5790 1805
rect 5400 1735 5685 1785
rect 5735 1735 5790 1785
rect 5400 1715 5790 1735
rect 4295 855 4315 905
rect 4365 855 4385 905
rect 4105 695 4195 715
rect 4105 645 4125 695
rect 4175 645 4195 695
rect 4105 625 4195 645
rect 2945 125 2965 175
rect 3015 125 3035 175
rect 2945 105 3035 125
rect 4105 175 4195 515
rect 4105 125 4125 175
rect 4175 125 4195 175
rect 4105 45 4195 125
rect 4295 175 4385 855
rect 5455 1635 5545 1715
rect 5455 1585 5475 1635
rect 5525 1585 5545 1635
rect 5455 865 5545 1585
rect 5455 815 5475 865
rect 5525 815 5545 865
rect 5455 795 5545 815
rect 5645 1635 5735 1655
rect 5645 1585 5665 1635
rect 5715 1585 5735 1635
rect 5645 865 5735 1585
rect 6750 1625 7140 1645
rect 6750 1575 7040 1625
rect 7090 1575 7140 1625
rect 6750 1555 7140 1575
rect 5645 815 5665 865
rect 5715 815 5735 865
rect 5455 655 5545 675
rect 5455 605 5475 655
rect 5525 605 5545 655
rect 5455 585 5545 605
rect 4295 125 4315 175
rect 4365 125 4385 175
rect 4295 105 4385 125
rect 5455 175 5545 475
rect 5455 125 5475 175
rect 5525 125 5545 175
rect 5455 45 5545 125
rect 5645 175 5735 815
rect 6805 1475 6895 1555
rect 6805 1425 6825 1475
rect 6875 1425 6895 1475
rect 6805 820 6895 1425
rect 6805 770 6825 820
rect 6875 770 6895 820
rect 6805 750 6895 770
rect 6995 1475 7085 1495
rect 6995 1425 7015 1475
rect 7065 1425 7085 1475
rect 6995 820 7085 1425
rect 8100 1465 8490 1485
rect 8100 1415 8385 1465
rect 8435 1415 8490 1465
rect 8100 1395 8490 1415
rect 6995 770 7015 820
rect 7065 770 7085 820
rect 6805 610 6895 630
rect 6805 560 6825 610
rect 6875 560 6895 610
rect 6805 540 6895 560
rect 5645 125 5665 175
rect 5715 125 5735 175
rect 5645 105 5735 125
rect 6805 175 6895 430
rect 6805 125 6825 175
rect 6875 125 6895 175
rect 6805 45 6895 125
rect 6995 175 7085 770
rect 8155 1315 8245 1395
rect 8155 1265 8175 1315
rect 8225 1265 8245 1315
rect 8155 780 8245 1265
rect 8155 730 8175 780
rect 8225 730 8245 780
rect 8155 710 8245 730
rect 8345 1315 8435 1335
rect 8345 1265 8365 1315
rect 8415 1265 8435 1315
rect 8345 780 8435 1265
rect 9450 1305 9840 1325
rect 9450 1255 9735 1305
rect 9785 1255 9840 1305
rect 9450 1235 9840 1255
rect 8345 730 8365 780
rect 8415 730 8435 780
rect 8155 570 8245 590
rect 8155 520 8175 570
rect 8225 520 8245 570
rect 8155 500 8245 520
rect 6995 125 7015 175
rect 7065 125 7085 175
rect 6995 105 7085 125
rect 8155 175 8245 390
rect 8155 125 8175 175
rect 8225 125 8245 175
rect 8155 45 8245 125
rect 8345 175 8435 730
rect 9505 1155 9595 1235
rect 9505 1105 9525 1155
rect 9575 1105 9595 1155
rect 9505 735 9595 1105
rect 9505 685 9525 735
rect 9575 685 9595 735
rect 9505 665 9595 685
rect 9695 1155 9785 1175
rect 9695 1105 9715 1155
rect 9765 1105 9785 1155
rect 9695 735 9785 1105
rect 10800 1145 11190 1165
rect 10800 1095 11070 1145
rect 11120 1095 11190 1145
rect 10800 1075 11190 1095
rect 9695 685 9715 735
rect 9765 685 9785 735
rect 9505 525 9595 545
rect 9505 475 9525 525
rect 9575 475 9595 525
rect 9505 455 9595 475
rect 8345 125 8365 175
rect 8415 125 8435 175
rect 8345 105 8435 125
rect 9505 175 9595 345
rect 9505 125 9525 175
rect 9575 125 9595 175
rect 9505 45 9595 125
rect 9695 175 9785 685
rect 10855 995 10945 1075
rect 10855 945 10875 995
rect 10925 945 10945 995
rect 10855 690 10945 945
rect 10855 640 10875 690
rect 10925 640 10945 690
rect 10855 620 10945 640
rect 11045 995 11135 1015
rect 11045 945 11065 995
rect 11115 945 11135 995
rect 11045 690 11135 945
rect 12150 985 12540 1005
rect 12150 935 12455 985
rect 12505 935 12540 985
rect 12150 915 12540 935
rect 11045 640 11065 690
rect 11115 640 11135 690
rect 10855 480 10945 500
rect 10855 430 10875 480
rect 10925 430 10945 480
rect 10855 410 10945 430
rect 9695 125 9715 175
rect 9765 125 9785 175
rect 9695 105 9785 125
rect 10855 175 10945 300
rect 10855 125 10875 175
rect 10925 125 10945 175
rect 10855 45 10945 125
rect 11045 175 11135 640
rect 12205 835 12295 915
rect 12205 785 12225 835
rect 12275 785 12295 835
rect 12205 645 12295 785
rect 12205 595 12225 645
rect 12275 595 12295 645
rect 12205 575 12295 595
rect 12395 835 12485 855
rect 12395 785 12415 835
rect 12465 785 12485 835
rect 12395 645 12485 785
rect 13650 825 14040 845
rect 13650 775 13955 825
rect 14005 775 14040 825
rect 13650 755 14040 775
rect 12395 595 12415 645
rect 12465 595 12485 645
rect 12205 435 12295 455
rect 12205 385 12225 435
rect 12275 385 12295 435
rect 12205 365 12295 385
rect 11045 125 11065 175
rect 11115 125 11135 175
rect 11045 105 11135 125
rect 12205 175 12295 255
rect 12205 125 12225 175
rect 12275 125 12295 175
rect 12205 45 12295 125
rect 12395 175 12485 595
rect 13705 600 13795 755
rect 13705 550 13725 600
rect 13775 550 13795 600
rect 13705 530 13795 550
rect 13895 600 13985 695
rect 13895 550 13915 600
rect 13965 550 13985 600
rect 13705 390 13795 410
rect 13705 340 13725 390
rect 13775 340 13795 390
rect 13705 320 13795 340
rect 12395 125 12415 175
rect 12465 125 12485 175
rect 12395 105 12485 125
rect 13705 175 13795 210
rect 13705 125 13725 175
rect 13775 125 13795 175
rect 13705 45 13795 125
rect 13895 175 13985 550
rect 13895 125 13915 175
rect 13965 125 13985 175
rect 13895 105 13985 125
rect 0 25 390 45
rect 0 -25 310 25
rect 360 -25 390 25
rect 0 -45 390 -25
rect 1350 25 1740 45
rect 1350 -25 1660 25
rect 1710 -25 1740 25
rect 1350 -45 1740 -25
rect 2700 25 3090 45
rect 2700 -25 2995 25
rect 3045 -25 3090 25
rect 2700 -45 3090 -25
rect 4050 25 4440 45
rect 4050 -25 4335 25
rect 4385 -25 4440 25
rect 4050 -45 4440 -25
rect 5400 25 5790 45
rect 5400 -25 5675 25
rect 5725 -25 5790 25
rect 5400 -45 5790 -25
rect 6750 25 7140 45
rect 6750 -25 7010 25
rect 7060 -25 7140 25
rect 6750 -45 7140 -25
rect 8100 25 8490 45
rect 8100 -25 8350 25
rect 8400 -25 8490 25
rect 8100 -45 8490 -25
rect 9450 25 9840 45
rect 9450 -25 9685 25
rect 9735 -25 9840 25
rect 9450 -45 9840 -25
rect 10800 25 11190 45
rect 10800 -25 11025 25
rect 11075 -25 11190 25
rect 10800 -45 11190 -25
rect 12150 25 12540 45
rect 12150 -25 12460 25
rect 12510 -25 12540 25
rect 12150 -45 12540 -25
rect 13650 -45 14040 45
<< via1 >>
rect 295 2375 345 2425
rect 1650 2215 1700 2265
rect 2990 2055 3040 2105
rect 4345 1895 4395 1945
rect 5685 1735 5735 1785
rect 7040 1575 7090 1625
rect 8385 1415 8435 1465
rect 9735 1255 9785 1305
rect 11070 1095 11120 1145
rect 12455 935 12505 985
rect 13955 775 14005 825
rect 310 -25 360 25
rect 1660 -25 1710 25
rect 2995 -25 3045 25
rect 4335 -25 4385 25
rect 5675 -25 5725 25
rect 7010 -25 7060 25
rect 8350 -25 8400 25
rect 9685 -25 9735 25
rect 11025 -25 11075 25
rect 12460 -25 12510 25
<< metal2 >>
rect -50 2425 12795 2445
rect -50 2375 295 2425
rect 345 2375 12795 2425
rect -50 2355 12795 2375
rect 12685 2285 12795 2355
rect -50 2265 12795 2285
rect -50 2215 1650 2265
rect 1700 2215 12795 2265
rect -50 2195 12795 2215
rect 12685 2125 12795 2195
rect -50 2105 12795 2125
rect -50 2055 2990 2105
rect 3040 2055 12795 2105
rect -50 2035 12795 2055
rect 12685 1965 12795 2035
rect -50 1945 12795 1965
rect -50 1895 4345 1945
rect 4395 1895 12795 1945
rect -50 1875 12795 1895
rect 12685 1805 12795 1875
rect -50 1785 12795 1805
rect -50 1735 5685 1785
rect 5735 1735 12795 1785
rect -50 1715 12795 1735
rect 12685 1645 12795 1715
rect -50 1625 12795 1645
rect -50 1575 7040 1625
rect 7090 1575 12795 1625
rect -50 1555 12795 1575
rect 12685 1485 12795 1555
rect -50 1465 12795 1485
rect -50 1415 8385 1465
rect 8435 1415 12795 1465
rect -50 1395 12795 1415
rect 12685 1325 12795 1395
rect -50 1305 12795 1325
rect -50 1255 9735 1305
rect 9785 1255 12795 1305
rect -50 1235 12795 1255
rect 12685 1165 12795 1235
rect -50 1145 12795 1165
rect -50 1095 11070 1145
rect 11120 1095 12795 1145
rect -50 1075 12795 1095
rect 12685 1005 12795 1075
rect -50 985 12795 1005
rect -50 935 12455 985
rect 12505 935 12795 985
rect -50 915 12795 935
rect -50 825 14065 845
rect -50 775 13955 825
rect 14005 775 14065 825
rect -50 755 14065 775
rect -50 595 12795 685
rect 12685 525 12795 595
rect -50 435 12795 525
rect 12685 365 12795 435
rect -50 275 12795 365
rect 12685 205 12795 275
rect -50 115 12795 205
rect 12685 45 12795 115
rect -50 25 14155 45
rect -50 -25 310 25
rect 360 -25 1660 25
rect 1710 -25 2995 25
rect 3045 -25 4335 25
rect 4385 -25 5675 25
rect 5725 -25 7010 25
rect 7060 -25 8350 25
rect 8400 -25 9685 25
rect 9735 -25 11025 25
rect 11075 -25 12460 25
rect 12510 -25 14155 25
rect -50 -45 14155 -25
<< labels >>
flabel nwell 365 855 365 855 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 65 2375 65 2375 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 75 -25 75 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 1425 -25 1425 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 2775 -25 2775 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 4125 -25 4125 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 5475 -25 5475 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 6825 -25 6825 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 8175 -25 8175 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 9525 -25 9525 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 10875 -25 10875 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 12225 -25 12225 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel nwell 1715 810 1715 810 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 1415 2215 1415 2215 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 2765 2055 2765 2055 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 4115 1895 4115 1895 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 5465 1735 5465 1735 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 6815 1575 6815 1575 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 8165 1415 8165 1415 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 9515 1255 9515 1255 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 10865 1095 10865 1095 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 12215 935 12215 935 2 FreeSans 400 0 0 0 vdd
port 11 ne
rlabel space 1390 690 1490 810 1 help
rlabel space 1390 690 1490 810 1 -h
flabel metal1 s 1425 720 1425 720 2 FreeSans 400 0 0 0 a1
port 1 ne
flabel metal1 s 1625 680 1625 680 2 FreeSans 400 0 0 0 z1
port 14 ne
flabel metal1 s 11075 380 11075 380 2 FreeSans 400 0 0 0 z8
port 22 ne
flabel metal1 s 10875 420 10875 420 2 FreeSans 400 0 0 0 a8
port 9 ne
flabel nwell 11165 510 11165 510 2 FreeSans 400 0 0 0 vdd
flabel nwell 9815 555 9815 555 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 9525 465 9525 465 2 FreeSans 400 0 0 0 a7
port 8 ne
flabel metal1 s 9725 425 9725 425 2 FreeSans 400 0 0 0 z7
port 21 ne
flabel nwell 5765 685 5765 685 2 FreeSans 400 0 0 0 vdd
flabel nwell 7115 640 7115 640 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 5475 595 5475 595 2 FreeSans 400 0 0 0 a4
port 5 ne
flabel metal1 s 5675 555 5675 555 2 FreeSans 400 0 0 0 z4
port 18 ne
flabel metal1 s 6825 550 6825 550 2 FreeSans 400 0 0 0 a5
port 6 ne
flabel metal1 s 7025 510 7025 510 2 FreeSans 400 0 0 0 z5
port 19 ne
flabel nwell 3065 770 3065 770 2 FreeSans 400 0 0 0 vdd
flabel nwell 4415 725 4415 725 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 2775 680 2775 680 2 FreeSans 400 0 0 0 a2
port 3 ne
flabel metal1 s 2975 640 2975 640 2 FreeSans 400 0 0 0 z2
port 16 ne
flabel metal1 s 4125 635 4125 635 2 FreeSans 400 0 0 0 a3
port 4 ne
flabel metal1 s 4325 595 4325 595 2 FreeSans 400 0 0 0 z3
port 17 ne
flabel metal1 s 8375 470 8375 470 2 FreeSans 400 0 0 0 z6
port 20 ne
flabel metal1 s 8175 510 8175 510 2 FreeSans 400 0 0 0 a6
port 7 ne
flabel nwell 8465 600 8465 600 2 FreeSans 400 0 0 0 vdd
flabel nwell 12515 465 12515 465 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 12225 375 12225 375 2 FreeSans 400 0 0 0 a9
port 10 ne
flabel metal1 s 12425 335 12425 335 2 FreeSans 400 0 0 0 z9
port 23 ne
flabel metal1 s 13725 -25 13725 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 13715 775 13715 775 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel nwell 14015 420 14015 420 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 13725 330 13725 330 2 FreeSans 400 0 0 0 a10
port 2 ne
flabel metal1 s 13925 290 13925 290 2 FreeSans 400 0 0 0 z10
port 15 ne
flabel metal1 s 75 765 75 765 2 FreeSans 400 0 0 0 a0
port 0 ne
flabel metal1 s 275 725 275 725 2 FreeSans 400 0 0 0 z0
port 13 ne
<< end >>
