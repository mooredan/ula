../../lef/amic5n_tech.lef