magic
tech scmos
timestamp 1593830479
<< metal1 >>
rect 74 11 268 25
<< metal2 >>
rect 511 25 551 96
rect 74 11 662 25
<< gv1 >>
rect 75 22 77 24
rect 80 22 82 24
rect 85 22 87 24
rect 90 22 92 24
rect 95 22 97 24
rect 100 22 102 24
rect 105 22 107 24
rect 110 22 112 24
rect 115 22 117 24
rect 120 22 122 24
rect 125 22 127 24
rect 130 22 132 24
rect 135 22 137 24
rect 140 22 142 24
rect 145 22 147 24
rect 150 22 152 24
rect 155 22 157 24
rect 160 22 162 24
rect 165 22 167 24
rect 170 22 172 24
rect 175 22 177 24
rect 180 22 182 24
rect 185 22 187 24
rect 190 22 192 24
rect 195 22 197 24
rect 200 22 202 24
rect 205 22 207 24
rect 210 22 212 24
rect 215 22 217 24
rect 220 22 222 24
rect 225 22 227 24
rect 230 22 232 24
rect 235 22 237 24
rect 240 22 242 24
rect 245 22 247 24
rect 250 22 252 24
rect 255 22 257 24
rect 260 22 262 24
rect 265 22 267 24
rect 75 17 77 19
rect 80 17 82 19
rect 85 17 87 19
rect 90 17 92 19
rect 95 17 97 19
rect 100 17 102 19
rect 105 17 107 19
rect 110 17 112 19
rect 115 17 117 19
rect 120 17 122 19
rect 125 17 127 19
rect 130 17 132 19
rect 135 17 137 19
rect 140 17 142 19
rect 145 17 147 19
rect 150 17 152 19
rect 155 17 157 19
rect 160 17 162 19
rect 165 17 167 19
rect 170 17 172 19
rect 175 17 177 19
rect 180 17 182 19
rect 185 17 187 19
rect 190 17 192 19
rect 195 17 197 19
rect 200 17 202 19
rect 205 17 207 19
rect 210 17 212 19
rect 215 17 217 19
rect 220 17 222 19
rect 225 17 227 19
rect 230 17 232 19
rect 235 17 237 19
rect 240 17 242 19
rect 245 17 247 19
rect 250 17 252 19
rect 255 17 257 19
rect 260 17 262 19
rect 265 17 267 19
rect 75 12 77 14
rect 80 12 82 14
rect 85 12 87 14
rect 90 12 92 14
rect 95 12 97 14
rect 100 12 102 14
rect 105 12 107 14
rect 110 12 112 14
rect 115 12 117 14
rect 120 12 122 14
rect 125 12 127 14
rect 130 12 132 14
rect 135 12 137 14
rect 140 12 142 14
rect 145 12 147 14
rect 150 12 152 14
rect 155 12 157 14
rect 160 12 162 14
rect 165 12 167 14
rect 170 12 172 14
rect 175 12 177 14
rect 180 12 182 14
rect 185 12 187 14
rect 190 12 192 14
rect 195 12 197 14
rect 200 12 202 14
rect 205 12 207 14
rect 210 12 212 14
rect 215 12 217 14
rect 220 12 222 14
rect 225 12 227 14
rect 230 12 232 14
rect 235 12 237 14
rect 240 12 242 14
rect 245 12 247 14
rect 250 12 252 14
rect 255 12 257 14
rect 260 12 262 14
rect 265 12 267 14
<< metal3 >>
rect 149 869 172 888
rect 469 876 492 895
use pad_in_top  pad_in_top_0
timestamp 1593798130
transform 1 0 -11 0 1 -12
box -3 -2 363 1037
use pad_x0_top  pad_x0_top_0
timestamp 1593808045
transform 1 0 349 0 1 -12
box -3 -2 363 1037
<< labels >>
rlabel metal3 s 478 885 478 885 2 x0
port 1 ne
rlabel metal3 s 156 879 156 879 2 x1
port 2 ne
rlabel metal2 s 445 16 445 16 2 n1
rlabel metal3 s 407 34 407 34 2 vdd
port 3 ne
rlabel metal3 s 377 33 377 33 2 vss
port 4 ne
<< end >>
