magic
tech amic5n
timestamp 1624143956
<< nwell >>
rect -130 550 1180 1495
<< ntransistor >>
rect 165 275 225 400
rect 375 95 435 400
rect 615 95 675 400
rect 825 275 885 400
<< ptransistor >>
rect 165 700 225 885
rect 375 700 435 1345
rect 615 700 675 1345
rect 825 700 885 885
<< nselect >>
rect 140 1115 255 1345
rect -10 0 1060 430
<< pselect >>
rect -10 1345 1060 1440
rect -10 1115 140 1345
rect 255 1115 1060 1345
rect -10 670 1060 1115
<< ndiffusion >>
rect 45 370 165 400
rect 45 320 75 370
rect 125 320 165 370
rect 45 275 165 320
rect 225 355 375 400
rect 225 305 285 355
rect 335 305 375 355
rect 225 275 375 305
rect 255 175 375 275
rect 255 125 285 175
rect 335 125 375 175
rect 255 95 375 125
rect 435 95 615 400
rect 675 345 825 400
rect 675 295 715 345
rect 765 295 825 345
rect 675 275 825 295
rect 885 370 1005 400
rect 885 320 925 370
rect 975 320 1005 370
rect 885 275 1005 320
rect 675 175 795 275
rect 675 125 715 175
rect 765 125 795 175
rect 675 95 795 125
<< pdiffusion >>
rect 255 1315 375 1345
rect 255 1265 285 1315
rect 335 1265 375 1315
rect 255 1200 375 1265
rect 255 1150 285 1200
rect 335 1150 375 1200
rect 255 1075 375 1150
rect 255 1025 285 1075
rect 335 1025 375 1075
rect 255 945 375 1025
rect 255 895 285 945
rect 335 895 375 945
rect 255 885 375 895
rect 45 815 165 885
rect 45 765 75 815
rect 125 765 165 815
rect 45 700 165 765
rect 225 825 375 885
rect 225 775 285 825
rect 335 775 375 825
rect 225 700 375 775
rect 435 1315 615 1345
rect 435 1265 500 1315
rect 550 1265 615 1315
rect 435 1180 615 1265
rect 435 1130 500 1180
rect 550 1130 615 1180
rect 435 1080 615 1130
rect 435 1030 500 1080
rect 550 1030 615 1080
rect 435 980 615 1030
rect 435 930 500 980
rect 550 930 615 980
rect 435 880 615 930
rect 435 830 500 880
rect 550 830 615 880
rect 435 780 615 830
rect 435 730 500 780
rect 550 730 615 780
rect 435 700 615 730
rect 675 1315 795 1345
rect 675 1265 715 1315
rect 765 1265 795 1315
rect 675 1200 795 1265
rect 675 1150 715 1200
rect 765 1150 795 1200
rect 675 1075 795 1150
rect 675 1025 715 1075
rect 765 1025 795 1075
rect 675 945 795 1025
rect 675 895 715 945
rect 765 895 795 945
rect 675 885 795 895
rect 675 825 825 885
rect 675 775 715 825
rect 765 775 825 825
rect 675 700 825 775
rect 885 815 1005 885
rect 885 765 925 815
rect 975 765 1005 815
rect 885 700 1005 765
<< nsubstratendiff >>
rect 140 1315 255 1345
rect 140 1265 170 1315
rect 220 1265 255 1315
rect 140 1195 255 1265
rect 140 1145 170 1195
rect 220 1145 255 1195
rect 140 1115 255 1145
<< nsubstratencontact >>
rect 170 1265 220 1315
rect 170 1145 220 1195
<< ndcontact >>
rect 75 320 125 370
rect 285 305 335 355
rect 285 125 335 175
rect 715 295 765 345
rect 925 320 975 370
rect 715 125 765 175
<< pdcontact >>
rect 285 1265 335 1315
rect 285 1150 335 1200
rect 285 1025 335 1075
rect 285 895 335 945
rect 75 765 125 815
rect 285 775 335 825
rect 500 1265 550 1315
rect 500 1130 550 1180
rect 500 1030 550 1080
rect 500 930 550 980
rect 500 830 550 880
rect 500 730 550 780
rect 715 1265 765 1315
rect 715 1150 765 1200
rect 715 1025 765 1075
rect 715 895 765 945
rect 715 775 765 825
rect 925 765 975 815
<< polysilicon >>
rect 375 1345 435 1410
rect 615 1345 675 1410
rect 165 885 225 950
rect 825 1145 940 1165
rect 825 1095 870 1145
rect 920 1095 940 1145
rect 825 1075 940 1095
rect 825 885 885 1075
rect 165 400 225 700
rect 375 525 435 700
rect 325 505 435 525
rect 325 455 345 505
rect 395 455 435 505
rect 325 435 435 455
rect 375 400 435 435
rect 615 525 675 700
rect 615 505 745 525
rect 615 455 675 505
rect 725 455 745 505
rect 615 435 745 455
rect 615 400 675 435
rect 825 400 885 700
rect 165 205 225 275
rect 55 185 225 205
rect 55 135 75 185
rect 125 135 225 185
rect 55 115 225 135
rect 825 210 885 275
rect 375 30 435 95
rect 615 30 675 95
<< polycontact >>
rect 870 1095 920 1145
rect 345 455 395 505
rect 675 455 725 505
rect 75 135 125 185
<< metal1 >>
rect 0 1395 1050 1485
rect 150 1315 355 1395
rect 150 1265 170 1315
rect 220 1265 285 1315
rect 335 1265 355 1315
rect 150 1200 355 1265
rect 150 1195 285 1200
rect 150 1145 170 1195
rect 220 1150 285 1195
rect 335 1150 355 1200
rect 220 1145 355 1150
rect 150 1125 355 1145
rect 265 1075 355 1125
rect 265 1025 285 1075
rect 335 1025 355 1075
rect 265 945 355 1025
rect 265 895 285 945
rect 335 895 355 945
rect 55 815 145 845
rect 55 765 75 815
rect 125 765 145 815
rect 55 525 145 765
rect 265 825 355 895
rect 265 775 285 825
rect 335 775 355 825
rect 265 745 355 775
rect 480 1315 570 1335
rect 480 1265 500 1315
rect 550 1265 570 1315
rect 480 1180 570 1265
rect 480 1130 500 1180
rect 550 1130 570 1180
rect 480 1080 570 1130
rect 480 1030 500 1080
rect 550 1030 570 1080
rect 480 980 570 1030
rect 480 930 500 980
rect 550 930 570 980
rect 480 880 570 930
rect 480 830 500 880
rect 550 830 570 880
rect 480 780 570 830
rect 480 730 500 780
rect 550 730 570 780
rect 695 1315 785 1395
rect 695 1265 715 1315
rect 765 1265 785 1315
rect 695 1200 785 1265
rect 695 1150 715 1200
rect 765 1150 785 1200
rect 695 1075 785 1150
rect 850 1145 1020 1165
rect 850 1095 870 1145
rect 920 1095 1020 1145
rect 850 1075 1020 1095
rect 695 1025 715 1075
rect 765 1025 785 1075
rect 695 945 785 1025
rect 695 895 715 945
rect 765 895 785 945
rect 695 825 785 895
rect 695 775 715 825
rect 765 775 785 825
rect 695 745 785 775
rect 905 815 995 845
rect 905 765 925 815
rect 975 765 995 815
rect 55 505 415 525
rect 55 455 345 505
rect 395 455 415 505
rect 55 435 415 455
rect 55 370 145 435
rect 480 375 570 730
rect 905 525 995 765
rect 655 505 995 525
rect 655 455 675 505
rect 725 455 995 505
rect 655 435 995 455
rect 55 320 75 370
rect 125 320 145 370
rect 55 300 145 320
rect 265 355 355 375
rect 265 305 285 355
rect 335 305 355 355
rect 30 185 145 205
rect 30 135 75 185
rect 125 135 145 185
rect 30 115 145 135
rect 265 175 355 305
rect 480 345 785 375
rect 480 295 715 345
rect 765 295 785 345
rect 480 275 785 295
rect 905 370 995 435
rect 905 320 925 370
rect 975 320 995 370
rect 905 285 995 320
rect 265 125 285 175
rect 335 125 355 175
rect 265 45 355 125
rect 695 175 785 275
rect 695 125 715 175
rect 765 125 785 175
rect 695 45 785 125
rect 0 -45 1050 45
<< labels >>
flabel metal1 s 245 1415 245 1415 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 510 470 510 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel nwell 230 600 230 600 8 FreeSans 400 180 0 0 vdd
flabel metal1 s 70 130 70 130 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 865 1085 865 1085 2 FreeSans 400 0 0 0 b
port 2 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 4 ne
<< end >>
