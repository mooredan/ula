* clamp2 normal power up testing
*
.lib device_models/AMI_C5N.lib TT
.include "clamp2.cir"

* Power
Vvdd vsrc 0 DC 0 PWL ( 0 0 1u 0 4u 5)
Rsrc vsrc vdd 0.010

* Ground
Vvss vss 0 DC 0

* Clamp(s)
XCLAMP  vdd vss clamp2
XCLAMP1 vdd vss clamp2
* XCLAMP2 vdd vss clamp2
* XCLAMP3 vdd vss clamp2


* DUT load
CDUT vdd vss 10p
RDUT vdd vss 10Meg


.save all
.tran 1n 10.0u 

.control
destroy all
run
plot v(vdd)
plot i(vvss)
plot v(xclamp.trig) v(xclamp.ntrig)


.endc
.end
