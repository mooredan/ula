magic
tech scmos
magscale 1 2
timestamp 1570494029
<< error_p >>
rect 1584 1322 1586 1324
rect 1582 1320 1584 1322
rect 1574 1312 1576 1314
rect 1572 1310 1574 1312
rect 1564 1302 1566 1304
rect 1562 1300 1564 1302
rect 1554 1292 1556 1294
rect 1552 1290 1554 1292
rect 1544 1282 1546 1284
rect 1542 1280 1544 1282
rect 1534 1272 1536 1274
rect 1532 1270 1534 1272
rect 1524 1262 1526 1264
rect 1522 1260 1524 1262
rect 1514 1252 1516 1254
rect 1512 1250 1514 1252
rect 1504 1242 1506 1244
rect 1502 1240 1504 1242
rect 1494 1232 1496 1234
rect 1492 1230 1494 1232
rect 1484 1222 1486 1224
rect 1482 1220 1484 1222
rect 1474 1212 1476 1214
rect 1472 1210 1474 1212
rect 1464 1202 1466 1204
rect 1462 1200 1464 1202
rect 1454 1192 1456 1194
rect 1452 1190 1454 1192
rect 1444 1182 1446 1184
rect 1442 1180 1444 1182
rect 1434 1172 1436 1174
rect 1432 1170 1434 1172
rect 1424 1162 1426 1164
rect 1422 1160 1424 1162
rect 1414 1152 1416 1154
rect 1412 1150 1414 1152
rect 1404 1142 1406 1144
rect 1402 1140 1404 1142
rect 1394 1132 1396 1134
rect 1392 1130 1394 1132
rect 1384 1122 1386 1124
rect 1382 1120 1384 1122
rect 1374 1112 1376 1114
rect 1372 1110 1374 1112
rect 1364 1102 1366 1104
rect 1362 1100 1364 1102
rect 1354 1092 1356 1094
rect 1352 1090 1354 1092
rect 1344 1082 1346 1084
rect 1342 1080 1344 1082
rect 1334 1072 1336 1074
rect 1332 1070 1334 1072
rect 1324 1062 1326 1064
rect 1322 1060 1324 1062
rect 1572 1054 1574 1056
rect 1592 1054 1594 1056
rect 1314 1052 1316 1054
rect 1570 1052 1572 1054
rect 1594 1052 1596 1054
rect 1312 1050 1314 1052
rect 1562 1044 1564 1046
rect 1304 1042 1306 1044
rect 1560 1042 1562 1044
rect 1302 1040 1304 1042
rect 1552 1034 1554 1036
rect 1294 1032 1296 1034
rect 1550 1032 1552 1034
rect 1292 1030 1294 1032
rect 1542 1024 1544 1026
rect 1284 1022 1286 1024
rect 1540 1022 1542 1024
rect 1594 1022 1596 1024
rect 1282 1020 1284 1022
rect 1592 1020 1594 1022
rect 1532 1014 1534 1016
rect 1274 1012 1276 1014
rect 1530 1012 1532 1014
rect 1584 1012 1586 1014
rect 1272 1010 1274 1012
rect 1582 1010 1584 1012
rect 1522 1004 1524 1006
rect 1264 1002 1266 1004
rect 1520 1002 1522 1004
rect 1574 1002 1576 1004
rect 1262 1000 1264 1002
rect 1572 1000 1574 1002
rect 1512 994 1514 996
rect 1254 992 1256 994
rect 1510 992 1512 994
rect 1564 992 1566 994
rect 1252 990 1254 992
rect 1562 990 1564 992
rect 1502 984 1504 986
rect 1244 982 1246 984
rect 1500 982 1502 984
rect 1554 982 1556 984
rect 1242 980 1244 982
rect 1552 980 1554 982
rect 1492 974 1494 976
rect 1234 972 1236 974
rect 1490 972 1492 974
rect 1544 972 1546 974
rect 1232 970 1234 972
rect 1542 970 1544 972
rect 1482 964 1484 966
rect 1224 962 1226 964
rect 1480 962 1482 964
rect 1534 962 1536 964
rect 1222 960 1224 962
rect 1532 960 1534 962
rect 1472 954 1474 956
rect 1214 952 1216 954
rect 1470 952 1472 954
rect 1524 952 1526 954
rect 1212 950 1214 952
rect 1522 950 1524 952
rect 1462 944 1464 946
rect 1204 942 1206 944
rect 1460 942 1462 944
rect 1514 942 1516 944
rect 1202 940 1204 942
rect 1512 940 1514 942
rect 1452 934 1454 936
rect 1194 932 1196 934
rect 1450 932 1452 934
rect 1504 932 1506 934
rect 1192 930 1194 932
rect 1502 930 1504 932
rect 1442 924 1444 926
rect 1184 922 1186 924
rect 1440 922 1442 924
rect 1494 922 1496 924
rect 1182 920 1184 922
rect 1492 920 1494 922
rect 1432 914 1434 916
rect 1174 912 1176 914
rect 1430 912 1432 914
rect 1484 912 1486 914
rect 1172 910 1174 912
rect 1482 910 1484 912
rect 1422 904 1424 906
rect 1164 902 1166 904
rect 1420 902 1422 904
rect 1474 902 1476 904
rect 1162 900 1164 902
rect 1472 900 1474 902
rect 1412 894 1414 896
rect 1154 892 1156 894
rect 1410 892 1412 894
rect 1464 892 1466 894
rect 1152 890 1154 892
rect 1462 890 1464 892
rect 1402 884 1404 886
rect 1702 884 1704 886
rect 1732 884 1734 886
rect 1144 882 1146 884
rect 1400 882 1402 884
rect 1454 882 1456 884
rect 1700 882 1702 884
rect 1734 882 1736 884
rect 1142 880 1144 882
rect 1452 880 1454 882
rect 1392 874 1394 876
rect 1692 874 1694 876
rect 1134 872 1136 874
rect 1390 872 1392 874
rect 1444 872 1446 874
rect 1690 872 1692 874
rect 1132 870 1134 872
rect 1442 870 1444 872
rect 1382 864 1384 866
rect 1682 864 1684 866
rect 1124 862 1126 864
rect 1380 862 1382 864
rect 1434 862 1436 864
rect 1680 862 1682 864
rect 1734 862 1736 864
rect 1122 860 1124 862
rect 1432 860 1434 862
rect 1732 860 1734 862
rect 1372 854 1374 856
rect 1672 854 1674 856
rect 1114 852 1116 854
rect 1370 852 1372 854
rect 1424 852 1426 854
rect 1670 852 1672 854
rect 1724 852 1726 854
rect 1112 850 1114 852
rect 1422 850 1424 852
rect 1722 850 1724 852
rect 1362 844 1364 846
rect 1662 844 1664 846
rect 1722 844 1724 846
rect 1732 844 1734 846
rect 1752 844 1754 846
rect 1762 844 1764 846
rect 1782 844 1784 846
rect 1792 844 1794 846
rect 1812 844 1814 846
rect 1822 844 1824 846
rect 1842 844 1844 846
rect 1852 844 1854 846
rect 1872 844 1874 846
rect 1882 844 1884 846
rect 1902 844 1904 846
rect 1912 844 1914 846
rect 1932 844 1934 846
rect 1942 844 1944 846
rect 1962 844 1964 846
rect 1972 844 1974 846
rect 1104 842 1106 844
rect 1360 842 1362 844
rect 1414 842 1416 844
rect 1660 842 1662 844
rect 1714 842 1716 844
rect 1720 842 1722 844
rect 1734 842 1736 844
rect 1750 842 1752 844
rect 1764 842 1766 844
rect 1780 842 1782 844
rect 1794 842 1796 844
rect 1810 842 1812 844
rect 1824 842 1826 844
rect 1840 842 1842 844
rect 1854 842 1856 844
rect 1870 842 1872 844
rect 1884 842 1886 844
rect 1900 842 1902 844
rect 1914 842 1916 844
rect 1930 842 1932 844
rect 1944 842 1946 844
rect 1960 842 1962 844
rect 1974 842 1976 844
rect 1102 840 1104 842
rect 1412 840 1414 842
rect 1712 840 1714 842
rect 1352 834 1354 836
rect 1652 834 1654 836
rect 1742 834 1744 836
rect 1772 834 1774 836
rect 1802 834 1804 836
rect 1832 834 1834 836
rect 1862 834 1864 836
rect 1892 834 1894 836
rect 1922 834 1924 836
rect 1952 834 1954 836
rect 1982 834 1984 836
rect 1094 832 1096 834
rect 1350 832 1352 834
rect 1404 832 1406 834
rect 1650 832 1652 834
rect 1704 832 1706 834
rect 1720 832 1722 834
rect 1744 832 1746 834
rect 1750 832 1752 834
rect 1774 832 1776 834
rect 1780 832 1782 834
rect 1804 832 1806 834
rect 1810 832 1812 834
rect 1834 832 1836 834
rect 1840 832 1842 834
rect 1864 832 1866 834
rect 1870 832 1872 834
rect 1894 832 1896 834
rect 1900 832 1902 834
rect 1924 832 1926 834
rect 1930 832 1932 834
rect 1954 832 1956 834
rect 1960 832 1962 834
rect 1984 832 1986 834
rect 1092 830 1094 832
rect 1402 830 1404 832
rect 1702 830 1704 832
rect 1722 830 1724 832
rect 1752 830 1754 832
rect 1782 830 1784 832
rect 1812 830 1814 832
rect 1842 830 1844 832
rect 1872 830 1874 832
rect 1902 830 1904 832
rect 1932 830 1934 832
rect 1962 830 1964 832
rect 1342 824 1344 826
rect 1642 824 1644 826
rect 1722 824 1724 826
rect 1752 824 1754 826
rect 1782 824 1784 826
rect 1812 824 1814 826
rect 1842 824 1844 826
rect 1872 824 1874 826
rect 1902 824 1904 826
rect 1932 824 1934 826
rect 1962 824 1964 826
rect 1084 822 1086 824
rect 1340 822 1342 824
rect 1394 822 1396 824
rect 1640 822 1642 824
rect 1694 822 1696 824
rect 1720 822 1722 824
rect 1744 822 1746 824
rect 1750 822 1752 824
rect 1774 822 1776 824
rect 1780 822 1782 824
rect 1804 822 1806 824
rect 1810 822 1812 824
rect 1834 822 1836 824
rect 1840 822 1842 824
rect 1864 822 1866 824
rect 1870 822 1872 824
rect 1894 822 1896 824
rect 1900 822 1902 824
rect 1924 822 1926 824
rect 1930 822 1932 824
rect 1954 822 1956 824
rect 1960 822 1962 824
rect 1984 822 1986 824
rect 1082 820 1084 822
rect 1392 820 1394 822
rect 1692 820 1694 822
rect 1742 820 1744 822
rect 1772 820 1774 822
rect 1802 820 1804 822
rect 1832 820 1834 822
rect 1862 820 1864 822
rect 1892 820 1894 822
rect 1922 820 1924 822
rect 1952 820 1954 822
rect 1982 820 1984 822
rect 1332 814 1334 816
rect 1632 814 1634 816
rect 1692 814 1694 816
rect 1702 814 1704 816
rect 1742 814 1744 816
rect 1772 814 1774 816
rect 1802 814 1804 816
rect 1832 814 1834 816
rect 1862 814 1864 816
rect 1892 814 1894 816
rect 1922 814 1924 816
rect 1952 814 1954 816
rect 1982 814 1984 816
rect 1074 812 1076 814
rect 1330 812 1332 814
rect 1384 812 1386 814
rect 1630 812 1632 814
rect 1684 812 1686 814
rect 1690 812 1692 814
rect 1704 812 1706 814
rect 1720 812 1722 814
rect 1744 812 1746 814
rect 1750 812 1752 814
rect 1774 812 1776 814
rect 1780 812 1782 814
rect 1804 812 1806 814
rect 1810 812 1812 814
rect 1834 812 1836 814
rect 1840 812 1842 814
rect 1864 812 1866 814
rect 1870 812 1872 814
rect 1894 812 1896 814
rect 1900 812 1902 814
rect 1924 812 1926 814
rect 1930 812 1932 814
rect 1954 812 1956 814
rect 1960 812 1962 814
rect 1984 812 1986 814
rect 1072 810 1074 812
rect 1382 810 1384 812
rect 1682 810 1684 812
rect 1722 810 1724 812
rect 1752 810 1754 812
rect 1782 810 1784 812
rect 1812 810 1814 812
rect 1842 810 1844 812
rect 1872 810 1874 812
rect 1902 810 1904 812
rect 1932 810 1934 812
rect 1962 810 1964 812
rect 1322 804 1324 806
rect 1622 804 1624 806
rect 1682 804 1684 806
rect 1722 804 1724 806
rect 1752 804 1754 806
rect 1782 804 1784 806
rect 1812 804 1814 806
rect 1842 804 1844 806
rect 1872 804 1874 806
rect 1902 804 1904 806
rect 1932 804 1934 806
rect 1962 804 1964 806
rect 1064 802 1066 804
rect 1320 802 1322 804
rect 1374 802 1376 804
rect 1620 802 1622 804
rect 1674 802 1676 804
rect 1680 802 1682 804
rect 1704 802 1706 804
rect 1720 802 1722 804
rect 1744 802 1746 804
rect 1750 802 1752 804
rect 1774 802 1776 804
rect 1780 802 1782 804
rect 1804 802 1806 804
rect 1810 802 1812 804
rect 1834 802 1836 804
rect 1840 802 1842 804
rect 1864 802 1866 804
rect 1870 802 1872 804
rect 1894 802 1896 804
rect 1900 802 1902 804
rect 1924 802 1926 804
rect 1930 802 1932 804
rect 1954 802 1956 804
rect 1960 802 1962 804
rect 1984 802 1986 804
rect 1062 800 1064 802
rect 1372 800 1374 802
rect 1672 800 1674 802
rect 1702 800 1704 802
rect 1742 800 1744 802
rect 1772 800 1774 802
rect 1802 800 1804 802
rect 1832 800 1834 802
rect 1862 800 1864 802
rect 1892 800 1894 802
rect 1922 800 1924 802
rect 1952 800 1954 802
rect 1982 800 1984 802
rect 1312 794 1314 796
rect 1612 794 1614 796
rect 1672 794 1674 796
rect 1702 794 1704 796
rect 1742 794 1744 796
rect 1772 794 1774 796
rect 1802 794 1804 796
rect 1832 794 1834 796
rect 1862 794 1864 796
rect 1892 794 1894 796
rect 1922 794 1924 796
rect 1952 794 1954 796
rect 1982 794 1984 796
rect 1054 792 1056 794
rect 1310 792 1312 794
rect 1364 792 1366 794
rect 1610 792 1612 794
rect 1664 792 1666 794
rect 1670 792 1672 794
rect 1704 792 1706 794
rect 1720 792 1722 794
rect 1744 792 1746 794
rect 1750 792 1752 794
rect 1774 792 1776 794
rect 1780 792 1782 794
rect 1804 792 1806 794
rect 1810 792 1812 794
rect 1834 792 1836 794
rect 1840 792 1842 794
rect 1864 792 1866 794
rect 1870 792 1872 794
rect 1894 792 1896 794
rect 1900 792 1902 794
rect 1924 792 1926 794
rect 1930 792 1932 794
rect 1954 792 1956 794
rect 1960 792 1962 794
rect 1984 792 1986 794
rect 1052 790 1054 792
rect 1362 790 1364 792
rect 1662 790 1664 792
rect 1722 790 1724 792
rect 1752 790 1754 792
rect 1782 790 1784 792
rect 1812 790 1814 792
rect 1842 790 1844 792
rect 1872 790 1874 792
rect 1902 790 1904 792
rect 1932 790 1934 792
rect 1962 790 1964 792
rect 1302 784 1304 786
rect 1602 784 1604 786
rect 1662 784 1664 786
rect 1722 784 1724 786
rect 1752 784 1754 786
rect 1782 784 1784 786
rect 1812 784 1814 786
rect 1842 784 1844 786
rect 1872 784 1874 786
rect 1902 784 1904 786
rect 1932 784 1934 786
rect 1962 784 1964 786
rect 1044 782 1046 784
rect 1300 782 1302 784
rect 1354 782 1356 784
rect 1600 782 1602 784
rect 1654 782 1656 784
rect 1660 782 1662 784
rect 1704 782 1706 784
rect 1720 782 1722 784
rect 1744 782 1746 784
rect 1750 782 1752 784
rect 1774 782 1776 784
rect 1780 782 1782 784
rect 1804 782 1806 784
rect 1810 782 1812 784
rect 1834 782 1836 784
rect 1840 782 1842 784
rect 1864 782 1866 784
rect 1870 782 1872 784
rect 1894 782 1896 784
rect 1900 782 1902 784
rect 1924 782 1926 784
rect 1930 782 1932 784
rect 1954 782 1956 784
rect 1960 782 1962 784
rect 1984 782 1986 784
rect 1042 780 1044 782
rect 1352 780 1354 782
rect 1652 780 1654 782
rect 1702 780 1704 782
rect 1742 780 1744 782
rect 1772 780 1774 782
rect 1802 780 1804 782
rect 1832 780 1834 782
rect 1862 780 1864 782
rect 1892 780 1894 782
rect 1922 780 1924 782
rect 1952 780 1954 782
rect 1982 780 1984 782
rect 1292 774 1294 776
rect 1592 774 1594 776
rect 1652 774 1654 776
rect 1742 774 1744 776
rect 1772 774 1774 776
rect 1802 774 1804 776
rect 1832 774 1834 776
rect 1862 774 1864 776
rect 1892 774 1894 776
rect 1922 774 1924 776
rect 1952 774 1954 776
rect 1982 774 1984 776
rect 1034 772 1036 774
rect 1290 772 1292 774
rect 1344 772 1346 774
rect 1590 772 1592 774
rect 1644 772 1646 774
rect 1650 772 1652 774
rect 1694 772 1696 774
rect 1720 772 1722 774
rect 1744 772 1746 774
rect 1750 772 1752 774
rect 1774 772 1776 774
rect 1780 772 1782 774
rect 1804 772 1806 774
rect 1810 772 1812 774
rect 1834 772 1836 774
rect 1840 772 1842 774
rect 1864 772 1866 774
rect 1870 772 1872 774
rect 1894 772 1896 774
rect 1900 772 1902 774
rect 1924 772 1926 774
rect 1930 772 1932 774
rect 1954 772 1956 774
rect 1960 772 1962 774
rect 1984 772 1986 774
rect 1032 770 1034 772
rect 1342 770 1344 772
rect 1642 770 1644 772
rect 1692 770 1694 772
rect 1722 770 1724 772
rect 1752 770 1754 772
rect 1782 770 1784 772
rect 1812 770 1814 772
rect 1842 770 1844 772
rect 1872 770 1874 772
rect 1902 770 1904 772
rect 1932 770 1934 772
rect 1962 770 1964 772
rect 1282 764 1284 766
rect 1582 764 1584 766
rect 1642 764 1644 766
rect 1692 764 1694 766
rect 1702 764 1704 766
rect 1722 764 1724 766
rect 1752 764 1754 766
rect 1782 764 1784 766
rect 1812 764 1814 766
rect 1842 764 1844 766
rect 1872 764 1874 766
rect 1902 764 1904 766
rect 1932 764 1934 766
rect 1962 764 1964 766
rect 1024 762 1026 764
rect 1280 762 1282 764
rect 1334 762 1336 764
rect 1580 762 1582 764
rect 1634 762 1636 764
rect 1640 762 1642 764
rect 1684 762 1686 764
rect 1690 762 1692 764
rect 1704 762 1706 764
rect 1720 762 1722 764
rect 1744 762 1746 764
rect 1750 762 1752 764
rect 1774 762 1776 764
rect 1780 762 1782 764
rect 1804 762 1806 764
rect 1810 762 1812 764
rect 1834 762 1836 764
rect 1840 762 1842 764
rect 1864 762 1866 764
rect 1870 762 1872 764
rect 1894 762 1896 764
rect 1900 762 1902 764
rect 1924 762 1926 764
rect 1930 762 1932 764
rect 1954 762 1956 764
rect 1960 762 1962 764
rect 1984 762 1986 764
rect 1022 760 1024 762
rect 1332 760 1334 762
rect 1632 760 1634 762
rect 1682 760 1684 762
rect 1742 760 1744 762
rect 1772 760 1774 762
rect 1802 760 1804 762
rect 1832 760 1834 762
rect 1862 760 1864 762
rect 1892 760 1894 762
rect 1922 760 1924 762
rect 1952 760 1954 762
rect 1982 760 1984 762
rect 1272 754 1274 756
rect 1572 754 1574 756
rect 1632 754 1634 756
rect 1682 754 1684 756
rect 1742 754 1744 756
rect 1772 754 1774 756
rect 1802 754 1804 756
rect 1832 754 1834 756
rect 1862 754 1864 756
rect 1892 754 1894 756
rect 1922 754 1924 756
rect 1952 754 1954 756
rect 1982 754 1984 756
rect 1014 752 1016 754
rect 1270 752 1272 754
rect 1324 752 1326 754
rect 1570 752 1572 754
rect 1624 752 1626 754
rect 1630 752 1632 754
rect 1674 752 1676 754
rect 1680 752 1682 754
rect 1704 752 1706 754
rect 1720 752 1722 754
rect 1744 752 1746 754
rect 1750 752 1752 754
rect 1774 752 1776 754
rect 1780 752 1782 754
rect 1804 752 1806 754
rect 1810 752 1812 754
rect 1834 752 1836 754
rect 1840 752 1842 754
rect 1864 752 1866 754
rect 1870 752 1872 754
rect 1894 752 1896 754
rect 1900 752 1902 754
rect 1924 752 1926 754
rect 1930 752 1932 754
rect 1954 752 1956 754
rect 1960 752 1962 754
rect 1984 752 1986 754
rect 1012 750 1014 752
rect 1322 750 1324 752
rect 1622 750 1624 752
rect 1672 750 1674 752
rect 1702 750 1704 752
rect 1722 750 1724 752
rect 1752 750 1754 752
rect 1782 750 1784 752
rect 1812 750 1814 752
rect 1842 750 1844 752
rect 1872 750 1874 752
rect 1902 750 1904 752
rect 1932 750 1934 752
rect 1962 750 1964 752
rect 1262 744 1264 746
rect 1562 744 1564 746
rect 1622 744 1624 746
rect 1672 744 1674 746
rect 1722 744 1724 746
rect 1752 744 1754 746
rect 1782 744 1784 746
rect 1812 744 1814 746
rect 1842 744 1844 746
rect 1872 744 1874 746
rect 1902 744 1904 746
rect 1932 744 1934 746
rect 1962 744 1964 746
rect 1004 742 1006 744
rect 1260 742 1262 744
rect 1314 742 1316 744
rect 1560 742 1562 744
rect 1614 742 1616 744
rect 1620 742 1622 744
rect 1664 742 1666 744
rect 1670 742 1672 744
rect 1694 742 1696 744
rect 1720 742 1722 744
rect 1744 742 1746 744
rect 1750 742 1752 744
rect 1774 742 1776 744
rect 1780 742 1782 744
rect 1804 742 1806 744
rect 1810 742 1812 744
rect 1834 742 1836 744
rect 1840 742 1842 744
rect 1864 742 1866 744
rect 1870 742 1872 744
rect 1894 742 1896 744
rect 1900 742 1902 744
rect 1924 742 1926 744
rect 1930 742 1932 744
rect 1954 742 1956 744
rect 1960 742 1962 744
rect 1984 742 1986 744
rect 1002 740 1004 742
rect 1312 740 1314 742
rect 1612 740 1614 742
rect 1662 740 1664 742
rect 1692 740 1694 742
rect 1742 740 1744 742
rect 1772 740 1774 742
rect 1802 740 1804 742
rect 1832 740 1834 742
rect 1862 740 1864 742
rect 1892 740 1894 742
rect 1922 740 1924 742
rect 1952 740 1954 742
rect 1982 740 1984 742
rect 1252 734 1254 736
rect 1552 734 1554 736
rect 1612 734 1614 736
rect 1662 734 1664 736
rect 1742 734 1744 736
rect 1772 734 1774 736
rect 1802 734 1804 736
rect 1832 734 1834 736
rect 1862 734 1864 736
rect 1892 734 1894 736
rect 1922 734 1924 736
rect 1952 734 1954 736
rect 1982 734 1984 736
rect 994 732 996 734
rect 1250 732 1252 734
rect 1304 732 1306 734
rect 1550 732 1552 734
rect 1604 732 1606 734
rect 1610 732 1612 734
rect 1654 732 1656 734
rect 1660 732 1662 734
rect 1684 732 1686 734
rect 1720 732 1722 734
rect 1744 732 1746 734
rect 1750 732 1752 734
rect 1774 732 1776 734
rect 1780 732 1782 734
rect 1804 732 1806 734
rect 1810 732 1812 734
rect 1834 732 1836 734
rect 1840 732 1842 734
rect 1864 732 1866 734
rect 1870 732 1872 734
rect 1894 732 1896 734
rect 1900 732 1902 734
rect 1924 732 1926 734
rect 1930 732 1932 734
rect 1954 732 1956 734
rect 1960 732 1962 734
rect 1984 732 1986 734
rect 992 730 994 732
rect 1302 730 1304 732
rect 1602 730 1604 732
rect 1652 730 1654 732
rect 1682 730 1684 732
rect 1722 730 1724 732
rect 1752 730 1754 732
rect 1782 730 1784 732
rect 1812 730 1814 732
rect 1842 730 1844 732
rect 1872 730 1874 732
rect 1902 730 1904 732
rect 1932 730 1934 732
rect 1962 730 1964 732
rect 1242 724 1244 726
rect 1542 724 1544 726
rect 1602 724 1604 726
rect 1652 724 1654 726
rect 1722 724 1724 726
rect 1752 724 1754 726
rect 1782 724 1784 726
rect 1812 724 1814 726
rect 1842 724 1844 726
rect 1872 724 1874 726
rect 1902 724 1904 726
rect 1932 724 1934 726
rect 1962 724 1964 726
rect 984 722 986 724
rect 1240 722 1242 724
rect 1294 722 1296 724
rect 1540 722 1542 724
rect 1594 722 1596 724
rect 1600 722 1602 724
rect 1644 722 1646 724
rect 1650 722 1652 724
rect 1674 722 1676 724
rect 1720 722 1722 724
rect 1744 722 1746 724
rect 1750 722 1752 724
rect 1774 722 1776 724
rect 1780 722 1782 724
rect 1804 722 1806 724
rect 1810 722 1812 724
rect 1834 722 1836 724
rect 1840 722 1842 724
rect 1864 722 1866 724
rect 1870 722 1872 724
rect 1894 722 1896 724
rect 1900 722 1902 724
rect 1924 722 1926 724
rect 1930 722 1932 724
rect 1954 722 1956 724
rect 1960 722 1962 724
rect 1984 722 1986 724
rect 982 720 984 722
rect 1292 720 1294 722
rect 1592 720 1594 722
rect 1642 720 1644 722
rect 1672 720 1674 722
rect 1742 720 1744 722
rect 1772 720 1774 722
rect 1802 720 1804 722
rect 1832 720 1834 722
rect 1862 720 1864 722
rect 1892 720 1894 722
rect 1922 720 1924 722
rect 1952 720 1954 722
rect 1982 720 1984 722
rect 1232 714 1234 716
rect 1532 714 1534 716
rect 1592 714 1594 716
rect 1642 714 1644 716
rect 1742 714 1744 716
rect 1772 714 1774 716
rect 1802 714 1804 716
rect 1832 714 1834 716
rect 1862 714 1864 716
rect 1892 714 1894 716
rect 1922 714 1924 716
rect 1952 714 1954 716
rect 1982 714 1984 716
rect 974 712 976 714
rect 1230 712 1232 714
rect 1284 712 1286 714
rect 1530 712 1532 714
rect 1584 712 1586 714
rect 1590 712 1592 714
rect 1634 712 1636 714
rect 1640 712 1642 714
rect 1664 712 1666 714
rect 1720 712 1722 714
rect 1744 712 1746 714
rect 1750 712 1752 714
rect 1774 712 1776 714
rect 1780 712 1782 714
rect 1804 712 1806 714
rect 1810 712 1812 714
rect 1834 712 1836 714
rect 1840 712 1842 714
rect 1864 712 1866 714
rect 1870 712 1872 714
rect 1894 712 1896 714
rect 1900 712 1902 714
rect 1924 712 1926 714
rect 1930 712 1932 714
rect 1954 712 1956 714
rect 1960 712 1962 714
rect 1984 712 1986 714
rect 972 710 974 712
rect 1282 710 1284 712
rect 1582 710 1584 712
rect 1632 710 1634 712
rect 1662 710 1664 712
rect 1722 710 1724 712
rect 1752 710 1754 712
rect 1782 710 1784 712
rect 1812 710 1814 712
rect 1842 710 1844 712
rect 1872 710 1874 712
rect 1902 710 1904 712
rect 1932 710 1934 712
rect 1962 710 1964 712
rect 1222 704 1224 706
rect 1522 704 1524 706
rect 1582 704 1584 706
rect 1632 704 1634 706
rect 1692 704 1694 706
rect 1702 704 1704 706
rect 1722 704 1724 706
rect 1752 704 1754 706
rect 1782 704 1784 706
rect 1812 704 1814 706
rect 1842 704 1844 706
rect 1872 704 1874 706
rect 1902 704 1904 706
rect 1932 704 1934 706
rect 1962 704 1964 706
rect 964 702 966 704
rect 1220 702 1222 704
rect 1274 702 1276 704
rect 1520 702 1522 704
rect 1574 702 1576 704
rect 1580 702 1582 704
rect 1624 702 1626 704
rect 1630 702 1632 704
rect 1654 702 1656 704
rect 1690 702 1692 704
rect 1704 702 1706 704
rect 1720 702 1722 704
rect 1744 702 1746 704
rect 1750 702 1752 704
rect 1774 702 1776 704
rect 1780 702 1782 704
rect 1804 702 1806 704
rect 1810 702 1812 704
rect 1834 702 1836 704
rect 1840 702 1842 704
rect 1864 702 1866 704
rect 1870 702 1872 704
rect 1894 702 1896 704
rect 1900 702 1902 704
rect 1924 702 1926 704
rect 1930 702 1932 704
rect 1954 702 1956 704
rect 1960 702 1962 704
rect 1984 702 1986 704
rect 962 700 964 702
rect 1272 700 1274 702
rect 1572 700 1574 702
rect 1622 700 1624 702
rect 1652 700 1654 702
rect 1742 700 1744 702
rect 1772 700 1774 702
rect 1802 700 1804 702
rect 1832 700 1834 702
rect 1862 700 1864 702
rect 1892 700 1894 702
rect 1922 700 1924 702
rect 1952 700 1954 702
rect 1982 700 1984 702
rect 1212 694 1214 696
rect 1512 694 1514 696
rect 1572 694 1574 696
rect 1622 694 1624 696
rect 1682 694 1684 696
rect 1712 694 1714 696
rect 1742 694 1744 696
rect 1772 694 1774 696
rect 954 692 956 694
rect 1210 692 1212 694
rect 1264 692 1266 694
rect 1510 692 1512 694
rect 1564 692 1566 694
rect 1570 692 1572 694
rect 1624 692 1626 694
rect 1680 692 1682 694
rect 1714 692 1716 694
rect 1740 692 1742 694
rect 1774 692 1776 694
rect 952 690 954 692
rect 1262 690 1264 692
rect 1562 690 1564 692
rect 1202 684 1204 686
rect 1502 684 1504 686
rect 1562 684 1564 686
rect 1672 684 1674 686
rect 944 682 946 684
rect 1200 682 1202 684
rect 1254 682 1256 684
rect 1500 682 1502 684
rect 1554 682 1556 684
rect 1560 682 1562 684
rect 1644 682 1646 684
rect 1670 682 1672 684
rect 942 680 944 682
rect 1252 680 1254 682
rect 1552 680 1554 682
rect 1642 680 1644 682
rect 1192 674 1194 676
rect 1492 674 1494 676
rect 1552 674 1554 676
rect 1662 674 1664 676
rect 934 672 936 674
rect 1190 672 1192 674
rect 1244 672 1246 674
rect 1490 672 1492 674
rect 1544 672 1546 674
rect 1550 672 1552 674
rect 1634 672 1636 674
rect 1660 672 1662 674
rect 932 670 934 672
rect 1242 670 1244 672
rect 1542 670 1544 672
rect 1632 670 1634 672
rect 1182 664 1184 666
rect 1482 664 1484 666
rect 1542 664 1544 666
rect 1652 664 1654 666
rect 924 662 926 664
rect 1180 662 1182 664
rect 1234 662 1236 664
rect 1480 662 1482 664
rect 1534 662 1536 664
rect 1540 662 1542 664
rect 1624 662 1626 664
rect 1650 662 1652 664
rect 922 660 924 662
rect 1232 660 1234 662
rect 1532 660 1534 662
rect 1622 660 1624 662
rect 1172 654 1174 656
rect 1472 654 1474 656
rect 1532 654 1534 656
rect 1642 654 1644 656
rect 914 652 916 654
rect 1170 652 1172 654
rect 1224 652 1226 654
rect 1470 652 1472 654
rect 1524 652 1526 654
rect 1530 652 1532 654
rect 1614 652 1616 654
rect 1640 652 1642 654
rect 912 650 914 652
rect 1222 650 1224 652
rect 1522 650 1524 652
rect 1612 650 1614 652
rect 1162 644 1164 646
rect 1462 644 1464 646
rect 1522 644 1524 646
rect 1632 644 1634 646
rect 904 642 906 644
rect 1160 642 1162 644
rect 1214 642 1216 644
rect 1460 642 1462 644
rect 1514 642 1516 644
rect 1520 642 1522 644
rect 1604 642 1606 644
rect 1630 642 1632 644
rect 902 640 904 642
rect 1212 640 1214 642
rect 1512 640 1514 642
rect 1602 640 1604 642
rect 1152 634 1154 636
rect 1452 634 1454 636
rect 1512 634 1514 636
rect 1622 634 1624 636
rect 1848 634 1850 636
rect 1878 634 1880 636
rect 1908 634 1910 636
rect 1938 634 1940 636
rect 1968 634 1970 636
rect 894 632 896 634
rect 1150 632 1152 634
rect 1204 632 1206 634
rect 1450 632 1452 634
rect 1504 632 1506 634
rect 1510 632 1512 634
rect 1594 632 1596 634
rect 1620 632 1622 634
rect 1820 632 1822 634
rect 1826 632 1828 634
rect 1850 632 1852 634
rect 1856 632 1858 634
rect 1880 632 1882 634
rect 1886 632 1888 634
rect 1910 632 1912 634
rect 1916 632 1918 634
rect 1940 632 1942 634
rect 1946 632 1948 634
rect 1970 632 1972 634
rect 1976 632 1978 634
rect 892 630 894 632
rect 1202 630 1204 632
rect 1502 630 1504 632
rect 1592 630 1594 632
rect 1818 630 1820 632
rect 1828 630 1830 632
rect 1858 630 1860 632
rect 1888 630 1890 632
rect 1918 630 1920 632
rect 1948 630 1950 632
rect 1978 630 1980 632
rect 1142 624 1144 626
rect 1442 624 1444 626
rect 1502 624 1504 626
rect 1612 624 1614 626
rect 1828 624 1830 626
rect 1858 624 1860 626
rect 1888 624 1890 626
rect 1918 624 1920 626
rect 1948 624 1950 626
rect 1978 624 1980 626
rect 884 622 886 624
rect 1140 622 1142 624
rect 1194 622 1196 624
rect 1440 622 1442 624
rect 1494 622 1496 624
rect 1500 622 1502 624
rect 1584 622 1586 624
rect 1610 622 1612 624
rect 1810 622 1812 624
rect 1826 622 1828 624
rect 1850 622 1852 624
rect 1856 622 1858 624
rect 1880 622 1882 624
rect 1886 622 1888 624
rect 1910 622 1912 624
rect 1916 622 1918 624
rect 1940 622 1942 624
rect 1946 622 1948 624
rect 1970 622 1972 624
rect 1976 622 1978 624
rect 882 620 884 622
rect 1192 620 1194 622
rect 1492 620 1494 622
rect 1582 620 1584 622
rect 1808 620 1810 622
rect 1848 620 1850 622
rect 1878 620 1880 622
rect 1908 620 1910 622
rect 1938 620 1940 622
rect 1968 620 1970 622
rect 1132 614 1134 616
rect 1432 614 1434 616
rect 1492 614 1494 616
rect 1602 614 1604 616
rect 1808 614 1810 616
rect 1818 614 1820 616
rect 1848 614 1850 616
rect 1878 614 1880 616
rect 1908 614 1910 616
rect 1938 614 1940 616
rect 1968 614 1970 616
rect 874 612 876 614
rect 1130 612 1132 614
rect 1184 612 1186 614
rect 1430 612 1432 614
rect 1484 612 1486 614
rect 1490 612 1492 614
rect 1574 612 1576 614
rect 1600 612 1602 614
rect 1800 612 1802 614
rect 1806 612 1808 614
rect 1820 612 1822 614
rect 1826 612 1828 614
rect 1850 612 1852 614
rect 1856 612 1858 614
rect 1880 612 1882 614
rect 1886 612 1888 614
rect 1910 612 1912 614
rect 1916 612 1918 614
rect 1940 612 1942 614
rect 1946 612 1948 614
rect 1970 612 1972 614
rect 1976 612 1978 614
rect 872 610 874 612
rect 1182 610 1184 612
rect 1482 610 1484 612
rect 1572 610 1574 612
rect 1798 610 1800 612
rect 1828 610 1830 612
rect 1858 610 1860 612
rect 1888 610 1890 612
rect 1918 610 1920 612
rect 1948 610 1950 612
rect 1978 610 1980 612
rect 1122 604 1124 606
rect 1422 604 1424 606
rect 1482 604 1484 606
rect 1592 604 1594 606
rect 1798 604 1800 606
rect 1828 604 1830 606
rect 1858 604 1860 606
rect 1888 604 1890 606
rect 1918 604 1920 606
rect 1948 604 1950 606
rect 1978 604 1980 606
rect 864 602 866 604
rect 1120 602 1122 604
rect 1174 602 1176 604
rect 1420 602 1422 604
rect 1474 602 1476 604
rect 1480 602 1482 604
rect 1564 602 1566 604
rect 1590 602 1592 604
rect 1790 602 1792 604
rect 1796 602 1798 604
rect 1820 602 1822 604
rect 1826 602 1828 604
rect 1850 602 1852 604
rect 1856 602 1858 604
rect 1880 602 1882 604
rect 1886 602 1888 604
rect 1910 602 1912 604
rect 1916 602 1918 604
rect 1940 602 1942 604
rect 1946 602 1948 604
rect 1970 602 1972 604
rect 1976 602 1978 604
rect 862 600 864 602
rect 1172 600 1174 602
rect 1472 600 1474 602
rect 1562 600 1564 602
rect 1788 600 1790 602
rect 1818 600 1820 602
rect 1848 600 1850 602
rect 1878 600 1880 602
rect 1908 600 1910 602
rect 1938 600 1940 602
rect 1968 600 1970 602
rect 1112 594 1114 596
rect 1412 594 1414 596
rect 1472 594 1474 596
rect 1582 594 1584 596
rect 1788 594 1790 596
rect 1848 594 1850 596
rect 1878 594 1880 596
rect 1908 594 1910 596
rect 1938 594 1940 596
rect 1968 594 1970 596
rect 854 592 856 594
rect 1110 592 1112 594
rect 1164 592 1166 594
rect 1410 592 1412 594
rect 1464 592 1466 594
rect 1470 592 1472 594
rect 1554 592 1556 594
rect 1580 592 1582 594
rect 1780 592 1782 594
rect 1786 592 1788 594
rect 1810 592 1812 594
rect 1826 592 1828 594
rect 1850 592 1852 594
rect 1856 592 1858 594
rect 1880 592 1882 594
rect 1886 592 1888 594
rect 1910 592 1912 594
rect 1916 592 1918 594
rect 1940 592 1942 594
rect 1946 592 1948 594
rect 1970 592 1972 594
rect 1976 592 1978 594
rect 852 590 854 592
rect 1162 590 1164 592
rect 1462 590 1464 592
rect 1552 590 1554 592
rect 1778 590 1780 592
rect 1808 590 1810 592
rect 1828 590 1830 592
rect 1858 590 1860 592
rect 1888 590 1890 592
rect 1918 590 1920 592
rect 1948 590 1950 592
rect 1978 590 1980 592
rect 1102 584 1104 586
rect 1402 584 1404 586
rect 1462 584 1464 586
rect 1572 584 1574 586
rect 1778 584 1780 586
rect 1808 584 1810 586
rect 1818 584 1820 586
rect 1828 584 1830 586
rect 1888 584 1890 586
rect 1918 584 1920 586
rect 1948 584 1950 586
rect 1978 584 1980 586
rect 844 582 846 584
rect 1100 582 1102 584
rect 1154 582 1156 584
rect 1400 582 1402 584
rect 1454 582 1456 584
rect 1460 582 1462 584
rect 1544 582 1546 584
rect 1570 582 1572 584
rect 1770 582 1772 584
rect 1776 582 1778 584
rect 1800 582 1802 584
rect 1806 582 1808 584
rect 1820 582 1822 584
rect 1826 582 1828 584
rect 1850 582 1852 584
rect 1866 582 1868 584
rect 1880 582 1882 584
rect 1886 582 1888 584
rect 1910 582 1912 584
rect 1916 582 1918 584
rect 1940 582 1942 584
rect 1946 582 1948 584
rect 1970 582 1972 584
rect 1976 582 1978 584
rect 842 580 844 582
rect 1152 580 1154 582
rect 1452 580 1454 582
rect 1542 580 1544 582
rect 1768 580 1770 582
rect 1798 580 1800 582
rect 1848 580 1850 582
rect 1868 580 1870 582
rect 1878 580 1880 582
rect 1908 580 1910 582
rect 1938 580 1940 582
rect 1968 580 1970 582
rect 1092 574 1094 576
rect 1392 574 1394 576
rect 1452 574 1454 576
rect 1562 574 1564 576
rect 1768 574 1770 576
rect 1798 574 1800 576
rect 1868 574 1870 576
rect 1878 574 1880 576
rect 1908 574 1910 576
rect 1938 574 1940 576
rect 1968 574 1970 576
rect 834 572 836 574
rect 1090 572 1092 574
rect 1144 572 1146 574
rect 1390 572 1392 574
rect 1444 572 1446 574
rect 1450 572 1452 574
rect 1534 572 1536 574
rect 1560 572 1562 574
rect 1760 572 1762 574
rect 1766 572 1768 574
rect 1790 572 1792 574
rect 1796 572 1798 574
rect 1820 572 1822 574
rect 1826 572 1828 574
rect 1840 572 1842 574
rect 1866 572 1868 574
rect 1880 572 1882 574
rect 1886 572 1888 574
rect 1910 572 1912 574
rect 1916 572 1918 574
rect 1940 572 1942 574
rect 1946 572 1948 574
rect 1970 572 1972 574
rect 1976 572 1978 574
rect 832 570 834 572
rect 1142 570 1144 572
rect 1442 570 1444 572
rect 1532 570 1534 572
rect 1758 570 1760 572
rect 1788 570 1790 572
rect 1818 570 1820 572
rect 1828 570 1830 572
rect 1838 570 1840 572
rect 1888 570 1890 572
rect 1918 570 1920 572
rect 1948 570 1950 572
rect 1978 570 1980 572
rect 1082 564 1084 566
rect 1382 564 1384 566
rect 1442 564 1444 566
rect 1552 564 1554 566
rect 1758 564 1760 566
rect 1788 564 1790 566
rect 1858 564 1860 566
rect 1888 564 1890 566
rect 1918 564 1920 566
rect 1948 564 1950 566
rect 1978 564 1980 566
rect 824 562 826 564
rect 1080 562 1082 564
rect 1134 562 1136 564
rect 1380 562 1382 564
rect 1434 562 1436 564
rect 1440 562 1442 564
rect 1524 562 1526 564
rect 1550 562 1552 564
rect 1750 562 1752 564
rect 1756 562 1758 564
rect 1780 562 1782 564
rect 1786 562 1788 564
rect 1810 562 1812 564
rect 1856 562 1858 564
rect 1880 562 1882 564
rect 1886 562 1888 564
rect 1910 562 1912 564
rect 1916 562 1918 564
rect 1940 562 1942 564
rect 1946 562 1948 564
rect 1970 562 1972 564
rect 1976 562 1978 564
rect 822 560 824 562
rect 1132 560 1134 562
rect 1432 560 1434 562
rect 1522 560 1524 562
rect 1748 560 1750 562
rect 1778 560 1780 562
rect 1808 560 1810 562
rect 1878 560 1880 562
rect 1908 560 1910 562
rect 1938 560 1940 562
rect 1968 560 1970 562
rect 1072 554 1074 556
rect 1372 554 1374 556
rect 1432 554 1434 556
rect 1542 554 1544 556
rect 1748 554 1750 556
rect 1778 554 1780 556
rect 1838 554 1840 556
rect 1848 554 1850 556
rect 1878 554 1880 556
rect 1908 554 1910 556
rect 1938 554 1940 556
rect 1968 554 1970 556
rect 814 552 816 554
rect 1070 552 1072 554
rect 1124 552 1126 554
rect 1370 552 1372 554
rect 1424 552 1426 554
rect 1430 552 1432 554
rect 1514 552 1516 554
rect 1540 552 1542 554
rect 1740 552 1742 554
rect 1746 552 1748 554
rect 1770 552 1772 554
rect 1776 552 1778 554
rect 1800 552 1802 554
rect 1836 552 1838 554
rect 1850 552 1852 554
rect 1856 552 1858 554
rect 1880 552 1882 554
rect 1886 552 1888 554
rect 1910 552 1912 554
rect 1916 552 1918 554
rect 1940 552 1942 554
rect 1946 552 1948 554
rect 1970 552 1972 554
rect 1976 552 1978 554
rect 812 550 814 552
rect 1122 550 1124 552
rect 1422 550 1424 552
rect 1512 550 1514 552
rect 1738 550 1740 552
rect 1768 550 1770 552
rect 1798 550 1800 552
rect 1858 550 1860 552
rect 1888 550 1890 552
rect 1918 550 1920 552
rect 1948 550 1950 552
rect 1978 550 1980 552
rect 1062 544 1064 546
rect 1362 544 1364 546
rect 1422 544 1424 546
rect 1532 544 1534 546
rect 1738 544 1740 546
rect 1768 544 1770 546
rect 1828 544 1830 546
rect 1858 544 1860 546
rect 1888 544 1890 546
rect 1918 544 1920 546
rect 1948 544 1950 546
rect 1978 544 1980 546
rect 804 542 806 544
rect 1060 542 1062 544
rect 1114 542 1116 544
rect 1360 542 1362 544
rect 1414 542 1416 544
rect 1420 542 1422 544
rect 1504 542 1506 544
rect 1530 542 1532 544
rect 1730 542 1732 544
rect 1736 542 1738 544
rect 1760 542 1762 544
rect 1766 542 1768 544
rect 1790 542 1792 544
rect 1826 542 1828 544
rect 1850 542 1852 544
rect 1856 542 1858 544
rect 1880 542 1882 544
rect 1886 542 1888 544
rect 1910 542 1912 544
rect 1916 542 1918 544
rect 1940 542 1942 544
rect 1946 542 1948 544
rect 1970 542 1972 544
rect 1976 542 1978 544
rect 802 540 804 542
rect 1112 540 1114 542
rect 1412 540 1414 542
rect 1502 540 1504 542
rect 1728 540 1730 542
rect 1758 540 1760 542
rect 1788 540 1790 542
rect 1848 540 1850 542
rect 1878 540 1880 542
rect 1908 540 1910 542
rect 1938 540 1940 542
rect 1968 540 1970 542
rect 1052 534 1054 536
rect 1352 534 1354 536
rect 1412 534 1414 536
rect 1522 534 1524 536
rect 1728 534 1730 536
rect 1758 534 1760 536
rect 1808 534 1810 536
rect 1818 534 1820 536
rect 1848 534 1850 536
rect 1878 534 1880 536
rect 1908 534 1910 536
rect 1938 534 1940 536
rect 1968 534 1970 536
rect 794 532 796 534
rect 1050 532 1052 534
rect 1104 532 1106 534
rect 1350 532 1352 534
rect 1404 532 1406 534
rect 1410 532 1412 534
rect 1494 532 1496 534
rect 1520 532 1522 534
rect 1720 532 1722 534
rect 1726 532 1728 534
rect 1750 532 1752 534
rect 1756 532 1758 534
rect 1780 532 1782 534
rect 792 530 794 532
rect 1102 530 1104 532
rect 1402 530 1404 532
rect 1492 530 1494 532
rect 1718 530 1720 532
rect 1748 530 1750 532
rect 1778 530 1780 532
rect 1806 531 1808 534
rect 1820 531 1822 534
rect 1826 532 1828 534
rect 1850 532 1852 534
rect 1856 532 1858 534
rect 1880 532 1882 534
rect 1886 532 1888 534
rect 1910 532 1912 534
rect 1916 532 1918 534
rect 1940 532 1942 534
rect 1946 532 1948 534
rect 1970 532 1972 534
rect 1976 532 1978 534
rect 1808 529 1810 531
rect 1818 529 1820 531
rect 1828 530 1830 532
rect 1858 530 1860 532
rect 1888 530 1890 532
rect 1918 530 1920 532
rect 1948 530 1950 532
rect 1978 530 1980 532
rect 1042 524 1044 526
rect 1342 524 1344 526
rect 1402 524 1404 526
rect 1512 524 1514 526
rect 1718 524 1720 526
rect 1748 524 1750 526
rect 784 522 786 524
rect 1040 522 1042 524
rect 1094 522 1096 524
rect 1340 522 1342 524
rect 1394 522 1396 524
rect 1400 522 1402 524
rect 1484 522 1486 524
rect 1510 522 1512 524
rect 1710 522 1712 524
rect 1716 522 1718 524
rect 1740 522 1742 524
rect 1746 522 1748 524
rect 1770 522 1772 524
rect 1808 523 1810 525
rect 1818 523 1820 525
rect 1828 524 1830 526
rect 1858 524 1860 526
rect 1888 524 1890 526
rect 1918 524 1920 526
rect 1948 524 1950 526
rect 1978 524 1980 526
rect 782 520 784 522
rect 1092 520 1094 522
rect 1392 520 1394 522
rect 1482 520 1484 522
rect 1708 520 1710 522
rect 1738 520 1740 522
rect 1768 520 1770 522
rect 1806 521 1808 523
rect 1820 521 1822 523
rect 1826 522 1828 524
rect 1850 522 1852 524
rect 1856 522 1858 524
rect 1880 522 1882 524
rect 1886 522 1888 524
rect 1910 522 1912 524
rect 1916 522 1918 524
rect 1940 522 1942 524
rect 1946 522 1948 524
rect 1970 522 1972 524
rect 1976 522 1978 524
rect 1848 520 1850 522
rect 1878 520 1880 522
rect 1908 520 1910 522
rect 1938 520 1940 522
rect 1968 520 1970 522
rect 1032 514 1034 516
rect 1332 514 1334 516
rect 1392 514 1394 516
rect 1502 514 1504 516
rect 1708 514 1710 516
rect 1738 514 1740 516
rect 1798 514 1800 516
rect 1848 514 1850 516
rect 1878 514 1880 516
rect 1908 514 1910 516
rect 1938 514 1940 516
rect 1968 514 1970 516
rect 774 512 776 514
rect 1030 512 1032 514
rect 1084 512 1086 514
rect 1330 512 1332 514
rect 1384 512 1386 514
rect 1390 512 1392 514
rect 1474 512 1476 514
rect 1500 512 1502 514
rect 1700 512 1702 514
rect 1706 512 1708 514
rect 1730 512 1732 514
rect 1736 512 1738 514
rect 1760 512 1762 514
rect 1796 512 1798 514
rect 1820 512 1822 514
rect 1826 512 1828 514
rect 1850 512 1852 514
rect 1856 512 1858 514
rect 1880 512 1882 514
rect 1886 512 1888 514
rect 1910 512 1912 514
rect 1916 512 1918 514
rect 1940 512 1942 514
rect 1946 512 1948 514
rect 1970 512 1972 514
rect 1976 512 1978 514
rect 772 510 774 512
rect 1082 510 1084 512
rect 1382 510 1384 512
rect 1472 510 1474 512
rect 1698 510 1700 512
rect 1728 510 1730 512
rect 1758 510 1760 512
rect 1818 510 1820 512
rect 1828 510 1830 512
rect 1858 510 1860 512
rect 1888 510 1890 512
rect 1918 510 1920 512
rect 1948 510 1950 512
rect 1978 510 1980 512
rect 1022 504 1024 506
rect 1322 504 1324 506
rect 1382 504 1384 506
rect 1492 504 1494 506
rect 764 502 766 504
rect 1020 502 1022 504
rect 1074 502 1076 504
rect 1320 502 1322 504
rect 1374 502 1376 504
rect 1380 502 1382 504
rect 1464 502 1466 504
rect 1490 502 1492 504
rect 1690 502 1692 504
rect 1706 502 1708 504
rect 1720 502 1722 504
rect 1736 502 1738 504
rect 1750 502 1752 504
rect 1796 502 1798 504
rect 1810 502 1812 504
rect 1836 502 1838 504
rect 1850 502 1852 504
rect 1866 502 1868 504
rect 1880 502 1882 504
rect 1896 502 1898 504
rect 1910 502 1912 504
rect 1926 502 1928 504
rect 1940 502 1942 504
rect 1956 502 1958 504
rect 1970 502 1972 504
rect 1986 502 1988 504
rect 762 500 764 502
rect 1072 500 1074 502
rect 1372 500 1374 502
rect 1462 500 1464 502
rect 1688 500 1690 502
rect 1708 500 1710 502
rect 1718 500 1720 502
rect 1738 500 1740 502
rect 1748 500 1750 502
rect 1798 500 1800 502
rect 1808 500 1810 502
rect 1838 500 1840 502
rect 1848 500 1850 502
rect 1868 500 1870 502
rect 1878 500 1880 502
rect 1898 500 1900 502
rect 1908 500 1910 502
rect 1928 500 1930 502
rect 1938 500 1940 502
rect 1958 500 1960 502
rect 1968 500 1970 502
rect 1988 500 1990 502
rect 1012 494 1014 496
rect 1312 494 1314 496
rect 1372 494 1374 496
rect 1482 494 1484 496
rect 1688 494 1690 496
rect 1698 494 1700 496
rect 1708 494 1710 496
rect 1718 494 1720 496
rect 1728 494 1730 496
rect 1738 494 1740 496
rect 1748 494 1750 496
rect 1788 494 1790 496
rect 1798 494 1800 496
rect 1808 494 1810 496
rect 1818 494 1820 496
rect 1828 494 1830 496
rect 1838 494 1840 496
rect 1848 494 1850 496
rect 1858 494 1860 496
rect 1868 494 1870 496
rect 1888 494 1890 496
rect 754 492 756 494
rect 1010 492 1012 494
rect 1064 492 1066 494
rect 1310 492 1312 494
rect 1364 492 1366 494
rect 1370 492 1372 494
rect 1454 492 1456 494
rect 1480 492 1482 494
rect 1690 492 1692 494
rect 1696 492 1698 494
rect 1710 492 1712 494
rect 1716 492 1718 494
rect 1730 492 1732 494
rect 1736 492 1738 494
rect 1750 492 1752 494
rect 1786 492 1788 494
rect 1800 492 1802 494
rect 1806 492 1808 494
rect 1820 492 1822 494
rect 1826 492 1828 494
rect 1840 492 1842 494
rect 1846 492 1848 494
rect 1860 492 1862 494
rect 1866 492 1868 494
rect 1890 492 1892 494
rect 752 490 754 492
rect 1062 490 1064 492
rect 1362 490 1364 492
rect 1452 490 1454 492
rect 1002 484 1004 486
rect 1302 484 1304 486
rect 1362 484 1364 486
rect 1472 484 1474 486
rect 1778 484 1780 486
rect 744 482 746 484
rect 1000 482 1002 484
rect 1054 482 1056 484
rect 1300 482 1302 484
rect 1354 482 1356 484
rect 1360 482 1362 484
rect 1444 482 1446 484
rect 1470 482 1472 484
rect 1750 482 1752 484
rect 1776 482 1778 484
rect 1890 482 1892 484
rect 742 480 744 482
rect 1052 480 1054 482
rect 1352 480 1354 482
rect 1442 480 1444 482
rect 1748 480 1750 482
rect 1888 480 1890 482
rect 992 474 994 476
rect 1292 474 1294 476
rect 1352 474 1354 476
rect 1462 474 1464 476
rect 1768 474 1770 476
rect 734 472 736 474
rect 990 472 992 474
rect 1044 472 1046 474
rect 1290 472 1292 474
rect 1344 472 1346 474
rect 1350 472 1352 474
rect 1434 472 1436 474
rect 1460 472 1462 474
rect 1740 472 1742 474
rect 1766 472 1768 474
rect 1880 472 1882 474
rect 732 470 734 472
rect 1042 470 1044 472
rect 1342 470 1344 472
rect 1432 470 1434 472
rect 1738 470 1740 472
rect 1878 470 1880 472
rect 982 464 984 466
rect 1282 464 1284 466
rect 1342 464 1344 466
rect 1452 464 1454 466
rect 1758 464 1760 466
rect 724 462 726 464
rect 980 462 982 464
rect 1034 462 1036 464
rect 1280 462 1282 464
rect 1334 462 1336 464
rect 1340 462 1342 464
rect 1424 462 1426 464
rect 1450 462 1452 464
rect 1730 462 1732 464
rect 1756 462 1758 464
rect 1870 462 1872 464
rect 722 460 724 462
rect 1032 460 1034 462
rect 1332 460 1334 462
rect 1422 460 1424 462
rect 1728 460 1730 462
rect 1868 460 1870 462
rect 972 454 974 456
rect 1272 454 1274 456
rect 1332 454 1334 456
rect 1442 454 1444 456
rect 1748 454 1750 456
rect 714 452 716 454
rect 970 452 972 454
rect 1024 452 1026 454
rect 1270 452 1272 454
rect 1324 452 1326 454
rect 1330 452 1332 454
rect 1414 452 1416 454
rect 1440 452 1442 454
rect 1720 452 1722 454
rect 1746 452 1748 454
rect 1860 452 1862 454
rect 712 450 714 452
rect 1022 450 1024 452
rect 1322 450 1324 452
rect 1412 450 1414 452
rect 1718 450 1720 452
rect 1858 450 1860 452
rect 962 444 964 446
rect 1262 444 1264 446
rect 1322 444 1324 446
rect 1432 444 1434 446
rect 1738 444 1740 446
rect 704 442 706 444
rect 960 442 962 444
rect 1014 442 1016 444
rect 1260 442 1262 444
rect 1314 442 1316 444
rect 1320 442 1322 444
rect 1404 442 1406 444
rect 1430 442 1432 444
rect 1710 442 1712 444
rect 1736 442 1738 444
rect 1850 442 1852 444
rect 702 440 704 442
rect 1012 440 1014 442
rect 1312 440 1314 442
rect 1402 440 1404 442
rect 1708 440 1710 442
rect 1848 440 1850 442
rect 952 434 954 436
rect 1252 434 1254 436
rect 1312 434 1314 436
rect 1422 434 1424 436
rect 1728 434 1730 436
rect 694 432 696 434
rect 950 432 952 434
rect 1004 432 1006 434
rect 1250 432 1252 434
rect 1304 432 1306 434
rect 1310 432 1312 434
rect 1394 432 1396 434
rect 1420 432 1422 434
rect 1700 432 1702 434
rect 1726 432 1728 434
rect 1840 432 1842 434
rect 692 430 694 432
rect 1002 430 1004 432
rect 1302 430 1304 432
rect 1392 430 1394 432
rect 1698 430 1700 432
rect 1838 430 1840 432
rect 942 424 944 426
rect 1242 424 1244 426
rect 1302 424 1304 426
rect 1412 424 1414 426
rect 1718 424 1720 426
rect 684 422 686 424
rect 940 422 942 424
rect 994 422 996 424
rect 1240 422 1242 424
rect 1294 422 1296 424
rect 1300 422 1302 424
rect 1384 422 1386 424
rect 1410 422 1412 424
rect 1690 422 1692 424
rect 1716 422 1718 424
rect 682 420 684 422
rect 992 420 994 422
rect 1292 420 1294 422
rect 1382 420 1384 422
rect 1688 420 1690 422
rect 932 414 934 416
rect 1232 414 1234 416
rect 1292 414 1294 416
rect 1402 414 1404 416
rect 1708 414 1710 416
rect 1838 414 1840 416
rect 674 412 676 414
rect 930 412 932 414
rect 984 412 986 414
rect 1230 412 1232 414
rect 1284 412 1286 414
rect 1290 412 1292 414
rect 1374 412 1376 414
rect 1400 412 1402 414
rect 1680 412 1682 414
rect 1706 412 1708 414
rect 1840 412 1842 414
rect 672 410 674 412
rect 982 410 984 412
rect 1282 410 1284 412
rect 1372 410 1374 412
rect 1678 410 1680 412
rect 1222 404 1224 406
rect 1282 404 1284 406
rect 1392 404 1394 406
rect 1698 404 1700 406
rect 974 402 976 404
rect 1220 402 1222 404
rect 1274 402 1276 404
rect 1280 402 1282 404
rect 1364 402 1366 404
rect 1390 402 1392 404
rect 1670 402 1672 404
rect 1696 402 1698 404
rect 1840 402 1842 404
rect 972 400 974 402
rect 1272 400 1274 402
rect 1362 400 1364 402
rect 1668 400 1670 402
rect 1838 400 1840 402
rect 1212 394 1214 396
rect 1272 394 1274 396
rect 1382 394 1384 396
rect 1688 394 1690 396
rect 964 392 966 394
rect 1210 392 1212 394
rect 1264 392 1266 394
rect 1270 392 1272 394
rect 1354 392 1356 394
rect 1380 392 1382 394
rect 1660 392 1662 394
rect 1686 392 1688 394
rect 1830 392 1832 394
rect 962 390 964 392
rect 1262 390 1264 392
rect 1352 390 1354 392
rect 1658 390 1660 392
rect 1828 390 1830 392
rect 1202 384 1204 386
rect 1262 384 1264 386
rect 1372 384 1374 386
rect 1678 384 1680 386
rect 930 382 932 384
rect 954 382 956 384
rect 1200 382 1202 384
rect 1254 382 1256 384
rect 1260 382 1262 384
rect 1344 382 1346 384
rect 1370 382 1372 384
rect 1650 382 1652 384
rect 1676 382 1678 384
rect 1820 382 1822 384
rect 932 380 934 382
rect 952 380 954 382
rect 1252 380 1254 382
rect 1342 380 1344 382
rect 1648 380 1650 382
rect 1818 380 1820 382
rect 1192 374 1194 376
rect 1252 374 1254 376
rect 1362 374 1364 376
rect 1668 374 1670 376
rect 1190 372 1192 374
rect 1244 372 1246 374
rect 1250 372 1252 374
rect 1334 372 1336 374
rect 1360 372 1362 374
rect 1640 372 1642 374
rect 1666 372 1668 374
rect 1810 372 1812 374
rect 1242 370 1244 372
rect 1332 370 1334 372
rect 1638 370 1640 372
rect 1808 370 1810 372
rect 1182 364 1184 366
rect 1242 364 1244 366
rect 1352 364 1354 366
rect 1658 364 1660 366
rect 1180 362 1182 364
rect 1234 362 1236 364
rect 1240 362 1242 364
rect 1324 362 1326 364
rect 1350 362 1352 364
rect 1630 362 1632 364
rect 1656 362 1658 364
rect 1800 362 1802 364
rect 1232 360 1234 362
rect 1322 360 1324 362
rect 1628 360 1630 362
rect 1798 360 1800 362
rect 1172 354 1174 356
rect 1232 354 1234 356
rect 1342 354 1344 356
rect 1648 354 1650 356
rect 1170 352 1172 354
rect 1224 352 1226 354
rect 1230 352 1232 354
rect 1314 352 1316 354
rect 1340 352 1342 354
rect 1620 352 1622 354
rect 1646 352 1648 354
rect 1790 352 1792 354
rect 1222 350 1224 352
rect 1312 350 1314 352
rect 1618 350 1620 352
rect 1788 350 1790 352
rect 1162 344 1164 346
rect 1222 344 1224 346
rect 1332 344 1334 346
rect 1638 344 1640 346
rect 1160 342 1162 344
rect 1214 342 1216 344
rect 1220 342 1222 344
rect 1304 342 1306 344
rect 1330 342 1332 344
rect 1610 342 1612 344
rect 1636 342 1638 344
rect 1780 342 1782 344
rect 1212 340 1214 342
rect 1302 340 1304 342
rect 1608 340 1610 342
rect 1778 340 1780 342
rect 1152 334 1154 336
rect 1212 334 1214 336
rect 1322 334 1324 336
rect 1628 334 1630 336
rect 1150 332 1152 334
rect 1204 332 1206 334
rect 1210 332 1212 334
rect 1294 332 1296 334
rect 1320 332 1322 334
rect 1600 332 1602 334
rect 1626 332 1628 334
rect 1770 332 1772 334
rect 1202 330 1204 332
rect 1292 330 1294 332
rect 1598 330 1600 332
rect 1768 330 1770 332
rect 1142 324 1144 326
rect 1202 324 1204 326
rect 1312 324 1314 326
rect 1618 324 1620 326
rect 1140 322 1142 324
rect 1194 322 1196 324
rect 1200 322 1202 324
rect 1284 322 1286 324
rect 1310 322 1312 324
rect 1590 322 1592 324
rect 1616 322 1618 324
rect 1760 322 1762 324
rect 1192 320 1194 322
rect 1282 320 1284 322
rect 1588 320 1590 322
rect 1758 320 1760 322
rect 1132 314 1134 316
rect 1192 314 1194 316
rect 1302 314 1304 316
rect 1608 314 1610 316
rect 1130 312 1132 314
rect 1184 312 1186 314
rect 1190 312 1192 314
rect 1274 312 1276 314
rect 1300 312 1302 314
rect 1580 312 1582 314
rect 1606 312 1608 314
rect 1750 312 1752 314
rect 1182 310 1184 312
rect 1272 310 1274 312
rect 1578 310 1580 312
rect 1748 310 1750 312
rect 1122 304 1124 306
rect 1182 304 1184 306
rect 1292 304 1294 306
rect 1598 304 1600 306
rect 1120 302 1122 304
rect 1174 302 1176 304
rect 1180 302 1182 304
rect 1264 302 1266 304
rect 1290 302 1292 304
rect 1570 302 1572 304
rect 1596 302 1598 304
rect 1740 302 1742 304
rect 1172 300 1174 302
rect 1262 300 1264 302
rect 1568 300 1570 302
rect 1112 294 1114 296
rect 1172 294 1174 296
rect 1282 294 1284 296
rect 1578 294 1580 302
rect 1738 300 1740 302
rect 1588 294 1590 296
rect 1110 292 1112 294
rect 1164 292 1166 294
rect 1170 292 1172 294
rect 1254 292 1256 294
rect 1280 292 1282 294
rect 1560 292 1562 294
rect 1576 292 1580 294
rect 1586 292 1588 294
rect 1730 292 1732 294
rect 1162 290 1164 292
rect 1252 290 1254 292
rect 1558 290 1560 292
rect 1574 290 1580 292
rect 1728 290 1730 292
rect 1162 284 1164 286
rect 1272 284 1274 286
rect 1578 284 1580 286
rect 1154 282 1156 284
rect 1160 282 1162 284
rect 1244 282 1246 284
rect 1270 282 1272 284
rect 1550 282 1552 284
rect 1576 282 1578 284
rect 1720 282 1722 284
rect 1152 280 1154 282
rect 1242 280 1244 282
rect 1268 278 1270 282
rect 1548 280 1550 282
rect 1718 280 1720 282
rect 1092 274 1094 276
rect 1152 274 1154 276
rect 1262 274 1264 276
rect 1568 274 1570 276
rect 1090 272 1092 274
rect 1144 272 1146 274
rect 1150 272 1152 274
rect 1234 272 1236 274
rect 1260 272 1262 274
rect 1540 272 1542 274
rect 1566 272 1568 274
rect 1710 272 1712 274
rect 1142 270 1144 272
rect 1232 270 1234 272
rect 1538 270 1540 272
rect 1708 270 1710 272
rect 1232 264 1234 266
rect 1242 264 1244 266
rect 1558 264 1560 266
rect 1190 262 1192 264
rect 1224 262 1226 264
rect 1230 262 1232 264
rect 1244 262 1246 264
rect 1280 262 1282 264
rect 1314 262 1316 264
rect 1340 262 1342 264
rect 1530 262 1532 264
rect 1556 262 1558 264
rect 1700 262 1702 264
rect 1192 260 1194 262
rect 1222 260 1224 262
rect 1282 260 1284 262
rect 1312 260 1314 262
rect 1342 260 1344 262
rect 1528 260 1530 262
rect 1698 260 1700 262
rect 1342 254 1344 256
rect 1548 254 1550 256
rect 1340 252 1342 254
rect 1520 252 1522 254
rect 1546 252 1548 254
rect 1690 252 1692 254
rect 1518 250 1520 252
rect 1688 250 1690 252
rect 1192 244 1194 246
rect 1222 244 1224 246
rect 1252 244 1254 246
rect 1282 244 1284 246
rect 1312 244 1314 246
rect 1538 244 1540 246
rect 1090 242 1092 244
rect 1134 242 1136 244
rect 1150 242 1152 244
rect 1184 242 1186 244
rect 1190 242 1192 244
rect 1214 242 1216 244
rect 1220 242 1222 244
rect 1244 242 1246 244
rect 1250 242 1252 244
rect 1274 242 1276 244
rect 1280 242 1282 244
rect 1304 242 1306 244
rect 1310 242 1312 244
rect 1510 242 1512 244
rect 1536 242 1538 244
rect 1680 242 1682 244
rect 1092 240 1094 242
rect 1132 240 1134 242
rect 1152 240 1154 242
rect 1182 240 1184 242
rect 1212 240 1214 242
rect 1242 240 1244 242
rect 1272 240 1274 242
rect 1302 240 1304 242
rect 1508 240 1510 242
rect 1678 240 1680 242
rect 1182 234 1184 236
rect 1212 234 1214 236
rect 1242 234 1244 236
rect 1272 234 1274 236
rect 1302 234 1304 236
rect 1528 234 1530 236
rect 1160 232 1162 234
rect 1184 232 1186 234
rect 1190 232 1192 234
rect 1214 232 1216 234
rect 1220 232 1222 234
rect 1244 232 1246 234
rect 1250 232 1252 234
rect 1274 232 1276 234
rect 1280 232 1282 234
rect 1304 232 1306 234
rect 1310 232 1312 234
rect 1500 232 1502 234
rect 1526 232 1528 234
rect 1670 232 1672 234
rect 1162 230 1164 232
rect 1192 230 1194 232
rect 1222 230 1224 232
rect 1252 230 1254 232
rect 1282 230 1284 232
rect 1312 230 1314 232
rect 1498 230 1500 232
rect 1668 230 1670 232
rect 1162 224 1164 226
rect 1192 224 1194 226
rect 1222 224 1224 226
rect 1252 224 1254 226
rect 1282 224 1284 226
rect 1312 224 1314 226
rect 1518 224 1520 226
rect 1160 222 1162 224
rect 1184 222 1186 224
rect 1190 222 1192 224
rect 1214 222 1216 224
rect 1220 222 1222 224
rect 1244 222 1246 224
rect 1250 222 1252 224
rect 1274 222 1276 224
rect 1280 222 1282 224
rect 1304 222 1306 224
rect 1310 222 1312 224
rect 1490 222 1492 224
rect 1516 222 1518 224
rect 1660 222 1662 224
rect 1182 220 1184 222
rect 1212 220 1214 222
rect 1242 220 1244 222
rect 1272 220 1274 222
rect 1302 220 1304 222
rect 1488 220 1490 222
rect 1658 220 1660 222
rect 1182 214 1184 216
rect 1212 214 1214 216
rect 1242 214 1244 216
rect 1272 214 1274 216
rect 1302 214 1304 216
rect 1508 214 1510 216
rect 1160 212 1162 214
rect 1184 212 1186 214
rect 1190 212 1192 214
rect 1214 212 1216 214
rect 1220 212 1222 214
rect 1244 212 1246 214
rect 1250 212 1252 214
rect 1274 212 1276 214
rect 1280 212 1282 214
rect 1304 212 1306 214
rect 1480 212 1482 214
rect 1506 212 1508 214
rect 1650 212 1652 214
rect 1162 210 1164 212
rect 1192 210 1194 212
rect 1222 210 1224 212
rect 1252 210 1254 212
rect 1282 210 1284 212
rect 1478 210 1480 212
rect 1648 210 1650 212
rect 1162 204 1164 206
rect 1192 204 1194 206
rect 1222 204 1224 206
rect 1252 204 1254 206
rect 1282 204 1284 206
rect 1498 204 1500 206
rect 1160 202 1162 204
rect 1184 202 1186 204
rect 1190 202 1192 204
rect 1214 202 1216 204
rect 1220 202 1222 204
rect 1244 202 1246 204
rect 1250 202 1252 204
rect 1274 202 1276 204
rect 1280 202 1282 204
rect 1304 202 1306 204
rect 1470 202 1472 204
rect 1496 202 1498 204
rect 1640 202 1642 204
rect 1182 200 1184 202
rect 1212 200 1214 202
rect 1242 200 1244 202
rect 1272 200 1274 202
rect 1302 200 1304 202
rect 1468 200 1470 202
rect 1638 200 1640 202
rect 1182 194 1184 196
rect 1212 194 1214 196
rect 1242 194 1244 196
rect 1272 194 1274 196
rect 1302 194 1304 196
rect 1488 194 1490 196
rect 1160 192 1162 194
rect 1184 192 1186 194
rect 1190 192 1192 194
rect 1214 192 1216 194
rect 1220 192 1222 194
rect 1244 192 1246 194
rect 1250 192 1252 194
rect 1274 192 1276 194
rect 1280 192 1282 194
rect 1304 192 1306 194
rect 1460 192 1462 194
rect 1486 192 1488 194
rect 1630 192 1632 194
rect 1162 190 1164 192
rect 1192 190 1194 192
rect 1222 190 1224 192
rect 1252 190 1254 192
rect 1282 190 1284 192
rect 1458 190 1460 192
rect 1628 190 1630 192
rect 1162 184 1164 186
rect 1192 184 1194 186
rect 1222 184 1224 186
rect 1252 184 1254 186
rect 1282 184 1284 186
rect 1160 182 1162 184
rect 1184 182 1186 184
rect 1190 182 1192 184
rect 1214 182 1216 184
rect 1220 182 1222 184
rect 1244 182 1246 184
rect 1250 182 1252 184
rect 1274 182 1276 184
rect 1280 182 1282 184
rect 1304 182 1306 184
rect 1370 182 1372 184
rect 1376 182 1378 184
rect 1390 182 1392 184
rect 1396 182 1398 184
rect 1410 182 1412 184
rect 1416 182 1418 184
rect 1430 182 1432 184
rect 1436 182 1438 184
rect 1450 182 1452 184
rect 1486 182 1488 184
rect 1500 182 1502 184
rect 1506 182 1508 184
rect 1520 182 1522 184
rect 1526 182 1528 184
rect 1540 182 1542 184
rect 1546 182 1548 184
rect 1560 182 1562 184
rect 1620 182 1622 184
rect 1182 180 1184 182
rect 1212 180 1214 182
rect 1242 180 1244 182
rect 1272 180 1274 182
rect 1302 180 1304 182
rect 1368 180 1370 182
rect 1378 180 1380 182
rect 1388 180 1390 182
rect 1398 180 1400 182
rect 1408 180 1410 182
rect 1418 180 1420 182
rect 1428 180 1430 182
rect 1438 180 1440 182
rect 1448 180 1450 182
rect 1488 180 1490 182
rect 1498 180 1500 182
rect 1508 180 1510 182
rect 1518 180 1520 182
rect 1528 180 1530 182
rect 1538 180 1540 182
rect 1548 180 1550 182
rect 1558 180 1560 182
rect 1618 180 1620 182
rect 1182 174 1184 176
rect 1212 174 1214 176
rect 1242 174 1244 176
rect 1272 174 1274 176
rect 1302 174 1304 176
rect 1368 174 1370 176
rect 1378 174 1380 176
rect 1388 174 1390 176
rect 1398 174 1400 176
rect 1408 174 1410 176
rect 1418 174 1420 176
rect 1428 174 1430 176
rect 1468 174 1470 176
rect 1478 174 1480 176
rect 1488 174 1490 176
rect 1498 174 1500 176
rect 1508 174 1510 176
rect 1518 174 1520 176
rect 1528 174 1530 176
rect 1538 174 1540 176
rect 1548 174 1550 176
rect 1160 172 1162 174
rect 1184 172 1186 174
rect 1190 172 1192 174
rect 1214 172 1216 174
rect 1220 172 1222 174
rect 1244 172 1246 174
rect 1250 172 1252 174
rect 1274 172 1276 174
rect 1280 172 1282 174
rect 1304 172 1306 174
rect 1370 172 1372 174
rect 1376 172 1378 174
rect 1390 172 1392 174
rect 1396 172 1398 174
rect 1410 172 1412 174
rect 1416 172 1418 174
rect 1430 172 1432 174
rect 1466 172 1468 174
rect 1480 172 1482 174
rect 1486 172 1488 174
rect 1500 172 1502 174
rect 1506 172 1508 174
rect 1520 172 1522 174
rect 1526 172 1528 174
rect 1540 172 1542 174
rect 1546 172 1548 174
rect 1610 172 1612 174
rect 1162 170 1164 172
rect 1192 170 1194 172
rect 1222 170 1224 172
rect 1252 170 1254 172
rect 1282 170 1284 172
rect 1608 170 1610 172
rect 1162 164 1164 166
rect 1192 164 1194 166
rect 1222 164 1224 166
rect 1252 164 1254 166
rect 1282 164 1284 166
rect 1160 162 1162 164
rect 1184 162 1186 164
rect 1190 162 1192 164
rect 1214 162 1216 164
rect 1220 162 1222 164
rect 1244 162 1246 164
rect 1250 162 1252 164
rect 1274 162 1276 164
rect 1280 162 1282 164
rect 1304 162 1306 164
rect 1600 162 1602 164
rect 1182 160 1184 162
rect 1212 160 1214 162
rect 1242 160 1244 162
rect 1272 160 1274 162
rect 1302 160 1304 162
rect 1598 160 1600 162
rect 1182 154 1184 156
rect 1212 154 1214 156
rect 1242 154 1244 156
rect 1272 154 1274 156
rect 1302 154 1304 156
rect 1160 152 1162 154
rect 1184 152 1186 154
rect 1190 152 1192 154
rect 1214 152 1216 154
rect 1220 152 1222 154
rect 1244 152 1246 154
rect 1250 152 1252 154
rect 1274 152 1276 154
rect 1280 152 1282 154
rect 1304 152 1306 154
rect 1590 152 1592 154
rect 1162 150 1164 152
rect 1192 150 1194 152
rect 1222 150 1224 152
rect 1252 150 1254 152
rect 1282 150 1284 152
rect 1588 150 1590 152
rect 1162 144 1164 146
rect 1192 144 1194 146
rect 1222 144 1224 146
rect 1252 144 1254 146
rect 1282 144 1284 146
rect 1438 144 1440 146
rect 1458 144 1460 146
rect 1160 142 1162 144
rect 1184 142 1186 144
rect 1190 142 1192 144
rect 1214 142 1216 144
rect 1220 142 1222 144
rect 1244 142 1246 144
rect 1250 142 1252 144
rect 1274 142 1276 144
rect 1280 142 1282 144
rect 1304 142 1306 144
rect 1356 142 1358 144
rect 1390 142 1392 144
rect 1416 142 1418 144
rect 1440 142 1442 144
rect 1456 142 1458 144
rect 1480 142 1482 144
rect 1506 142 1508 144
rect 1520 142 1522 144
rect 1526 142 1528 144
rect 1540 142 1542 144
rect 1546 142 1548 144
rect 1580 142 1582 144
rect 1182 140 1184 142
rect 1212 140 1214 142
rect 1242 140 1244 142
rect 1272 140 1274 142
rect 1302 140 1304 142
rect 1358 140 1360 142
rect 1388 140 1390 142
rect 1418 140 1420 142
rect 1478 140 1480 142
rect 1508 140 1510 142
rect 1518 140 1520 142
rect 1528 140 1530 142
rect 1538 140 1540 142
rect 1548 140 1550 142
rect 1578 140 1580 142
rect 1182 134 1184 136
rect 1212 134 1214 136
rect 1242 134 1244 136
rect 1272 134 1274 136
rect 1302 134 1304 136
rect 1358 134 1360 136
rect 1388 134 1390 136
rect 1418 134 1420 136
rect 1448 134 1450 136
rect 1478 134 1480 136
rect 1160 132 1162 134
rect 1184 132 1186 134
rect 1190 132 1192 134
rect 1214 132 1216 134
rect 1220 132 1222 134
rect 1244 132 1246 134
rect 1250 132 1252 134
rect 1274 132 1276 134
rect 1280 132 1282 134
rect 1304 132 1306 134
rect 1356 132 1358 134
rect 1380 132 1382 134
rect 1386 132 1388 134
rect 1410 132 1412 134
rect 1416 132 1418 134
rect 1440 132 1442 134
rect 1446 132 1448 134
rect 1470 132 1472 134
rect 1476 132 1478 134
rect 1500 132 1502 134
rect 1162 130 1164 132
rect 1192 130 1194 132
rect 1222 130 1224 132
rect 1252 130 1254 132
rect 1282 130 1284 132
rect 1378 130 1380 132
rect 1408 130 1410 132
rect 1438 130 1440 132
rect 1468 130 1470 132
rect 1498 130 1500 132
rect 1162 124 1164 126
rect 1192 124 1194 126
rect 1222 124 1224 126
rect 1252 124 1254 126
rect 1282 124 1284 126
rect 1378 124 1380 126
rect 1408 124 1410 126
rect 1438 124 1440 126
rect 1468 124 1470 126
rect 1498 124 1500 126
rect 1160 122 1162 124
rect 1184 122 1186 124
rect 1190 122 1192 124
rect 1214 122 1216 124
rect 1220 122 1222 124
rect 1244 122 1246 124
rect 1250 122 1252 124
rect 1274 122 1276 124
rect 1280 122 1282 124
rect 1304 122 1306 124
rect 1356 122 1358 124
rect 1380 122 1382 124
rect 1386 122 1388 124
rect 1410 122 1412 124
rect 1416 122 1418 124
rect 1440 122 1442 124
rect 1446 122 1448 124
rect 1470 122 1472 124
rect 1476 122 1478 124
rect 1500 122 1502 124
rect 1182 120 1184 122
rect 1212 120 1214 122
rect 1242 120 1244 122
rect 1272 120 1274 122
rect 1302 120 1304 122
rect 1358 120 1360 122
rect 1388 120 1390 122
rect 1418 120 1420 122
rect 1448 120 1450 122
rect 1478 120 1480 122
rect 1182 114 1184 116
rect 1212 114 1214 116
rect 1242 114 1244 116
rect 1272 114 1274 116
rect 1302 114 1304 116
rect 1358 114 1360 116
rect 1388 114 1390 116
rect 1418 114 1420 116
rect 1448 114 1450 116
rect 1478 114 1480 116
rect 1160 112 1162 114
rect 1184 112 1186 114
rect 1190 112 1192 114
rect 1214 112 1216 114
rect 1220 112 1222 114
rect 1244 112 1246 114
rect 1250 112 1252 114
rect 1274 112 1276 114
rect 1280 112 1282 114
rect 1304 112 1306 114
rect 1356 112 1358 114
rect 1380 112 1382 114
rect 1386 112 1388 114
rect 1410 112 1412 114
rect 1416 112 1418 114
rect 1440 112 1442 114
rect 1446 112 1448 114
rect 1470 112 1472 114
rect 1476 112 1478 114
rect 1500 112 1502 114
rect 1162 110 1164 112
rect 1192 110 1194 112
rect 1222 110 1224 112
rect 1252 110 1254 112
rect 1282 110 1284 112
rect 1378 110 1380 112
rect 1408 110 1410 112
rect 1438 110 1440 112
rect 1468 110 1470 112
rect 1498 110 1500 112
rect 1162 104 1164 106
rect 1192 104 1194 106
rect 1222 104 1224 106
rect 1252 104 1254 106
rect 1282 104 1284 106
rect 1378 104 1380 106
rect 1408 104 1410 106
rect 1438 104 1440 106
rect 1468 104 1470 106
rect 1498 104 1500 106
rect 1160 102 1162 104
rect 1184 102 1186 104
rect 1190 102 1192 104
rect 1214 102 1216 104
rect 1220 102 1222 104
rect 1244 102 1246 104
rect 1250 102 1252 104
rect 1274 102 1276 104
rect 1280 102 1282 104
rect 1304 102 1306 104
rect 1356 102 1358 104
rect 1380 102 1382 104
rect 1386 102 1388 104
rect 1410 102 1412 104
rect 1416 102 1418 104
rect 1440 102 1442 104
rect 1446 102 1448 104
rect 1470 102 1472 104
rect 1476 102 1478 104
rect 1500 102 1502 104
rect 1182 100 1184 102
rect 1212 100 1214 102
rect 1242 100 1244 102
rect 1272 100 1274 102
rect 1302 100 1304 102
rect 1358 100 1360 102
rect 1388 100 1390 102
rect 1418 100 1420 102
rect 1448 100 1450 102
rect 1478 100 1480 102
rect 1182 94 1184 96
rect 1212 94 1214 96
rect 1242 94 1244 96
rect 1272 94 1274 96
rect 1302 94 1304 96
rect 1358 94 1360 96
rect 1388 94 1390 96
rect 1418 94 1420 96
rect 1448 94 1450 96
rect 1478 94 1480 96
rect 1160 92 1162 94
rect 1184 92 1186 94
rect 1190 92 1192 94
rect 1214 92 1216 94
rect 1220 92 1222 94
rect 1244 92 1246 94
rect 1250 92 1252 94
rect 1274 92 1276 94
rect 1280 92 1282 94
rect 1304 92 1306 94
rect 1356 92 1358 94
rect 1380 92 1382 94
rect 1386 92 1388 94
rect 1410 92 1412 94
rect 1416 92 1418 94
rect 1440 92 1442 94
rect 1446 92 1448 94
rect 1470 92 1472 94
rect 1476 92 1478 94
rect 1500 92 1502 94
rect 1162 90 1164 92
rect 1192 90 1194 92
rect 1222 90 1224 92
rect 1252 90 1254 92
rect 1282 90 1284 92
rect 1378 90 1380 92
rect 1408 90 1410 92
rect 1438 90 1440 92
rect 1468 90 1470 92
rect 1498 90 1500 92
rect 1162 84 1164 86
rect 1192 84 1194 86
rect 1222 84 1224 86
rect 1252 84 1254 86
rect 1282 84 1284 86
rect 1378 84 1380 86
rect 1408 84 1410 86
rect 1438 84 1440 86
rect 1468 84 1470 86
rect 1498 84 1500 86
rect 1160 82 1162 84
rect 1184 82 1186 84
rect 1190 82 1192 84
rect 1214 82 1216 84
rect 1220 82 1222 84
rect 1244 82 1246 84
rect 1250 82 1252 84
rect 1274 82 1276 84
rect 1280 82 1282 84
rect 1304 82 1306 84
rect 1356 82 1358 84
rect 1380 82 1382 84
rect 1386 82 1388 84
rect 1410 82 1412 84
rect 1416 82 1418 84
rect 1440 82 1442 84
rect 1446 82 1448 84
rect 1470 82 1472 84
rect 1476 82 1478 84
rect 1500 82 1502 84
rect 1182 80 1184 82
rect 1212 80 1214 82
rect 1242 80 1244 82
rect 1272 80 1274 82
rect 1302 80 1304 82
rect 1358 80 1360 82
rect 1388 80 1390 82
rect 1418 80 1420 82
rect 1448 80 1450 82
rect 1478 80 1480 82
rect 1182 74 1184 76
rect 1212 74 1214 76
rect 1242 74 1244 76
rect 1272 74 1274 76
rect 1302 74 1304 76
rect 1358 74 1360 76
rect 1388 74 1390 76
rect 1418 74 1420 76
rect 1448 74 1450 76
rect 1478 74 1480 76
rect 1160 72 1162 74
rect 1184 72 1186 74
rect 1190 72 1192 74
rect 1214 72 1216 74
rect 1220 72 1222 74
rect 1244 72 1246 74
rect 1250 72 1252 74
rect 1274 72 1276 74
rect 1280 72 1282 74
rect 1304 72 1306 74
rect 1356 72 1358 74
rect 1380 72 1382 74
rect 1386 72 1388 74
rect 1410 72 1412 74
rect 1416 72 1418 74
rect 1440 72 1442 74
rect 1446 72 1448 74
rect 1470 72 1472 74
rect 1476 72 1478 74
rect 1500 72 1502 74
rect 1162 70 1164 72
rect 1192 70 1194 72
rect 1222 70 1224 72
rect 1252 70 1254 72
rect 1282 70 1284 72
rect 1378 70 1380 72
rect 1408 70 1410 72
rect 1438 70 1440 72
rect 1468 70 1470 72
rect 1498 70 1500 72
rect 1162 64 1164 66
rect 1192 64 1194 66
rect 1222 64 1224 66
rect 1252 64 1254 66
rect 1282 64 1284 66
rect 1378 64 1380 66
rect 1408 64 1410 66
rect 1438 64 1440 66
rect 1468 64 1470 66
rect 1498 64 1500 66
rect 1160 62 1162 64
rect 1184 62 1186 64
rect 1190 62 1192 64
rect 1214 62 1216 64
rect 1220 62 1222 64
rect 1244 62 1246 64
rect 1250 62 1252 64
rect 1274 62 1276 64
rect 1280 62 1282 64
rect 1304 62 1306 64
rect 1356 62 1358 64
rect 1380 62 1382 64
rect 1386 62 1388 64
rect 1410 62 1412 64
rect 1416 62 1418 64
rect 1440 62 1442 64
rect 1446 62 1448 64
rect 1470 62 1472 64
rect 1476 62 1478 64
rect 1500 62 1502 64
rect 1182 60 1184 62
rect 1212 60 1214 62
rect 1242 60 1244 62
rect 1272 60 1274 62
rect 1302 60 1304 62
rect 1358 60 1360 62
rect 1388 60 1390 62
rect 1418 60 1420 62
rect 1448 60 1450 62
rect 1478 60 1480 62
rect 1182 54 1184 56
rect 1212 54 1214 56
rect 1242 54 1244 56
rect 1272 54 1274 56
rect 1302 54 1304 56
rect 1358 54 1360 56
rect 1388 54 1390 56
rect 1418 54 1420 56
rect 1448 54 1450 56
rect 1478 54 1480 56
rect 1160 52 1162 54
rect 1184 52 1186 54
rect 1190 52 1192 54
rect 1214 52 1216 54
rect 1220 52 1222 54
rect 1244 52 1246 54
rect 1250 52 1252 54
rect 1274 52 1276 54
rect 1280 52 1282 54
rect 1304 52 1306 54
rect 1356 52 1358 54
rect 1380 52 1382 54
rect 1386 52 1388 54
rect 1410 52 1412 54
rect 1416 52 1418 54
rect 1440 52 1442 54
rect 1446 52 1448 54
rect 1470 52 1472 54
rect 1476 52 1478 54
rect 1500 52 1502 54
rect 1162 50 1164 52
rect 1192 50 1194 52
rect 1222 50 1224 52
rect 1252 50 1254 52
rect 1282 50 1284 52
rect 1378 50 1380 52
rect 1408 50 1410 52
rect 1438 50 1440 52
rect 1468 50 1470 52
rect 1498 50 1500 52
rect 1162 44 1164 46
rect 1192 44 1194 46
rect 1222 44 1224 46
rect 1252 44 1254 46
rect 1282 44 1284 46
rect 1378 44 1380 46
rect 1408 44 1410 46
rect 1438 44 1440 46
rect 1468 44 1470 46
rect 1498 44 1500 46
rect 1160 42 1162 44
rect 1184 42 1186 44
rect 1190 42 1192 44
rect 1214 42 1216 44
rect 1220 42 1222 44
rect 1244 42 1246 44
rect 1250 42 1252 44
rect 1274 42 1276 44
rect 1280 42 1282 44
rect 1304 42 1306 44
rect 1356 42 1358 44
rect 1380 42 1382 44
rect 1386 42 1388 44
rect 1410 42 1412 44
rect 1416 42 1418 44
rect 1440 42 1442 44
rect 1446 42 1448 44
rect 1470 42 1472 44
rect 1476 42 1478 44
rect 1500 42 1502 44
rect 1182 40 1184 42
rect 1212 40 1214 42
rect 1242 40 1244 42
rect 1272 40 1274 42
rect 1302 40 1304 42
rect 1358 40 1360 42
rect 1388 40 1390 42
rect 1418 40 1420 42
rect 1448 40 1450 42
rect 1478 40 1480 42
rect 1182 34 1184 36
rect 1212 34 1214 36
rect 1242 34 1244 36
rect 1272 34 1274 36
rect 1302 34 1304 36
rect 1358 34 1360 36
rect 1388 34 1390 36
rect 1418 34 1420 36
rect 1448 34 1450 36
rect 1478 34 1480 36
rect 1160 32 1162 34
rect 1184 32 1186 34
rect 1190 32 1192 34
rect 1214 32 1216 34
rect 1220 32 1222 34
rect 1244 32 1246 34
rect 1250 32 1252 34
rect 1274 32 1276 34
rect 1280 32 1282 34
rect 1304 32 1306 34
rect 1356 32 1358 34
rect 1380 32 1382 34
rect 1386 32 1388 34
rect 1410 32 1412 34
rect 1416 32 1418 34
rect 1440 32 1442 34
rect 1446 32 1448 34
rect 1470 32 1472 34
rect 1476 32 1478 34
rect 1500 32 1502 34
rect 1162 30 1164 32
rect 1192 30 1194 32
rect 1222 30 1224 32
rect 1252 30 1254 32
rect 1282 30 1284 32
rect 1378 30 1380 32
rect 1408 30 1410 32
rect 1438 30 1440 32
rect 1468 30 1470 32
rect 1498 30 1500 32
rect 1162 24 1164 26
rect 1192 24 1194 26
rect 1222 24 1224 26
rect 1252 24 1254 26
rect 1282 24 1284 26
rect 1378 24 1380 26
rect 1408 24 1410 26
rect 1438 24 1440 26
rect 1468 24 1470 26
rect 1498 24 1500 26
rect 1160 22 1162 24
rect 1184 22 1186 24
rect 1190 22 1192 24
rect 1214 22 1216 24
rect 1220 22 1222 24
rect 1244 22 1246 24
rect 1250 22 1252 24
rect 1274 22 1276 24
rect 1280 22 1282 24
rect 1304 22 1306 24
rect 1356 22 1358 24
rect 1380 22 1382 24
rect 1386 22 1388 24
rect 1410 22 1412 24
rect 1416 22 1418 24
rect 1440 22 1442 24
rect 1446 22 1448 24
rect 1470 22 1472 24
rect 1476 22 1478 24
rect 1500 22 1502 24
rect 1182 20 1184 22
rect 1212 20 1214 22
rect 1242 20 1244 22
rect 1272 20 1274 22
rect 1302 20 1304 22
rect 1358 20 1360 22
rect 1388 20 1390 22
rect 1418 20 1420 22
rect 1448 20 1450 22
rect 1478 20 1480 22
rect 1182 14 1184 16
rect 1212 14 1214 16
rect 1242 14 1244 16
rect 1272 14 1274 16
rect 1302 14 1304 16
rect 1358 14 1360 16
rect 1388 14 1390 16
rect 1418 14 1420 16
rect 1448 14 1450 16
rect 1478 14 1480 16
rect 1160 12 1162 14
rect 1184 12 1186 14
rect 1190 12 1192 14
rect 1214 12 1216 14
rect 1220 12 1222 14
rect 1244 12 1246 14
rect 1250 12 1252 14
rect 1274 12 1276 14
rect 1280 12 1282 14
rect 1304 12 1306 14
rect 1356 12 1358 14
rect 1380 12 1382 14
rect 1386 12 1388 14
rect 1410 12 1412 14
rect 1416 12 1418 14
rect 1440 12 1442 14
rect 1446 12 1448 14
rect 1470 12 1472 14
rect 1476 12 1478 14
rect 1500 12 1502 14
rect 1162 10 1164 12
rect 1192 10 1194 12
rect 1222 10 1224 12
rect 1252 10 1254 12
rect 1282 10 1284 12
rect 1378 10 1380 12
rect 1408 10 1410 12
rect 1438 10 1440 12
rect 1468 10 1470 12
rect 1498 10 1500 12
<< nwell >>
tri 1340 182 1818 660 se
rect 1818 182 2006 660
rect 1340 -6 2006 182
<< psubstratepdiff >>
tri 1580 1338 1582 1340 se
rect 1582 1338 2000 1340
tri 1574 1332 1580 1338 se
rect 1580 1332 2000 1338
tri 1568 1326 1574 1332 se
rect 1574 1326 1584 1332
tri 1562 1320 1568 1326 se
rect 1568 1322 1584 1326
rect 1568 1320 1574 1322
tri 1556 1314 1562 1320 se
rect 1562 1314 1574 1320
tri 1550 1308 1556 1314 se
rect 1556 1312 1574 1314
rect 1556 1308 1564 1312
tri 1544 1302 1550 1308 se
rect 1550 1302 1564 1308
tri 1538 1296 1544 1302 se
rect 1544 1296 1554 1302
tri 1532 1290 1538 1296 se
rect 1538 1292 1554 1296
rect 1538 1290 1544 1292
tri 1528 1286 1532 1290 se
rect 1532 1286 1544 1290
tri 1522 1280 1528 1286 se
rect 1528 1282 1544 1286
rect 1528 1280 1534 1282
tri 1516 1274 1522 1280 se
rect 1522 1274 1534 1280
tri 1510 1268 1516 1274 se
rect 1516 1272 1534 1274
rect 1516 1268 1524 1272
tri 1504 1262 1510 1268 se
rect 1510 1262 1524 1268
tri 1498 1256 1504 1262 se
rect 1504 1256 1514 1262
tri 1492 1250 1498 1256 se
rect 1498 1252 1514 1256
rect 1498 1250 1504 1252
tri 1486 1244 1492 1250 se
rect 1492 1244 1504 1250
tri 1480 1238 1486 1244 se
rect 1486 1242 1504 1244
rect 1486 1238 1494 1242
tri 1474 1232 1480 1238 se
rect 1480 1232 1494 1238
tri 1468 1226 1474 1232 se
rect 1474 1226 1484 1232
tri 1462 1220 1468 1226 se
rect 1468 1222 1484 1226
rect 1468 1220 1474 1222
tri 1456 1214 1462 1220 se
rect 1462 1214 1474 1220
tri 1450 1208 1456 1214 se
rect 1456 1212 1474 1214
rect 1456 1208 1464 1212
tri 1444 1202 1450 1208 se
rect 1450 1202 1464 1208
tri 1438 1196 1444 1202 se
rect 1444 1196 1454 1202
tri 1432 1190 1438 1196 se
rect 1438 1192 1454 1196
rect 1438 1190 1444 1192
tri 1426 1184 1432 1190 se
rect 1432 1184 1444 1190
tri 1420 1178 1426 1184 se
rect 1426 1182 1444 1184
rect 1426 1178 1434 1182
tri 1414 1172 1420 1178 se
rect 1420 1172 1434 1178
tri 1408 1166 1414 1172 se
rect 1414 1166 1424 1172
tri 1402 1160 1408 1166 se
rect 1408 1162 1424 1166
rect 1408 1160 1414 1162
tri 1396 1154 1402 1160 se
rect 1402 1154 1414 1160
tri 1390 1148 1396 1154 se
rect 1396 1152 1414 1154
rect 1396 1148 1404 1152
tri 1384 1142 1390 1148 se
rect 1390 1142 1404 1148
tri 1378 1136 1384 1142 se
rect 1384 1136 1394 1142
tri 1372 1130 1378 1136 se
rect 1378 1132 1394 1136
rect 1378 1130 1384 1132
tri 1366 1124 1372 1130 se
rect 1372 1124 1384 1130
tri 1360 1118 1366 1124 se
rect 1366 1122 1384 1124
rect 1366 1118 1374 1122
tri 1354 1112 1360 1118 se
rect 1360 1112 1374 1118
tri 1348 1106 1354 1112 se
rect 1354 1106 1364 1112
tri 1342 1100 1348 1106 se
rect 1348 1102 1364 1106
rect 1348 1100 1354 1102
tri 1336 1094 1342 1100 se
rect 1342 1094 1354 1100
tri 1330 1088 1336 1094 se
rect 1336 1092 1354 1094
rect 1336 1088 1344 1092
tri 1324 1082 1330 1088 se
rect 1330 1082 1344 1088
tri 1318 1076 1324 1082 se
rect 1324 1076 1334 1082
tri 1312 1070 1318 1076 se
rect 1318 1072 1334 1076
rect 1318 1070 1324 1072
tri 1306 1064 1312 1070 se
rect 1312 1064 1324 1070
tri 1300 1058 1306 1064 se
rect 1306 1062 1324 1064
rect 1306 1058 1314 1062
tri 1294 1052 1300 1058 se
rect 1300 1052 1314 1058
tri 1288 1046 1294 1052 se
rect 1294 1046 1304 1052
tri 1282 1040 1288 1046 se
rect 1288 1042 1304 1046
rect 1572 1044 1594 1054
rect 1288 1040 1294 1042
tri 1276 1034 1282 1040 se
rect 1282 1034 1294 1040
rect 1562 1034 1594 1044
tri 1270 1028 1276 1034 se
rect 1276 1032 1294 1034
rect 1276 1028 1284 1032
tri 1264 1022 1270 1028 se
rect 1270 1022 1284 1028
rect 1552 1024 1594 1034
rect 1542 1022 1594 1024
tri 1258 1016 1264 1022 se
rect 1264 1016 1274 1022
tri 1252 1010 1258 1016 se
rect 1258 1012 1274 1016
rect 1542 1014 1584 1022
rect 1532 1012 1584 1014
rect 1258 1010 1264 1012
tri 1246 1004 1252 1010 se
rect 1252 1004 1264 1010
rect 1532 1004 1574 1012
tri 1240 998 1246 1004 se
rect 1246 1002 1264 1004
rect 1522 1002 1574 1004
rect 1246 998 1254 1002
tri 1234 992 1240 998 se
rect 1240 992 1254 998
rect 1522 994 1564 1002
rect 1512 992 1564 994
tri 1228 986 1234 992 se
rect 1234 986 1244 992
tri 1222 980 1228 986 se
rect 1228 982 1244 986
rect 1512 984 1554 992
rect 1502 982 1554 984
rect 1228 980 1234 982
tri 1216 974 1222 980 se
rect 1222 974 1234 980
rect 1502 974 1544 982
tri 1210 968 1216 974 se
rect 1216 972 1234 974
rect 1492 972 1544 974
rect 1216 968 1224 972
tri 1208 966 1210 968 se
rect 1210 966 1224 968
tri 1202 960 1208 966 se
rect 1208 962 1224 966
rect 1492 964 1534 972
rect 1482 962 1534 964
rect 1208 960 1214 962
tri 1196 954 1202 960 se
rect 1202 954 1214 960
rect 1482 954 1524 962
tri 1190 948 1196 954 se
rect 1196 952 1214 954
rect 1472 952 1524 954
rect 1196 948 1204 952
tri 1184 942 1190 948 se
rect 1190 942 1204 948
rect 1472 944 1514 952
rect 1462 942 1514 944
tri 1178 936 1184 942 se
rect 1184 936 1194 942
tri 1172 930 1178 936 se
rect 1178 932 1194 936
rect 1462 934 1504 942
rect 1452 932 1504 934
rect 1178 930 1184 932
tri 1166 924 1172 930 se
rect 1172 924 1184 930
rect 1452 924 1494 932
tri 1160 918 1166 924 se
rect 1166 922 1184 924
rect 1442 922 1494 924
rect 1166 918 1174 922
tri 1154 912 1160 918 se
rect 1160 912 1174 918
rect 1442 914 1484 922
rect 1432 912 1484 914
tri 1148 906 1154 912 se
rect 1154 906 1164 912
tri 1142 900 1148 906 se
rect 1148 902 1164 906
rect 1432 904 1474 912
rect 1422 902 1474 904
rect 1148 900 1154 902
tri 1136 894 1142 900 se
rect 1142 894 1154 900
rect 1422 894 1464 902
tri 1130 888 1136 894 se
rect 1136 892 1154 894
rect 1412 892 1464 894
rect 1136 888 1144 892
tri 1124 882 1130 888 se
rect 1130 882 1144 888
rect 1412 884 1454 892
rect 1402 882 1454 884
tri 1118 876 1124 882 se
rect 1124 876 1134 882
tri 1112 870 1118 876 se
rect 1118 872 1134 876
rect 1402 874 1444 882
rect 1702 874 1734 884
rect 1392 872 1444 874
rect 1118 870 1124 872
tri 1106 864 1112 870 se
rect 1112 864 1124 870
rect 1392 864 1434 872
rect 1692 864 1734 874
tri 1100 858 1106 864 se
rect 1106 862 1124 864
rect 1382 862 1434 864
rect 1682 862 1734 864
rect 1106 858 1114 862
tri 1094 852 1100 858 se
rect 1100 852 1114 858
rect 1382 854 1424 862
rect 1682 854 1724 862
rect 1372 852 1424 854
rect 1672 852 1724 854
tri 1088 846 1094 852 se
rect 1094 846 1104 852
tri 1082 840 1088 846 se
rect 1088 842 1104 846
rect 1372 844 1414 852
rect 1672 844 1714 852
rect 1362 842 1414 844
rect 1662 842 1714 844
rect 1088 840 1094 842
tri 1076 834 1082 840 se
rect 1082 834 1094 840
rect 1362 834 1404 842
rect 1662 834 1704 842
tri 1070 828 1076 834 se
rect 1076 832 1094 834
rect 1352 832 1404 834
rect 1652 832 1704 834
rect 1722 834 1734 844
rect 1752 834 1764 844
rect 1782 834 1794 844
rect 1812 834 1824 844
rect 1842 834 1854 844
rect 1872 834 1884 844
rect 1902 834 1914 844
rect 1932 834 1944 844
rect 1962 834 1974 844
rect 1722 832 1744 834
rect 1752 832 1774 834
rect 1782 832 1804 834
rect 1812 832 1834 834
rect 1842 832 1864 834
rect 1872 832 1894 834
rect 1902 832 1924 834
rect 1932 832 1954 834
rect 1962 832 1984 834
rect 1076 828 1084 832
tri 1064 822 1070 828 se
rect 1070 822 1084 828
rect 1352 824 1394 832
rect 1652 824 1694 832
rect 1732 824 1744 832
rect 1762 824 1774 832
rect 1792 824 1804 832
rect 1822 824 1834 832
rect 1852 824 1864 832
rect 1882 824 1894 832
rect 1912 824 1924 832
rect 1942 824 1954 832
rect 1972 824 1984 832
rect 1342 822 1394 824
rect 1642 822 1694 824
rect 1722 822 1744 824
rect 1752 822 1774 824
rect 1782 822 1804 824
rect 1812 822 1834 824
rect 1842 822 1864 824
rect 1872 822 1894 824
rect 1902 822 1924 824
rect 1932 822 1954 824
rect 1962 822 1984 824
tri 1058 816 1064 822 se
rect 1064 816 1074 822
tri 1052 810 1058 816 se
rect 1058 812 1074 816
rect 1342 814 1384 822
rect 1642 814 1684 822
rect 1722 814 1734 822
rect 1752 814 1764 822
rect 1782 814 1794 822
rect 1812 814 1824 822
rect 1842 814 1854 822
rect 1872 814 1884 822
rect 1902 814 1914 822
rect 1932 814 1944 822
rect 1962 814 1974 822
rect 1332 812 1384 814
rect 1632 812 1684 814
rect 1058 810 1064 812
tri 1046 804 1052 810 se
rect 1052 804 1064 810
rect 1332 804 1374 812
rect 1632 804 1674 812
rect 1692 804 1704 814
rect 1722 812 1744 814
rect 1752 812 1774 814
rect 1782 812 1804 814
rect 1812 812 1834 814
rect 1842 812 1864 814
rect 1872 812 1894 814
rect 1902 812 1924 814
rect 1932 812 1954 814
rect 1962 812 1984 814
rect 1732 804 1744 812
rect 1762 804 1774 812
rect 1792 804 1804 812
rect 1822 804 1834 812
rect 1852 804 1864 812
rect 1882 804 1894 812
rect 1912 804 1924 812
rect 1942 804 1954 812
rect 1972 804 1984 812
tri 1040 798 1046 804 se
rect 1046 802 1064 804
rect 1322 802 1374 804
rect 1622 802 1674 804
rect 1682 802 1704 804
rect 1722 802 1744 804
rect 1752 802 1774 804
rect 1782 802 1804 804
rect 1812 802 1834 804
rect 1842 802 1864 804
rect 1872 802 1894 804
rect 1902 802 1924 804
rect 1932 802 1954 804
rect 1962 802 1984 804
rect 1046 798 1054 802
tri 1034 792 1040 798 se
rect 1040 792 1054 798
rect 1322 794 1364 802
rect 1622 794 1664 802
rect 1682 794 1694 802
rect 1722 794 1734 802
rect 1752 794 1764 802
rect 1782 794 1794 802
rect 1812 794 1824 802
rect 1842 794 1854 802
rect 1872 794 1884 802
rect 1902 794 1914 802
rect 1932 794 1944 802
rect 1962 794 1974 802
rect 1312 792 1364 794
rect 1612 792 1664 794
rect 1672 792 1704 794
rect 1722 792 1744 794
rect 1752 792 1774 794
rect 1782 792 1804 794
rect 1812 792 1834 794
rect 1842 792 1864 794
rect 1872 792 1894 794
rect 1902 792 1924 794
rect 1932 792 1954 794
rect 1962 792 1984 794
tri 1028 786 1034 792 se
rect 1034 786 1044 792
tri 1022 780 1028 786 se
rect 1028 782 1044 786
rect 1312 784 1354 792
rect 1612 784 1654 792
rect 1672 784 1684 792
rect 1692 784 1704 792
rect 1732 784 1744 792
rect 1762 784 1774 792
rect 1792 784 1804 792
rect 1822 784 1834 792
rect 1852 784 1864 792
rect 1882 784 1894 792
rect 1912 784 1924 792
rect 1942 784 1954 792
rect 1972 784 1984 792
rect 1302 782 1354 784
rect 1602 782 1654 784
rect 1662 782 1704 784
rect 1722 782 1744 784
rect 1752 782 1774 784
rect 1782 782 1804 784
rect 1812 782 1834 784
rect 1842 782 1864 784
rect 1872 782 1894 784
rect 1902 782 1924 784
rect 1932 782 1954 784
rect 1962 782 1984 784
rect 1028 780 1034 782
tri 1016 774 1022 780 se
rect 1022 774 1034 780
rect 1302 774 1344 782
rect 1602 774 1644 782
rect 1662 774 1674 782
rect 1682 774 1694 782
tri 1010 768 1016 774 se
rect 1016 772 1034 774
rect 1292 772 1344 774
rect 1592 772 1644 774
rect 1652 772 1694 774
rect 1722 774 1734 782
rect 1752 774 1764 782
rect 1782 774 1794 782
rect 1812 774 1824 782
rect 1842 774 1854 782
rect 1872 774 1884 782
rect 1902 774 1914 782
rect 1932 774 1944 782
rect 1962 774 1974 782
rect 1722 772 1744 774
rect 1752 772 1774 774
rect 1782 772 1804 774
rect 1812 772 1834 774
rect 1842 772 1864 774
rect 1872 772 1894 774
rect 1902 772 1924 774
rect 1932 772 1954 774
rect 1962 772 1984 774
rect 1016 768 1024 772
tri 1004 762 1010 768 se
rect 1010 762 1024 768
rect 1292 764 1334 772
rect 1592 764 1634 772
rect 1652 764 1664 772
rect 1672 764 1684 772
rect 1732 764 1744 772
rect 1762 764 1774 772
rect 1792 764 1804 772
rect 1822 764 1834 772
rect 1852 764 1864 772
rect 1882 764 1894 772
rect 1912 764 1924 772
rect 1942 764 1954 772
rect 1972 764 1984 772
rect 1282 762 1334 764
rect 1582 762 1634 764
rect 1642 762 1684 764
tri 998 756 1004 762 se
rect 1004 756 1014 762
tri 992 750 998 756 se
rect 998 752 1014 756
rect 1282 754 1324 762
rect 1582 754 1624 762
rect 1642 754 1654 762
rect 1662 754 1674 762
rect 1692 754 1704 764
rect 1272 752 1324 754
rect 1572 752 1624 754
rect 1632 752 1674 754
rect 1682 752 1704 754
rect 1722 762 1744 764
rect 1752 762 1774 764
rect 1782 762 1804 764
rect 1812 762 1834 764
rect 1842 762 1864 764
rect 1872 762 1894 764
rect 1902 762 1924 764
rect 1932 762 1954 764
rect 1962 762 1984 764
rect 1722 754 1734 762
rect 1752 754 1764 762
rect 1782 754 1794 762
rect 1812 754 1824 762
rect 1842 754 1854 762
rect 1872 754 1884 762
rect 1902 754 1914 762
rect 1932 754 1944 762
rect 1962 754 1974 762
rect 1722 752 1744 754
rect 1752 752 1774 754
rect 1782 752 1804 754
rect 1812 752 1834 754
rect 1842 752 1864 754
rect 1872 752 1894 754
rect 1902 752 1924 754
rect 1932 752 1954 754
rect 1962 752 1984 754
rect 998 750 1004 752
tri 986 744 992 750 se
rect 992 744 1004 750
rect 1272 744 1314 752
rect 1572 744 1614 752
rect 1632 744 1644 752
rect 1652 744 1664 752
rect 1682 744 1694 752
rect 1732 744 1744 752
rect 1762 744 1774 752
rect 1792 744 1804 752
rect 1822 744 1834 752
rect 1852 744 1864 752
rect 1882 744 1894 752
rect 1912 744 1924 752
rect 1942 744 1954 752
rect 1972 744 1984 752
tri 980 738 986 744 se
rect 986 742 1004 744
rect 1262 742 1314 744
rect 1562 742 1614 744
rect 1622 742 1664 744
rect 1672 742 1694 744
rect 1722 742 1744 744
rect 1752 742 1774 744
rect 1782 742 1804 744
rect 1812 742 1834 744
rect 1842 742 1864 744
rect 1872 742 1894 744
rect 1902 742 1924 744
rect 1932 742 1954 744
rect 1962 742 1984 744
rect 986 738 994 742
tri 974 732 980 738 se
rect 980 732 994 738
rect 1262 734 1304 742
rect 1562 734 1604 742
rect 1622 734 1634 742
rect 1642 734 1654 742
rect 1672 734 1684 742
rect 1252 732 1304 734
rect 1552 732 1604 734
rect 1612 732 1654 734
rect 1662 732 1684 734
rect 1722 734 1734 742
rect 1752 734 1764 742
rect 1782 734 1794 742
rect 1812 734 1824 742
rect 1842 734 1854 742
rect 1872 734 1884 742
rect 1902 734 1914 742
rect 1932 734 1944 742
rect 1962 734 1974 742
rect 1722 732 1744 734
rect 1752 732 1774 734
rect 1782 732 1804 734
rect 1812 732 1834 734
rect 1842 732 1864 734
rect 1872 732 1894 734
rect 1902 732 1924 734
rect 1932 732 1954 734
rect 1962 732 1984 734
tri 968 726 974 732 se
rect 974 726 984 732
tri 962 720 968 726 se
rect 968 722 984 726
rect 1252 724 1294 732
rect 1552 724 1594 732
rect 1612 724 1624 732
rect 1632 724 1644 732
rect 1662 724 1674 732
rect 1732 724 1744 732
rect 1762 724 1774 732
rect 1792 724 1804 732
rect 1822 724 1834 732
rect 1852 724 1864 732
rect 1882 724 1894 732
rect 1912 724 1924 732
rect 1942 724 1954 732
rect 1972 724 1984 732
rect 1242 722 1294 724
rect 1542 722 1594 724
rect 1602 722 1644 724
rect 1652 722 1674 724
rect 1722 722 1744 724
rect 1752 722 1774 724
rect 1782 722 1804 724
rect 1812 722 1834 724
rect 1842 722 1864 724
rect 1872 722 1894 724
rect 1902 722 1924 724
rect 1932 722 1954 724
rect 1962 722 1984 724
rect 968 720 974 722
tri 956 714 962 720 se
rect 962 714 974 720
rect 1242 714 1284 722
rect 1542 714 1584 722
rect 1602 714 1614 722
rect 1622 714 1634 722
rect 1652 714 1664 722
tri 950 708 956 714 se
rect 956 712 974 714
rect 1232 712 1284 714
rect 1532 712 1584 714
rect 1592 712 1634 714
rect 1642 712 1664 714
rect 1722 714 1734 722
rect 1752 714 1764 722
rect 1782 714 1794 722
rect 1812 714 1824 722
rect 1842 714 1854 722
rect 1872 714 1884 722
rect 1902 714 1914 722
rect 1932 714 1944 722
rect 1962 714 1974 722
rect 1722 712 1744 714
rect 1752 712 1774 714
rect 1782 712 1804 714
rect 1812 712 1834 714
rect 1842 712 1864 714
rect 1872 712 1894 714
rect 1902 712 1924 714
rect 1932 712 1954 714
rect 1962 712 1984 714
rect 956 708 964 712
tri 944 702 950 708 se
rect 950 702 964 708
rect 1232 704 1274 712
rect 1532 704 1574 712
rect 1592 704 1604 712
rect 1612 704 1624 712
rect 1642 704 1654 712
rect 1732 704 1744 712
rect 1762 704 1774 712
rect 1792 704 1804 712
rect 1822 704 1834 712
rect 1852 704 1864 712
rect 1882 704 1894 712
rect 1912 704 1924 712
rect 1942 704 1954 712
rect 1972 704 1984 712
rect 1222 702 1274 704
rect 1522 702 1574 704
rect 1582 702 1624 704
rect 1632 702 1654 704
tri 938 696 944 702 se
rect 944 696 954 702
tri 932 690 938 696 se
rect 938 692 954 696
rect 1222 694 1264 702
rect 1522 694 1564 702
rect 1582 694 1594 702
rect 1602 694 1614 702
rect 1212 692 1264 694
rect 1512 692 1564 694
rect 1572 692 1624 694
rect 938 690 944 692
tri 926 684 932 690 se
rect 932 684 944 690
rect 1212 684 1254 692
rect 1512 684 1554 692
rect 1572 684 1584 692
rect 1592 684 1604 692
rect 1612 684 1624 692
rect 1632 684 1644 702
rect 1692 694 1704 704
rect 1722 702 1744 704
rect 1752 702 1774 704
rect 1782 702 1804 704
rect 1812 702 1834 704
rect 1842 702 1864 704
rect 1872 702 1894 704
rect 1902 702 1924 704
rect 1932 702 1954 704
rect 1962 702 1984 704
rect 1682 692 1714 694
rect 1682 684 1694 692
rect 1702 684 1714 692
rect 1722 684 1734 702
rect 1752 694 1764 702
rect 1782 694 1794 702
rect 1812 694 1824 702
rect 1842 694 1854 702
rect 1872 694 1884 702
rect 1902 694 1914 702
rect 1932 694 1944 702
rect 1962 694 1974 702
rect 1992 694 2000 1332
rect 1742 692 1774 694
rect 1742 684 1754 692
rect 1762 684 1774 692
rect 1782 686 2000 694
rect 1782 684 1784 686
tri 920 678 926 684 se
rect 926 682 944 684
rect 1202 682 1254 684
rect 1502 682 1554 684
rect 1562 682 1644 684
rect 1672 682 1784 684
rect 926 678 934 682
tri 914 672 920 678 se
rect 920 672 934 678
rect 1202 674 1244 682
rect 1502 674 1544 682
rect 1562 674 1574 682
rect 1582 674 1594 682
rect 1602 674 1614 682
rect 1622 674 1634 682
rect 1672 674 1684 682
rect 1692 674 1704 682
rect 1712 674 1724 682
rect 1732 674 1744 682
rect 1752 674 1764 682
rect 1772 680 1784 682
tri 1784 680 1790 686 nw
rect 1772 674 1776 680
rect 1192 672 1244 674
rect 1492 672 1544 674
rect 1552 672 1634 674
rect 1662 672 1776 674
tri 1776 672 1784 680 nw
tri 908 666 914 672 se
rect 914 666 924 672
tri 902 660 908 666 se
rect 908 662 924 666
rect 1192 664 1234 672
rect 1492 664 1534 672
rect 1552 664 1564 672
rect 1572 664 1584 672
rect 1592 664 1604 672
rect 1612 664 1624 672
rect 1662 664 1674 672
rect 1682 664 1694 672
rect 1702 664 1714 672
rect 1722 664 1734 672
rect 1742 664 1754 672
rect 1762 664 1768 672
tri 1768 664 1776 672 nw
rect 1182 662 1234 664
rect 1482 662 1534 664
rect 1542 662 1624 664
rect 1652 662 1766 664
tri 1766 662 1768 664 nw
rect 908 660 914 662
tri 896 654 902 660 se
rect 902 654 914 660
rect 1182 654 1224 662
rect 1482 654 1524 662
rect 1542 654 1554 662
rect 1562 654 1574 662
rect 1582 654 1594 662
rect 1602 654 1614 662
rect 1652 654 1664 662
rect 1672 654 1684 662
rect 1692 654 1704 662
rect 1712 654 1724 662
rect 1732 654 1744 662
rect 1752 660 1764 662
tri 1764 660 1766 662 nw
rect 1752 658 1762 660
tri 1762 658 1764 660 nw
rect 1752 654 1758 658
tri 1758 654 1762 658 nw
tri 894 652 896 654 se
rect 896 652 914 654
rect 1172 652 1224 654
rect 1472 652 1524 654
rect 1532 652 1614 654
rect 1642 652 1756 654
tri 1756 652 1758 654 nw
tri 892 650 894 652 se
rect 894 650 904 652
tri 890 648 892 650 se
rect 892 648 904 650
tri 888 646 890 648 se
rect 890 646 904 648
tri 884 642 888 646 se
rect 888 642 904 646
rect 1172 644 1214 652
rect 1472 644 1514 652
rect 1532 644 1544 652
rect 1552 644 1564 652
rect 1572 644 1584 652
rect 1592 644 1604 652
rect 1642 644 1654 652
rect 1662 644 1674 652
rect 1682 644 1694 652
rect 1702 644 1714 652
rect 1722 644 1734 652
rect 1742 650 1754 652
tri 1754 650 1756 652 nw
rect 1742 646 1750 650
tri 1750 646 1754 650 nw
rect 1742 644 1744 646
rect 1162 642 1214 644
rect 1462 642 1514 644
rect 1522 642 1604 644
rect 1632 642 1744 644
tri 882 640 884 642 se
rect 884 640 894 642
tri 878 636 882 640 se
rect 882 636 894 640
tri 876 634 878 636 se
rect 878 634 894 636
rect 1162 634 1204 642
rect 1462 634 1504 642
rect 1522 634 1534 642
rect 1542 634 1554 642
rect 1562 634 1574 642
rect 1582 634 1594 642
rect 1632 634 1644 642
rect 1652 634 1664 642
rect 1672 634 1684 642
rect 1692 634 1704 642
rect 1712 634 1724 642
rect 1732 640 1744 642
tri 1744 640 1750 646 nw
rect 1732 638 1742 640
tri 1742 638 1744 640 nw
rect 1732 634 1738 638
tri 1738 634 1742 638 nw
tri 872 630 876 634 se
rect 876 632 894 634
rect 1152 632 1204 634
rect 1452 632 1504 634
rect 1512 632 1594 634
rect 1622 632 1734 634
rect 876 630 884 632
tri 870 628 872 630 se
rect 872 628 884 630
tri 866 624 870 628 se
rect 870 624 884 628
rect 1152 624 1194 632
rect 1452 624 1494 632
rect 1512 624 1524 632
rect 1532 624 1544 632
rect 1552 624 1564 632
rect 1572 624 1584 632
rect 1622 624 1634 632
rect 1642 624 1654 632
rect 1662 624 1674 632
rect 1682 624 1694 632
rect 1702 624 1714 632
rect 1722 630 1734 632
tri 1734 630 1738 634 nw
rect 1722 628 1732 630
tri 1732 628 1734 630 nw
rect 1722 624 1728 628
tri 1728 624 1732 628 nw
tri 864 622 866 624 se
rect 866 622 884 624
rect 1142 622 1194 624
rect 1442 622 1494 624
rect 1502 622 1584 624
rect 1612 622 1726 624
tri 1726 622 1728 624 nw
tri 860 618 864 622 se
rect 864 618 874 622
tri 858 616 860 618 se
rect 860 616 874 618
tri 854 612 858 616 se
rect 858 612 874 616
rect 1142 614 1184 622
rect 1442 614 1484 622
rect 1502 614 1514 622
rect 1522 614 1534 622
rect 1542 614 1554 622
rect 1562 614 1574 622
rect 1612 614 1624 622
rect 1632 614 1644 622
rect 1652 614 1664 622
rect 1672 614 1684 622
rect 1692 614 1704 622
rect 1712 616 1720 622
tri 1720 616 1726 622 nw
rect 1712 614 1718 616
tri 1718 614 1720 616 nw
rect 1132 612 1184 614
rect 1432 612 1484 614
rect 1492 612 1574 614
rect 1602 612 1714 614
tri 852 610 854 612 se
rect 854 610 864 612
tri 848 606 852 610 se
rect 852 606 864 610
tri 846 604 848 606 se
rect 848 604 864 606
rect 1132 604 1174 612
rect 1432 604 1474 612
rect 1492 604 1504 612
rect 1512 604 1524 612
rect 1532 604 1544 612
rect 1552 604 1564 612
rect 1602 604 1614 612
rect 1622 604 1634 612
rect 1642 604 1654 612
rect 1662 604 1674 612
rect 1682 604 1694 612
rect 1702 610 1714 612
tri 1714 610 1718 614 nw
rect 1702 606 1710 610
tri 1710 606 1714 610 nw
rect 1702 604 1708 606
tri 1708 604 1710 606 nw
tri 842 600 846 604 se
rect 846 602 864 604
rect 1122 602 1174 604
rect 1422 602 1474 604
rect 1482 602 1564 604
rect 1592 602 1702 604
rect 846 600 854 602
tri 840 598 842 600 se
rect 842 598 854 600
tri 836 594 840 598 se
rect 840 594 854 598
rect 1122 594 1164 602
rect 1422 594 1464 602
rect 1482 594 1494 602
rect 1502 594 1514 602
rect 1522 594 1534 602
rect 1542 594 1554 602
rect 1592 594 1604 602
rect 1612 594 1624 602
rect 1632 594 1644 602
rect 1652 594 1664 602
rect 1672 594 1684 602
rect 1692 598 1702 602
tri 1702 598 1708 604 nw
rect 1692 594 1696 598
tri 834 592 836 594 se
rect 836 592 854 594
rect 1112 592 1164 594
rect 1412 592 1464 594
rect 1472 592 1554 594
rect 1582 592 1696 594
tri 1696 592 1702 598 nw
tri 830 588 834 592 se
rect 834 588 844 592
tri 824 582 830 588 se
rect 830 582 844 588
rect 1112 584 1154 592
rect 1412 584 1454 592
rect 1472 584 1484 592
rect 1492 584 1504 592
rect 1512 584 1524 592
rect 1532 584 1544 592
rect 1582 584 1594 592
rect 1602 584 1614 592
rect 1622 584 1634 592
rect 1642 584 1654 592
rect 1662 584 1674 592
rect 1682 590 1694 592
tri 1694 590 1696 592 nw
rect 1682 588 1692 590
tri 1692 588 1694 590 nw
rect 1682 584 1686 588
rect 1102 582 1154 584
rect 1402 582 1454 584
rect 1462 582 1544 584
rect 1572 582 1686 584
tri 1686 582 1692 588 nw
tri 818 576 824 582 se
rect 824 576 834 582
tri 812 570 818 576 se
rect 818 572 834 576
rect 1102 574 1144 582
rect 1402 574 1444 582
rect 1462 574 1474 582
rect 1482 574 1494 582
rect 1502 574 1514 582
rect 1522 574 1534 582
rect 1572 574 1584 582
rect 1592 574 1604 582
rect 1612 574 1624 582
rect 1632 574 1644 582
rect 1652 574 1664 582
rect 1672 576 1680 582
tri 1680 576 1686 582 nw
rect 1672 574 1678 576
tri 1678 574 1680 576 nw
rect 1092 572 1144 574
rect 1392 572 1444 574
rect 1452 572 1534 574
rect 1562 572 1674 574
rect 818 570 824 572
tri 806 564 812 570 se
rect 812 564 824 570
rect 1092 564 1134 572
rect 1392 564 1434 572
rect 1452 564 1464 572
rect 1472 564 1484 572
rect 1492 564 1504 572
rect 1512 564 1524 572
rect 1562 564 1574 572
rect 1582 564 1594 572
rect 1602 564 1614 572
rect 1622 564 1634 572
rect 1642 564 1654 572
rect 1662 570 1674 572
tri 1674 570 1678 574 nw
rect 1662 566 1670 570
tri 1670 566 1674 570 nw
rect 1662 564 1668 566
tri 1668 564 1670 566 nw
tri 800 558 806 564 se
rect 806 562 824 564
rect 1082 562 1134 564
rect 1382 562 1434 564
rect 1442 562 1524 564
rect 1552 562 1662 564
rect 806 558 814 562
tri 794 552 800 558 se
rect 800 552 814 558
rect 1082 554 1124 562
rect 1382 554 1424 562
rect 1442 554 1454 562
rect 1462 554 1474 562
rect 1482 554 1494 562
rect 1502 554 1514 562
rect 1552 554 1564 562
rect 1572 554 1584 562
rect 1592 554 1604 562
rect 1612 554 1624 562
rect 1632 554 1644 562
rect 1652 558 1662 562
tri 1662 558 1668 564 nw
rect 1652 554 1656 558
rect 1072 552 1124 554
rect 1372 552 1424 554
rect 1432 552 1514 554
rect 1542 552 1656 554
tri 1656 552 1662 558 nw
tri 788 546 794 552 se
rect 794 546 804 552
tri 782 540 788 546 se
rect 788 542 804 546
rect 1072 544 1114 552
rect 1372 544 1414 552
rect 1432 544 1444 552
rect 1452 544 1464 552
rect 1472 544 1484 552
rect 1492 544 1504 552
rect 1542 544 1554 552
rect 1562 544 1574 552
rect 1582 544 1594 552
rect 1602 544 1614 552
rect 1622 544 1634 552
rect 1642 550 1654 552
tri 1654 550 1656 552 nw
rect 1642 546 1650 550
tri 1650 546 1654 550 nw
rect 1642 544 1644 546
rect 1062 542 1114 544
rect 1362 542 1414 544
rect 1422 542 1504 544
rect 1532 542 1644 544
rect 788 540 794 542
tri 776 534 782 540 se
rect 782 534 794 540
rect 1062 534 1104 542
rect 1362 534 1404 542
rect 1422 534 1434 542
rect 1442 534 1454 542
rect 1462 534 1474 542
rect 1482 534 1494 542
rect 1532 534 1544 542
rect 1552 534 1564 542
rect 1572 534 1584 542
rect 1592 534 1604 542
rect 1612 534 1624 542
rect 1632 540 1644 542
tri 1644 540 1650 546 nw
rect 1632 538 1642 540
tri 1642 538 1644 540 nw
rect 1632 534 1638 538
tri 1638 534 1642 538 nw
tri 770 528 776 534 se
rect 776 532 794 534
rect 1052 532 1104 534
rect 1352 532 1404 534
rect 1412 532 1494 534
rect 1522 532 1634 534
rect 776 528 784 532
tri 764 522 770 528 se
rect 770 522 784 528
rect 1052 524 1094 532
rect 1352 524 1394 532
rect 1412 524 1424 532
rect 1432 524 1444 532
rect 1452 524 1464 532
rect 1472 524 1484 532
rect 1522 524 1534 532
rect 1542 524 1554 532
rect 1562 524 1574 532
rect 1582 524 1594 532
rect 1602 524 1614 532
rect 1622 530 1634 532
tri 1634 530 1638 534 nw
rect 1622 528 1632 530
tri 1632 528 1634 530 nw
rect 1622 524 1626 528
rect 1042 522 1094 524
rect 1342 522 1394 524
rect 1402 522 1484 524
rect 1512 522 1626 524
tri 1626 522 1632 528 nw
tri 758 516 764 522 se
rect 764 516 774 522
tri 754 512 758 516 se
rect 758 512 774 516
rect 1042 514 1084 522
rect 1342 514 1384 522
rect 1402 514 1414 522
rect 1422 514 1434 522
rect 1442 514 1454 522
rect 1462 514 1474 522
rect 1512 514 1524 522
rect 1532 514 1544 522
rect 1552 514 1564 522
rect 1572 514 1584 522
rect 1592 514 1604 522
rect 1612 516 1620 522
tri 1620 516 1626 522 nw
rect 1612 514 1618 516
tri 1618 514 1620 516 nw
rect 1032 512 1084 514
rect 1332 512 1384 514
rect 1392 512 1474 514
rect 1502 512 1616 514
tri 1616 512 1618 514 nw
tri 752 510 754 512 se
rect 754 510 764 512
tri 748 506 752 510 se
rect 752 506 764 510
tri 746 504 748 506 se
rect 748 504 764 506
rect 1032 504 1074 512
rect 1332 504 1374 512
rect 1392 504 1404 512
rect 1412 504 1424 512
rect 1432 504 1444 512
rect 1452 504 1464 512
rect 1502 504 1514 512
rect 1522 504 1534 512
rect 1542 504 1554 512
rect 1562 504 1574 512
rect 1582 504 1594 512
rect 1602 506 1610 512
tri 1610 506 1616 512 nw
rect 1602 504 1604 506
tri 742 500 746 504 se
rect 746 502 764 504
rect 1022 502 1074 504
rect 1322 502 1374 504
rect 1382 502 1464 504
rect 1492 502 1604 504
rect 746 500 754 502
tri 740 498 742 500 se
rect 742 498 754 500
tri 736 494 740 498 se
rect 740 494 754 498
rect 1022 494 1064 502
rect 1322 494 1364 502
rect 1382 494 1394 502
rect 1402 494 1414 502
rect 1422 494 1434 502
rect 1442 494 1454 502
rect 1492 494 1504 502
rect 1512 494 1524 502
rect 1532 494 1544 502
rect 1552 494 1564 502
rect 1572 494 1584 502
rect 1592 500 1604 502
tri 1604 500 1610 506 nw
rect 1592 498 1602 500
tri 1602 498 1604 500 nw
rect 1592 494 1598 498
tri 1598 494 1602 498 nw
tri 734 492 736 494 se
rect 736 492 754 494
rect 1012 492 1064 494
rect 1312 492 1364 494
rect 1372 492 1454 494
rect 1482 492 1594 494
tri 730 488 734 492 se
rect 734 488 744 492
tri 728 486 730 488 se
rect 730 486 744 488
tri 724 482 728 486 se
rect 728 482 744 486
rect 1012 484 1054 492
rect 1312 484 1354 492
rect 1372 484 1384 492
rect 1392 484 1404 492
rect 1412 484 1424 492
rect 1432 484 1444 492
rect 1482 484 1494 492
rect 1502 484 1514 492
rect 1522 484 1534 492
rect 1542 484 1554 492
rect 1562 484 1574 492
rect 1582 490 1594 492
tri 1594 490 1598 494 nw
rect 1582 488 1592 490
tri 1592 488 1594 490 nw
rect 1582 484 1586 488
rect 1002 482 1054 484
rect 1302 482 1354 484
rect 1362 482 1444 484
rect 1472 482 1586 484
tri 1586 482 1592 488 nw
tri 722 480 724 482 se
rect 724 480 734 482
tri 718 476 722 480 se
rect 722 476 734 480
tri 716 474 718 476 se
rect 718 474 734 476
rect 1002 474 1044 482
rect 1302 474 1344 482
rect 1362 474 1374 482
rect 1382 474 1394 482
rect 1402 474 1414 482
rect 1422 474 1434 482
rect 1472 474 1484 482
rect 1492 474 1504 482
rect 1512 474 1524 482
rect 1532 474 1544 482
rect 1552 474 1564 482
rect 1572 476 1580 482
tri 1580 476 1586 482 nw
rect 1572 474 1578 476
tri 1578 474 1580 476 nw
tri 712 470 716 474 se
rect 716 472 734 474
rect 992 472 1044 474
rect 1292 472 1344 474
rect 1352 472 1434 474
rect 1462 472 1574 474
rect 716 470 724 472
tri 710 468 712 470 se
rect 712 468 724 470
tri 706 464 710 468 se
rect 710 464 724 468
rect 992 464 1034 472
rect 1292 464 1334 472
rect 1352 464 1364 472
rect 1372 464 1384 472
rect 1392 464 1404 472
rect 1412 464 1424 472
rect 1462 464 1474 472
rect 1482 464 1494 472
rect 1502 464 1514 472
rect 1522 464 1534 472
rect 1542 464 1554 472
rect 1562 470 1574 472
tri 1574 470 1578 474 nw
rect 1562 466 1570 470
tri 1570 466 1574 470 nw
rect 1562 464 1568 466
tri 1568 464 1570 466 nw
tri 704 462 706 464 se
rect 706 462 724 464
rect 982 462 1034 464
rect 1282 462 1334 464
rect 1342 462 1424 464
rect 1452 462 1562 464
tri 700 458 704 462 se
rect 704 458 714 462
tri 698 456 700 458 se
rect 700 456 714 458
tri 694 452 698 456 se
rect 698 452 714 456
rect 982 454 1024 462
rect 1282 454 1324 462
rect 1342 454 1354 462
rect 1362 454 1374 462
rect 1382 454 1394 462
rect 1402 454 1414 462
rect 1452 454 1464 462
rect 1472 454 1484 462
rect 1492 454 1504 462
rect 1512 454 1524 462
rect 1532 454 1544 462
rect 1552 458 1562 462
tri 1562 458 1568 464 nw
rect 1552 454 1556 458
rect 972 452 1024 454
rect 1272 452 1324 454
rect 1332 452 1414 454
rect 1442 452 1556 454
tri 1556 452 1562 458 nw
tri 692 450 694 452 se
rect 694 450 704 452
tri 690 448 692 450 se
rect 692 448 704 450
tri 686 444 690 448 se
rect 690 444 704 448
rect 972 444 1014 452
rect 1272 444 1314 452
rect 1332 444 1344 452
rect 1352 444 1364 452
rect 1372 444 1384 452
rect 1392 444 1404 452
rect 1442 444 1454 452
rect 1462 444 1474 452
rect 1482 444 1494 452
rect 1502 444 1514 452
rect 1522 444 1534 452
rect 1542 448 1552 452
tri 1552 448 1556 452 nw
rect 1542 444 1548 448
tri 1548 444 1552 448 nw
tri 684 442 686 444 se
rect 686 442 704 444
rect 962 442 1014 444
rect 1262 442 1314 444
rect 1322 442 1404 444
rect 1432 442 1546 444
tri 1546 442 1548 444 nw
tri 680 438 684 442 se
rect 684 438 694 442
tri 678 436 680 438 se
rect 680 436 694 438
tri 674 432 678 436 se
rect 678 432 694 436
rect 962 434 1004 442
rect 1262 434 1304 442
rect 1322 434 1334 442
rect 1342 434 1354 442
rect 1362 434 1374 442
rect 1382 434 1394 442
rect 1432 434 1444 442
rect 1452 434 1464 442
rect 1472 434 1484 442
rect 1492 434 1504 442
rect 1512 434 1524 442
rect 1532 436 1540 442
tri 1540 436 1546 442 nw
rect 1532 434 1534 436
rect 952 432 1004 434
rect 1252 432 1304 434
rect 1312 432 1394 434
rect 1422 432 1534 434
tri 672 430 674 432 se
rect 674 430 684 432
tri 668 426 672 430 se
rect 672 426 684 430
tri 666 424 668 426 se
rect 668 424 684 426
rect 952 424 994 432
rect 1252 424 1294 432
rect 1312 424 1324 432
rect 1332 424 1344 432
rect 1352 424 1364 432
rect 1372 424 1384 432
rect 1422 424 1434 432
rect 1442 424 1454 432
rect 1462 424 1474 432
rect 1482 424 1494 432
rect 1502 424 1514 432
rect 1522 430 1534 432
tri 1534 430 1540 436 nw
rect 1522 428 1532 430
tri 1532 428 1534 430 nw
rect 1522 424 1528 428
tri 1528 424 1532 428 nw
tri 662 420 666 424 se
rect 666 422 684 424
rect 942 422 994 424
rect 1242 422 1294 424
rect 1302 422 1384 424
rect 1412 422 1524 424
rect 666 420 674 422
tri 660 418 662 420 se
rect 662 418 674 420
rect 660 412 674 418
rect 942 414 984 422
rect 1242 414 1284 422
rect 1302 414 1314 422
rect 1322 414 1334 422
rect 1342 414 1354 422
rect 1362 414 1374 422
rect 1412 414 1424 422
rect 1432 414 1444 422
rect 1452 414 1464 422
rect 1472 414 1484 422
rect 1492 414 1504 422
rect 1512 420 1524 422
tri 1524 420 1528 424 nw
rect 1512 418 1522 420
tri 1522 418 1524 420 nw
rect 1512 414 1516 418
rect 932 412 984 414
rect 1232 412 1284 414
rect 1292 412 1374 414
rect 1402 412 1516 414
tri 1516 412 1522 418 nw
rect 660 4 664 412
rect 932 402 974 412
rect 1232 404 1274 412
rect 1292 404 1304 412
rect 1312 404 1324 412
rect 1332 404 1344 412
rect 1352 404 1364 412
rect 1402 404 1414 412
rect 1422 404 1434 412
rect 1442 404 1454 412
rect 1462 404 1474 412
rect 1482 404 1494 412
rect 1502 410 1514 412
tri 1514 410 1516 412 nw
rect 1502 406 1510 410
tri 1510 406 1514 410 nw
rect 1502 404 1506 406
rect 1222 402 1274 404
rect 1282 402 1364 404
rect 1392 402 1506 404
tri 1506 402 1510 406 nw
rect 932 392 964 402
rect 1222 394 1264 402
rect 1282 394 1294 402
rect 1302 394 1314 402
rect 1322 394 1334 402
rect 1342 394 1354 402
rect 1392 394 1404 402
rect 1412 394 1424 402
rect 1432 394 1444 402
rect 1452 394 1464 402
rect 1472 394 1484 402
rect 1492 400 1504 402
tri 1504 400 1506 402 nw
rect 1492 394 1498 400
tri 1498 394 1504 400 nw
rect 1212 392 1264 394
rect 1272 392 1354 394
rect 1382 392 1492 394
rect 932 382 954 392
rect 1212 384 1254 392
rect 1272 384 1284 392
rect 1292 384 1304 392
rect 1312 384 1324 392
rect 1332 384 1344 392
rect 1382 384 1394 392
rect 1402 384 1414 392
rect 1422 384 1434 392
rect 1442 384 1454 392
rect 1462 384 1474 392
rect 1482 388 1492 392
tri 1492 388 1498 394 nw
rect 1482 386 1490 388
tri 1490 386 1492 388 nw
rect 1482 384 1488 386
tri 1488 384 1490 386 nw
rect 1202 382 1254 384
rect 1262 382 1344 384
rect 1372 382 1482 384
rect 1202 374 1244 382
rect 1262 374 1274 382
rect 1282 374 1294 382
rect 1302 374 1314 382
rect 1322 374 1334 382
rect 1372 374 1384 382
rect 1392 374 1404 382
rect 1412 374 1424 382
rect 1432 374 1444 382
rect 1452 374 1464 382
rect 1472 378 1482 382
tri 1482 378 1488 384 nw
rect 1472 374 1476 378
rect 1192 372 1244 374
rect 1252 372 1334 374
rect 1362 372 1476 374
tri 1476 372 1482 378 nw
rect 1192 364 1234 372
rect 1252 364 1264 372
rect 1272 364 1284 372
rect 1292 364 1304 372
rect 1312 364 1324 372
rect 1362 364 1374 372
rect 1382 364 1394 372
rect 1402 364 1414 372
rect 1422 364 1434 372
rect 1442 364 1454 372
rect 1462 370 1474 372
tri 1474 370 1476 372 nw
rect 1462 366 1470 370
tri 1470 366 1474 370 nw
rect 1462 364 1468 366
tri 1468 364 1470 366 nw
rect 1182 362 1234 364
rect 1242 362 1324 364
rect 1352 362 1466 364
tri 1466 362 1468 364 nw
rect 1182 354 1224 362
rect 1242 354 1254 362
rect 1262 354 1274 362
rect 1282 354 1294 362
rect 1302 354 1314 362
rect 1352 354 1364 362
rect 1372 354 1384 362
rect 1392 354 1404 362
rect 1412 354 1424 362
rect 1432 354 1444 362
rect 1452 360 1464 362
tri 1464 360 1466 362 nw
rect 1452 354 1458 360
tri 1458 354 1464 360 nw
rect 1172 352 1224 354
rect 1232 352 1314 354
rect 1342 352 1452 354
rect 1172 344 1214 352
rect 1232 344 1244 352
rect 1252 344 1264 352
rect 1272 344 1284 352
rect 1292 344 1304 352
rect 1342 344 1354 352
rect 1362 344 1374 352
rect 1382 344 1394 352
rect 1402 344 1414 352
rect 1422 344 1434 352
rect 1442 348 1452 352
tri 1452 348 1458 354 nw
rect 1442 346 1450 348
tri 1450 346 1452 348 nw
rect 1442 344 1446 346
rect 1162 342 1214 344
rect 1222 342 1304 344
rect 1332 342 1446 344
tri 1446 342 1450 346 nw
rect 1162 334 1204 342
rect 1222 334 1234 342
rect 1242 334 1254 342
rect 1262 334 1274 342
rect 1282 334 1294 342
rect 1332 334 1344 342
rect 1352 334 1364 342
rect 1372 334 1384 342
rect 1392 334 1404 342
rect 1412 334 1424 342
rect 1432 338 1442 342
tri 1442 338 1446 342 nw
rect 1432 336 1440 338
tri 1440 336 1442 338 nw
rect 1432 334 1434 336
rect 1152 332 1204 334
rect 1212 332 1294 334
rect 1322 332 1434 334
rect 1152 324 1194 332
rect 1212 324 1224 332
rect 1232 324 1244 332
rect 1252 324 1264 332
rect 1272 324 1284 332
rect 1322 324 1334 332
rect 1342 324 1354 332
rect 1362 324 1374 332
rect 1382 324 1394 332
rect 1402 324 1414 332
rect 1422 330 1434 332
tri 1434 330 1440 336 nw
rect 1422 324 1428 330
tri 1428 324 1434 330 nw
rect 1142 322 1194 324
rect 1202 322 1284 324
rect 1312 322 1426 324
tri 1426 322 1428 324 nw
rect 1142 314 1184 322
rect 1202 314 1214 322
rect 1222 314 1234 322
rect 1242 314 1254 322
rect 1262 314 1274 322
rect 1312 314 1324 322
rect 1332 314 1344 322
rect 1352 314 1364 322
rect 1372 314 1384 322
rect 1392 314 1404 322
rect 1412 320 1424 322
tri 1424 320 1426 322 nw
rect 1412 314 1418 320
tri 1418 314 1424 320 nw
rect 1132 312 1184 314
rect 1192 312 1274 314
rect 1302 312 1412 314
rect 1132 304 1174 312
rect 1192 304 1204 312
rect 1212 304 1224 312
rect 1232 304 1244 312
rect 1252 304 1264 312
rect 1302 304 1314 312
rect 1322 304 1334 312
rect 1342 304 1354 312
rect 1362 304 1374 312
rect 1382 304 1394 312
rect 1402 308 1412 312
tri 1412 308 1418 314 nw
rect 1402 306 1410 308
tri 1410 306 1412 308 nw
rect 1402 304 1406 306
rect 1122 302 1174 304
rect 1182 302 1264 304
rect 1292 302 1406 304
tri 1406 302 1410 306 nw
rect 1122 294 1164 302
rect 1182 294 1194 302
rect 1202 294 1214 302
rect 1222 294 1234 302
rect 1242 294 1254 302
rect 1292 294 1304 302
rect 1312 294 1324 302
rect 1332 294 1344 302
rect 1352 294 1364 302
rect 1372 294 1384 302
rect 1392 298 1402 302
tri 1402 298 1406 302 nw
rect 1392 296 1400 298
tri 1400 296 1402 298 nw
rect 1392 294 1394 296
rect 1112 292 1164 294
rect 1172 292 1254 294
rect 1282 292 1394 294
rect 1112 282 1154 292
rect 1172 284 1184 292
rect 1192 284 1204 292
rect 1212 284 1224 292
rect 1232 284 1244 292
rect 1282 284 1294 292
rect 1302 284 1314 292
rect 1322 284 1334 292
rect 1342 284 1354 292
rect 1362 284 1374 292
rect 1382 290 1394 292
tri 1394 290 1400 296 nw
rect 1382 284 1388 290
tri 1388 284 1394 290 nw
rect 1162 282 1244 284
rect 1272 282 1386 284
tri 1386 282 1388 284 nw
rect 1112 274 1144 282
rect 1162 274 1174 282
rect 1182 274 1194 282
rect 1202 274 1214 282
rect 1222 274 1234 282
rect 1272 274 1284 282
rect 1292 274 1304 282
rect 1312 274 1324 282
rect 1332 274 1344 282
rect 1352 274 1364 282
rect 1372 280 1384 282
tri 1384 280 1386 282 nw
rect 1372 274 1378 280
tri 1378 274 1384 280 nw
rect 1092 272 1144 274
rect 1152 272 1234 274
rect 1262 272 1372 274
rect 1092 242 1134 272
rect 1152 244 1164 272
rect 1172 244 1184 272
rect 1192 264 1204 272
rect 1212 264 1224 272
rect 1192 262 1224 264
rect 1202 244 1214 262
rect 1232 244 1244 264
rect 1262 244 1274 272
rect 1282 264 1294 272
rect 1302 264 1314 272
rect 1282 262 1314 264
rect 1292 244 1304 262
rect 1322 244 1334 272
rect 1342 264 1354 272
rect 1362 268 1372 272
tri 1372 268 1378 274 nw
rect 1362 266 1370 268
tri 1370 266 1372 268 nw
rect 1362 264 1366 266
rect 1342 262 1366 264
tri 1366 262 1370 266 nw
rect 1352 258 1362 262
tri 1362 258 1366 262 nw
rect 1352 256 1360 258
tri 1360 256 1362 258 nw
rect 1352 254 1354 256
rect 1342 250 1354 254
tri 1354 250 1360 256 nw
rect 1342 244 1348 250
tri 1348 244 1354 250 nw
rect 1152 242 1184 244
rect 1192 242 1214 244
rect 1222 242 1244 244
rect 1252 242 1274 244
rect 1282 242 1304 244
rect 1312 242 1346 244
tri 1346 242 1348 244 nw
rect 1162 234 1174 242
rect 1192 234 1204 242
rect 1222 234 1234 242
rect 1252 234 1264 242
rect 1282 234 1294 242
rect 1312 234 1324 242
rect 1332 240 1344 242
tri 1344 240 1346 242 nw
rect 1332 238 1342 240
tri 1342 238 1344 240 nw
rect 1332 236 1340 238
tri 1340 236 1342 238 nw
rect 1332 234 1338 236
tri 1338 234 1340 236 nw
rect 1162 232 1184 234
rect 1192 232 1214 234
rect 1222 232 1244 234
rect 1252 232 1274 234
rect 1282 232 1304 234
rect 1312 232 1334 234
rect 1172 224 1184 232
rect 1202 224 1214 232
rect 1232 224 1244 232
rect 1262 224 1274 232
rect 1292 224 1304 232
rect 1322 230 1334 232
tri 1334 230 1338 234 nw
rect 1322 228 1332 230
tri 1332 228 1334 230 nw
rect 1322 224 1326 228
rect 1162 222 1184 224
rect 1192 222 1214 224
rect 1222 222 1244 224
rect 1252 222 1274 224
rect 1282 222 1304 224
rect 1312 222 1326 224
tri 1326 222 1332 228 nw
rect 1162 214 1174 222
rect 1192 214 1204 222
rect 1222 214 1234 222
rect 1252 214 1264 222
rect 1282 214 1294 222
rect 1312 216 1320 222
tri 1320 216 1326 222 nw
rect 1312 214 1318 216
tri 1318 214 1320 216 nw
rect 1162 212 1184 214
rect 1192 212 1214 214
rect 1222 212 1244 214
rect 1252 212 1274 214
rect 1282 212 1304 214
rect 1172 204 1184 212
rect 1202 204 1214 212
rect 1232 204 1244 212
rect 1262 204 1274 212
rect 1292 204 1304 212
rect 1162 202 1184 204
rect 1192 202 1214 204
rect 1222 202 1244 204
rect 1252 202 1274 204
rect 1282 202 1304 204
rect 1162 194 1174 202
rect 1192 194 1204 202
rect 1222 194 1234 202
rect 1252 194 1264 202
rect 1282 194 1294 202
rect 1162 192 1184 194
rect 1192 192 1214 194
rect 1222 192 1244 194
rect 1252 192 1274 194
rect 1282 192 1304 194
rect 1172 184 1184 192
rect 1202 184 1214 192
rect 1232 184 1244 192
rect 1262 184 1274 192
rect 1292 184 1304 192
rect 1162 182 1184 184
rect 1192 182 1214 184
rect 1222 182 1244 184
rect 1252 182 1274 184
rect 1282 182 1304 184
rect 1162 174 1174 182
rect 1192 174 1204 182
rect 1222 174 1234 182
rect 1252 174 1264 182
rect 1282 174 1294 182
rect 1162 172 1184 174
rect 1192 172 1214 174
rect 1222 172 1244 174
rect 1252 172 1274 174
rect 1282 172 1304 174
rect 1172 164 1184 172
rect 1202 164 1214 172
rect 1232 164 1244 172
rect 1262 164 1274 172
rect 1292 164 1304 172
rect 1162 162 1184 164
rect 1192 162 1214 164
rect 1222 162 1244 164
rect 1252 162 1274 164
rect 1282 162 1304 164
rect 1162 154 1174 162
rect 1192 154 1204 162
rect 1222 154 1234 162
rect 1252 154 1264 162
rect 1282 154 1294 162
rect 1162 152 1184 154
rect 1192 152 1214 154
rect 1222 152 1244 154
rect 1252 152 1274 154
rect 1282 152 1304 154
rect 1172 144 1184 152
rect 1202 144 1214 152
rect 1232 144 1244 152
rect 1262 144 1274 152
rect 1292 144 1304 152
rect 1162 142 1184 144
rect 1192 142 1214 144
rect 1222 142 1244 144
rect 1252 142 1274 144
rect 1282 142 1304 144
rect 1162 134 1174 142
rect 1192 134 1204 142
rect 1222 134 1234 142
rect 1252 134 1264 142
rect 1282 134 1294 142
rect 1162 132 1184 134
rect 1192 132 1214 134
rect 1222 132 1244 134
rect 1252 132 1274 134
rect 1282 132 1304 134
rect 1172 124 1184 132
rect 1202 124 1214 132
rect 1232 124 1244 132
rect 1262 124 1274 132
rect 1292 124 1304 132
rect 1162 122 1184 124
rect 1192 122 1214 124
rect 1222 122 1244 124
rect 1252 122 1274 124
rect 1282 122 1304 124
rect 1162 114 1174 122
rect 1192 114 1204 122
rect 1222 114 1234 122
rect 1252 114 1264 122
rect 1282 114 1294 122
rect 1162 112 1184 114
rect 1192 112 1214 114
rect 1222 112 1244 114
rect 1252 112 1274 114
rect 1282 112 1304 114
rect 1172 104 1184 112
rect 1202 104 1214 112
rect 1232 104 1244 112
rect 1262 104 1274 112
rect 1292 104 1304 112
rect 1162 102 1184 104
rect 1192 102 1214 104
rect 1222 102 1244 104
rect 1252 102 1274 104
rect 1282 102 1304 104
rect 1162 94 1174 102
rect 1192 94 1204 102
rect 1222 94 1234 102
rect 1252 94 1264 102
rect 1282 94 1294 102
rect 1162 92 1184 94
rect 1192 92 1214 94
rect 1222 92 1244 94
rect 1252 92 1274 94
rect 1282 92 1304 94
rect 1172 84 1184 92
rect 1202 84 1214 92
rect 1232 84 1244 92
rect 1262 84 1274 92
rect 1292 84 1304 92
rect 1162 82 1184 84
rect 1192 82 1214 84
rect 1222 82 1244 84
rect 1252 82 1274 84
rect 1282 82 1304 84
rect 1162 74 1174 82
rect 1192 74 1204 82
rect 1222 74 1234 82
rect 1252 74 1264 82
rect 1282 74 1294 82
rect 1162 72 1184 74
rect 1192 72 1214 74
rect 1222 72 1244 74
rect 1252 72 1274 74
rect 1282 72 1304 74
rect 1172 64 1184 72
rect 1202 64 1214 72
rect 1232 64 1244 72
rect 1262 64 1274 72
rect 1292 64 1304 72
rect 1162 62 1184 64
rect 1192 62 1214 64
rect 1222 62 1244 64
rect 1252 62 1274 64
rect 1282 62 1304 64
rect 1162 54 1174 62
rect 1192 54 1204 62
rect 1222 54 1234 62
rect 1252 54 1264 62
rect 1282 54 1294 62
rect 1162 52 1184 54
rect 1192 52 1214 54
rect 1222 52 1244 54
rect 1252 52 1274 54
rect 1282 52 1304 54
rect 1172 44 1184 52
rect 1202 44 1214 52
rect 1232 44 1244 52
rect 1262 44 1274 52
rect 1292 44 1304 52
rect 1162 42 1184 44
rect 1192 42 1214 44
rect 1222 42 1244 44
rect 1252 42 1274 44
rect 1282 42 1304 44
rect 1162 34 1174 42
rect 1192 34 1204 42
rect 1222 34 1234 42
rect 1252 34 1264 42
rect 1282 34 1294 42
rect 1162 32 1184 34
rect 1192 32 1214 34
rect 1222 32 1244 34
rect 1252 32 1274 34
rect 1282 32 1304 34
rect 1172 24 1184 32
rect 1202 24 1214 32
rect 1232 24 1244 32
rect 1262 24 1274 32
rect 1292 24 1304 32
rect 1162 22 1184 24
rect 1192 22 1214 24
rect 1222 22 1244 24
rect 1252 22 1274 24
rect 1282 22 1304 24
rect 1162 14 1174 22
rect 1192 14 1204 22
rect 1222 14 1234 22
rect 1252 14 1264 22
rect 1282 14 1294 22
rect 1162 12 1184 14
rect 1192 12 1214 14
rect 1222 12 1244 14
rect 1252 12 1274 14
rect 1282 12 1304 14
rect 1172 4 1184 12
rect 1202 4 1214 12
rect 1232 4 1244 12
rect 1262 4 1274 12
rect 1292 4 1304 12
rect 1312 4 1314 214
tri 1314 210 1318 214 nw
rect 660 0 1314 4
<< nsubstratendiff >>
tri 1820 652 1822 654 se
rect 1822 652 2000 654
tri 1818 650 1820 652 se
rect 1820 650 2000 652
tri 1814 646 1818 650 se
rect 1818 646 2000 650
tri 1808 640 1814 646 se
rect 1814 642 2000 646
rect 1814 640 1820 642
tri 1802 634 1808 640 se
rect 1808 634 1820 640
tri 1796 628 1802 634 se
rect 1802 632 1820 634
rect 1828 634 1840 642
rect 1858 634 1870 642
rect 1888 634 1900 642
rect 1918 634 1930 642
rect 1948 634 1960 642
rect 1978 634 1990 642
rect 1998 634 2000 642
rect 1828 632 1850 634
rect 1858 632 1880 634
rect 1888 632 1910 634
rect 1918 632 1940 634
rect 1948 632 1970 634
rect 1978 632 2000 634
rect 1802 628 1810 632
tri 1792 624 1796 628 se
rect 1796 624 1810 628
rect 1838 624 1850 632
rect 1868 624 1880 632
rect 1898 624 1910 632
rect 1928 624 1940 632
rect 1958 624 1970 632
rect 1988 624 2000 632
tri 1790 622 1792 624 se
rect 1792 622 1810 624
rect 1828 622 1850 624
rect 1858 622 1880 624
rect 1888 622 1910 624
rect 1918 622 1940 624
rect 1948 622 1970 624
rect 1978 622 2000 624
tri 1784 616 1790 622 se
rect 1790 616 1800 622
tri 1778 610 1784 616 se
rect 1784 612 1800 616
rect 1828 614 1840 622
rect 1858 614 1870 622
rect 1888 614 1900 622
rect 1918 614 1930 622
rect 1948 614 1960 622
rect 1978 614 1990 622
rect 1998 614 2000 622
rect 1784 610 1790 612
tri 1772 604 1778 610 se
rect 1778 604 1790 610
rect 1808 604 1820 614
rect 1828 612 1850 614
rect 1858 612 1880 614
rect 1888 612 1910 614
rect 1918 612 1940 614
rect 1948 612 1970 614
rect 1978 612 2000 614
rect 1838 604 1850 612
rect 1868 604 1880 612
rect 1898 604 1910 612
rect 1928 604 1940 612
rect 1958 604 1970 612
rect 1988 604 2000 612
tri 1766 598 1772 604 se
rect 1772 602 1790 604
rect 1798 602 1820 604
rect 1828 602 1850 604
rect 1858 602 1880 604
rect 1888 602 1910 604
rect 1918 602 1940 604
rect 1948 602 1970 604
rect 1978 602 2000 604
rect 1772 598 1780 602
tri 1760 592 1766 598 se
rect 1766 592 1780 598
rect 1798 594 1810 602
rect 1788 592 1810 594
rect 1828 594 1840 602
rect 1858 594 1870 602
rect 1888 594 1900 602
rect 1918 594 1930 602
rect 1948 594 1960 602
rect 1978 594 1990 602
rect 1998 594 2000 602
rect 1828 592 1850 594
rect 1858 592 1880 594
rect 1888 592 1910 594
rect 1918 592 1940 594
rect 1948 592 1970 594
rect 1978 592 2000 594
tri 1756 588 1760 592 se
rect 1760 588 1770 592
tri 1750 582 1756 588 se
rect 1756 582 1770 588
rect 1788 584 1800 592
rect 1838 584 1850 592
rect 1778 582 1800 584
tri 1744 576 1750 582 se
rect 1750 576 1760 582
tri 1738 570 1744 576 se
rect 1744 572 1760 576
rect 1778 574 1790 582
rect 1808 574 1820 584
rect 1768 572 1790 574
rect 1798 572 1820 574
rect 1828 582 1850 584
rect 1868 582 1880 592
rect 1898 584 1910 592
rect 1928 584 1940 592
rect 1958 584 1970 592
rect 1988 584 2000 592
rect 1888 582 1910 584
rect 1918 582 1940 584
rect 1948 582 1970 584
rect 1978 582 2000 584
rect 1828 572 1840 582
rect 1888 574 1900 582
rect 1918 574 1930 582
rect 1948 574 1960 582
rect 1978 574 1990 582
rect 1998 574 2000 582
rect 1744 570 1750 572
tri 1732 564 1738 570 se
rect 1738 564 1750 570
rect 1768 564 1780 572
rect 1798 564 1810 572
rect 1868 564 1880 574
rect 1888 572 1910 574
rect 1918 572 1940 574
rect 1948 572 1970 574
rect 1978 572 2000 574
rect 1898 564 1910 572
rect 1928 564 1940 572
rect 1958 564 1970 572
rect 1988 564 2000 572
tri 1726 558 1732 564 se
rect 1732 562 1750 564
rect 1758 562 1780 564
rect 1788 562 1810 564
rect 1858 562 1880 564
rect 1888 562 1910 564
rect 1918 562 1940 564
rect 1948 562 1970 564
rect 1978 562 2000 564
rect 1732 558 1740 562
tri 1720 552 1726 558 se
rect 1726 552 1740 558
rect 1758 554 1770 562
rect 1788 554 1800 562
rect 1858 554 1870 562
rect 1888 554 1900 562
rect 1918 554 1930 562
rect 1948 554 1960 562
rect 1978 554 1990 562
rect 1998 554 2000 562
rect 1748 552 1770 554
rect 1778 552 1800 554
tri 1714 546 1720 552 se
rect 1720 546 1730 552
tri 1708 540 1714 546 se
rect 1714 542 1730 546
rect 1748 544 1760 552
rect 1778 544 1790 552
rect 1838 544 1850 554
rect 1858 552 1880 554
rect 1888 552 1910 554
rect 1918 552 1940 554
rect 1948 552 1970 554
rect 1978 552 2000 554
rect 1868 544 1880 552
rect 1898 544 1910 552
rect 1928 544 1940 552
rect 1958 544 1970 552
rect 1988 544 2000 552
rect 1738 542 1760 544
rect 1768 542 1790 544
rect 1828 542 1850 544
rect 1858 542 1880 544
rect 1888 542 1910 544
rect 1918 542 1940 544
rect 1948 542 1970 544
rect 1978 542 2000 544
rect 1714 540 1720 542
tri 1702 534 1708 540 se
rect 1708 534 1720 540
rect 1738 534 1750 542
rect 1768 534 1780 542
rect 1828 534 1840 542
rect 1858 534 1870 542
rect 1888 534 1900 542
rect 1918 534 1930 542
rect 1948 534 1960 542
rect 1978 534 1990 542
rect 1998 534 2000 542
tri 1696 528 1702 534 se
rect 1702 532 1720 534
rect 1728 532 1750 534
rect 1758 532 1780 534
rect 1702 528 1710 532
tri 1690 522 1696 528 se
rect 1696 522 1710 528
rect 1728 524 1740 532
rect 1758 524 1770 532
rect 1808 531 1820 534
rect 1828 532 1850 534
rect 1858 532 1880 534
rect 1888 532 1910 534
rect 1918 532 1940 534
rect 1948 532 1970 534
rect 1978 532 2000 534
rect 1838 524 1850 532
rect 1868 524 1880 532
rect 1898 524 1910 532
rect 1928 524 1940 532
rect 1958 524 1970 532
rect 1988 524 2000 532
rect 1718 522 1740 524
rect 1748 522 1770 524
tri 1684 516 1690 522 se
rect 1690 516 1700 522
tri 1680 512 1684 516 se
rect 1684 512 1700 516
rect 1718 514 1730 522
rect 1748 514 1760 522
rect 1808 514 1820 523
rect 1708 512 1730 514
rect 1738 512 1760 514
rect 1798 512 1820 514
rect 1828 522 1850 524
rect 1858 522 1880 524
rect 1888 522 1910 524
rect 1918 522 1940 524
rect 1948 522 1970 524
rect 1978 522 2000 524
rect 1828 514 1840 522
rect 1858 514 1870 522
rect 1888 514 1900 522
rect 1918 514 1930 522
rect 1948 514 1960 522
rect 1978 514 1990 522
rect 1998 514 2000 522
rect 1828 512 1850 514
rect 1858 512 1880 514
rect 1888 512 1910 514
rect 1918 512 1940 514
rect 1948 512 1970 514
rect 1978 512 2000 514
tri 1674 506 1680 512 se
rect 1680 506 1690 512
tri 1668 500 1674 506 se
rect 1674 502 1690 506
rect 1708 502 1720 512
rect 1738 502 1750 512
rect 1798 502 1810 512
rect 1838 502 1850 512
rect 1868 502 1880 512
rect 1898 502 1910 512
rect 1928 502 1940 512
rect 1958 502 1970 512
rect 1988 502 2000 512
rect 1674 500 1680 502
tri 1662 494 1668 500 se
rect 1668 494 1680 500
tri 1656 488 1662 494 se
rect 1662 492 1690 494
rect 1662 488 1670 492
tri 1650 482 1656 488 se
rect 1656 484 1670 488
rect 1678 484 1690 492
rect 1698 484 1710 494
rect 1718 484 1730 494
rect 1738 484 1750 494
rect 1788 484 1800 494
rect 1808 484 1820 494
rect 1828 484 1840 494
rect 1848 484 1860 494
rect 1868 484 1890 494
rect 1656 482 1750 484
rect 1778 482 1890 484
tri 1644 476 1650 482 se
rect 1650 476 1660 482
tri 1638 470 1644 476 se
rect 1644 474 1660 476
rect 1668 474 1680 482
rect 1688 474 1700 482
rect 1708 474 1720 482
rect 1728 474 1740 482
rect 1778 474 1790 482
rect 1798 474 1810 482
rect 1818 474 1830 482
rect 1838 474 1850 482
rect 1858 474 1880 482
rect 1644 472 1740 474
rect 1768 472 1880 474
rect 1644 470 1650 472
tri 1632 464 1638 470 se
rect 1638 464 1650 470
rect 1658 464 1670 472
rect 1678 464 1690 472
rect 1698 464 1710 472
rect 1718 464 1730 472
rect 1768 464 1780 472
rect 1788 464 1800 472
rect 1808 464 1820 472
rect 1828 464 1840 472
rect 1848 464 1870 472
tri 1626 458 1632 464 se
rect 1632 462 1730 464
rect 1758 462 1870 464
rect 1632 458 1640 462
tri 1620 452 1626 458 se
rect 1626 454 1640 458
rect 1648 454 1660 462
rect 1668 454 1680 462
rect 1688 454 1700 462
rect 1708 454 1720 462
rect 1758 454 1770 462
rect 1778 454 1790 462
rect 1798 454 1810 462
rect 1818 454 1830 462
rect 1838 454 1860 462
rect 1626 452 1720 454
rect 1748 452 1860 454
tri 1616 448 1620 452 se
rect 1620 448 1630 452
tri 1610 442 1616 448 se
rect 1616 444 1630 448
rect 1638 444 1650 452
rect 1658 444 1670 452
rect 1678 444 1690 452
rect 1698 444 1710 452
rect 1748 444 1760 452
rect 1768 444 1780 452
rect 1788 444 1800 452
rect 1808 444 1820 452
rect 1828 444 1850 452
rect 1616 442 1710 444
rect 1738 442 1850 444
tri 1604 436 1610 442 se
rect 1610 436 1620 442
tri 1598 430 1604 436 se
rect 1604 434 1620 436
rect 1628 434 1640 442
rect 1648 434 1660 442
rect 1668 434 1680 442
rect 1688 434 1700 442
rect 1738 434 1750 442
rect 1758 434 1770 442
rect 1778 434 1790 442
rect 1798 434 1810 442
rect 1818 434 1840 442
rect 1604 432 1700 434
rect 1728 432 1840 434
rect 1604 430 1610 432
tri 1592 424 1598 430 se
rect 1598 424 1610 430
rect 1618 424 1630 432
rect 1638 424 1650 432
rect 1658 424 1670 432
rect 1678 424 1690 432
rect 1728 424 1740 432
rect 1748 424 1760 432
rect 1768 424 1780 432
rect 1788 424 1800 432
rect 1808 424 1830 432
tri 1588 420 1592 424 se
rect 1592 422 1690 424
rect 1718 422 1830 424
rect 1592 420 1600 422
tri 1586 418 1588 420 se
rect 1588 418 1600 420
tri 1580 412 1586 418 se
rect 1586 414 1600 418
rect 1608 414 1620 422
rect 1628 414 1640 422
rect 1648 414 1660 422
rect 1668 414 1680 422
rect 1718 414 1730 422
rect 1738 414 1750 422
rect 1758 414 1770 422
rect 1778 414 1790 422
rect 1798 414 1830 422
rect 1586 412 1680 414
rect 1708 412 1840 414
tri 1574 406 1580 412 se
rect 1580 406 1590 412
tri 1568 400 1574 406 se
rect 1574 404 1590 406
rect 1598 404 1610 412
rect 1618 404 1630 412
rect 1638 404 1650 412
rect 1658 404 1670 412
rect 1708 404 1720 412
rect 1728 404 1740 412
rect 1748 404 1760 412
rect 1768 404 1780 412
rect 1788 404 1840 412
rect 1574 402 1670 404
rect 1698 402 1840 404
rect 1574 400 1580 402
tri 1562 394 1568 400 se
rect 1568 394 1580 400
rect 1588 394 1600 402
rect 1608 394 1620 402
rect 1628 394 1640 402
rect 1648 394 1660 402
rect 1698 394 1710 402
rect 1718 394 1730 402
rect 1738 394 1750 402
rect 1758 394 1770 402
rect 1778 394 1830 402
tri 1556 388 1562 394 se
rect 1562 392 1660 394
rect 1688 392 1830 394
rect 1562 388 1570 392
tri 1552 384 1556 388 se
rect 1556 384 1570 388
rect 1578 384 1590 392
rect 1598 384 1610 392
rect 1618 384 1630 392
rect 1638 384 1650 392
rect 1688 384 1700 392
rect 1708 384 1720 392
rect 1728 384 1740 392
rect 1748 384 1760 392
rect 1768 384 1820 392
tri 1546 378 1552 384 se
rect 1552 382 1650 384
rect 1678 382 1820 384
rect 1552 378 1560 382
tri 1540 372 1546 378 se
rect 1546 374 1560 378
rect 1568 374 1580 382
rect 1588 374 1600 382
rect 1608 374 1620 382
rect 1628 374 1640 382
rect 1678 374 1690 382
rect 1698 374 1710 382
rect 1718 374 1730 382
rect 1738 374 1750 382
rect 1758 374 1810 382
rect 1546 372 1640 374
rect 1668 372 1810 374
tri 1534 366 1540 372 se
rect 1540 366 1550 372
tri 1532 364 1534 366 se
rect 1534 364 1550 366
rect 1558 364 1570 372
rect 1578 364 1590 372
rect 1598 364 1610 372
rect 1618 364 1630 372
rect 1668 364 1680 372
rect 1688 364 1700 372
rect 1708 364 1720 372
rect 1728 364 1740 372
rect 1748 364 1800 372
tri 1528 360 1532 364 se
rect 1532 362 1630 364
rect 1658 362 1800 364
rect 1532 360 1540 362
tri 1522 354 1528 360 se
rect 1528 354 1540 360
rect 1548 354 1560 362
rect 1568 354 1580 362
rect 1588 354 1600 362
rect 1608 354 1620 362
rect 1658 354 1670 362
rect 1678 354 1690 362
rect 1698 354 1710 362
rect 1718 354 1730 362
rect 1738 354 1790 362
tri 1516 348 1522 354 se
rect 1522 352 1620 354
rect 1648 352 1790 354
rect 1522 348 1530 352
tri 1510 342 1516 348 se
rect 1516 344 1530 348
rect 1538 344 1550 352
rect 1558 344 1570 352
rect 1578 344 1590 352
rect 1598 344 1610 352
rect 1648 344 1660 352
rect 1668 344 1680 352
rect 1688 344 1700 352
rect 1708 344 1720 352
rect 1728 344 1780 352
rect 1516 342 1610 344
rect 1638 342 1780 344
tri 1504 336 1510 342 se
rect 1510 336 1520 342
tri 1498 330 1504 336 se
rect 1504 334 1520 336
rect 1528 334 1540 342
rect 1548 334 1560 342
rect 1568 334 1580 342
rect 1588 334 1600 342
rect 1638 334 1650 342
rect 1658 334 1670 342
rect 1678 334 1690 342
rect 1698 334 1710 342
rect 1718 334 1770 342
rect 1504 332 1600 334
rect 1628 332 1770 334
rect 1504 330 1510 332
tri 1492 324 1498 330 se
rect 1498 324 1510 330
rect 1518 324 1530 332
rect 1538 324 1550 332
rect 1558 324 1570 332
rect 1578 324 1590 332
rect 1628 324 1640 332
rect 1648 324 1660 332
rect 1668 324 1680 332
rect 1688 324 1700 332
rect 1708 324 1760 332
tri 1488 320 1492 324 se
rect 1492 322 1590 324
rect 1618 322 1760 324
rect 1492 320 1500 322
tri 1482 314 1488 320 se
rect 1488 314 1500 320
rect 1508 314 1520 322
rect 1528 314 1540 322
rect 1548 314 1560 322
rect 1568 314 1580 322
rect 1618 314 1630 322
rect 1638 314 1650 322
rect 1658 314 1670 322
rect 1678 314 1690 322
rect 1698 314 1750 322
tri 1476 308 1482 314 se
rect 1482 312 1580 314
rect 1608 312 1750 314
rect 1482 308 1490 312
tri 1470 302 1476 308 se
rect 1476 304 1490 308
rect 1498 304 1510 312
rect 1518 304 1530 312
rect 1538 304 1550 312
rect 1558 304 1570 312
rect 1608 304 1620 312
rect 1628 304 1640 312
rect 1648 304 1660 312
rect 1668 304 1680 312
rect 1688 304 1740 312
rect 1476 302 1570 304
rect 1598 302 1740 304
tri 1464 296 1470 302 se
rect 1470 296 1480 302
tri 1458 290 1464 296 se
rect 1464 294 1480 296
rect 1488 294 1500 302
rect 1508 294 1520 302
rect 1528 294 1540 302
rect 1548 294 1560 302
rect 1598 294 1610 302
rect 1618 294 1630 302
rect 1638 294 1650 302
rect 1658 294 1670 302
rect 1678 294 1730 302
rect 1464 292 1560 294
rect 1588 292 1730 294
rect 1464 290 1470 292
tri 1452 284 1458 290 se
rect 1458 284 1470 290
rect 1478 284 1490 292
rect 1498 284 1510 292
rect 1518 284 1530 292
rect 1538 284 1550 292
rect 1588 284 1600 292
rect 1608 284 1620 292
rect 1628 284 1640 292
rect 1648 284 1660 292
rect 1668 284 1720 292
tri 1448 280 1452 284 se
rect 1452 282 1550 284
rect 1578 282 1720 284
rect 1452 280 1460 282
tri 1442 274 1448 280 se
rect 1448 274 1460 280
rect 1468 274 1480 282
rect 1488 274 1500 282
rect 1508 274 1520 282
rect 1528 274 1540 282
rect 1578 274 1590 282
rect 1598 274 1610 282
rect 1618 274 1630 282
rect 1638 274 1650 282
rect 1658 274 1710 282
tri 1436 268 1442 274 se
rect 1442 272 1540 274
rect 1568 272 1710 274
rect 1442 268 1450 272
tri 1430 262 1436 268 se
rect 1436 264 1450 268
rect 1458 264 1470 272
rect 1478 264 1490 272
rect 1498 264 1510 272
rect 1518 264 1530 272
rect 1568 264 1580 272
rect 1588 264 1600 272
rect 1608 264 1620 272
rect 1628 264 1640 272
rect 1648 264 1700 272
rect 1436 262 1530 264
rect 1558 262 1700 264
tri 1424 256 1430 262 se
rect 1430 256 1440 262
tri 1418 250 1424 256 se
rect 1424 254 1440 256
rect 1448 254 1460 262
rect 1468 254 1480 262
rect 1488 254 1500 262
rect 1508 254 1520 262
rect 1558 254 1570 262
rect 1578 254 1590 262
rect 1598 254 1610 262
rect 1618 254 1630 262
rect 1638 254 1690 262
rect 1424 252 1520 254
rect 1548 252 1690 254
rect 1424 250 1430 252
tri 1412 244 1418 250 se
rect 1418 244 1430 250
rect 1438 244 1450 252
rect 1458 244 1470 252
rect 1478 244 1490 252
rect 1498 244 1510 252
rect 1548 244 1560 252
rect 1568 244 1580 252
rect 1588 244 1600 252
rect 1608 244 1620 252
rect 1628 244 1680 252
tri 1408 240 1412 244 se
rect 1412 242 1510 244
rect 1538 242 1680 244
rect 1412 240 1420 242
tri 1402 234 1408 240 se
rect 1408 234 1420 240
rect 1428 234 1440 242
rect 1448 234 1460 242
rect 1468 234 1480 242
rect 1488 234 1500 242
rect 1538 234 1550 242
rect 1558 234 1570 242
rect 1578 234 1590 242
rect 1598 234 1610 242
rect 1618 234 1670 242
tri 1396 228 1402 234 se
rect 1402 232 1500 234
rect 1528 232 1670 234
rect 1402 228 1410 232
tri 1390 222 1396 228 se
rect 1396 224 1410 228
rect 1418 224 1430 232
rect 1438 224 1450 232
rect 1458 224 1470 232
rect 1478 224 1490 232
rect 1528 224 1540 232
rect 1548 224 1560 232
rect 1568 224 1580 232
rect 1588 224 1600 232
rect 1608 224 1660 232
rect 1396 222 1490 224
rect 1518 222 1660 224
tri 1384 216 1390 222 se
rect 1390 216 1400 222
tri 1378 210 1384 216 se
rect 1384 214 1400 216
rect 1408 214 1420 222
rect 1428 214 1440 222
rect 1448 214 1460 222
rect 1468 214 1480 222
rect 1518 214 1530 222
rect 1538 214 1550 222
rect 1558 214 1570 222
rect 1578 214 1590 222
rect 1598 214 1650 222
rect 1384 212 1480 214
rect 1508 212 1650 214
rect 1384 210 1390 212
tri 1374 206 1378 210 se
rect 1378 206 1390 210
tri 1372 204 1374 206 se
rect 1374 204 1390 206
rect 1398 204 1410 212
rect 1418 204 1430 212
rect 1438 204 1450 212
rect 1458 204 1470 212
rect 1508 204 1520 212
rect 1528 204 1540 212
rect 1548 204 1560 212
rect 1568 204 1580 212
rect 1588 204 1640 212
tri 1366 198 1372 204 se
rect 1372 202 1470 204
rect 1498 202 1640 204
rect 1372 198 1380 202
tri 1360 192 1366 198 se
rect 1366 194 1380 198
rect 1388 194 1400 202
rect 1408 194 1420 202
rect 1428 194 1440 202
rect 1448 194 1460 202
rect 1498 194 1510 202
rect 1518 194 1530 202
rect 1538 194 1550 202
rect 1558 194 1570 202
rect 1578 194 1630 202
rect 1366 192 1460 194
rect 1488 192 1630 194
tri 1354 186 1360 192 se
rect 1360 186 1370 192
tri 1350 182 1354 186 se
rect 1354 182 1370 186
rect 1378 182 1390 192
rect 1398 182 1410 192
rect 1418 182 1430 192
rect 1438 182 1450 192
rect 1488 182 1500 192
rect 1508 182 1520 192
rect 1528 182 1540 192
rect 1548 182 1560 192
rect 1568 182 1620 192
tri 1348 180 1350 182 se
rect 1350 180 1360 182
tri 1346 178 1348 180 se
rect 1348 178 1360 180
rect 1346 174 1360 178
rect 1568 174 1610 182
rect 1346 172 1370 174
rect 1346 4 1350 172
rect 1358 144 1370 172
rect 1378 144 1390 174
rect 1358 142 1390 144
rect 1368 134 1380 142
rect 1398 134 1410 174
rect 1418 144 1430 174
rect 1468 144 1480 174
rect 1418 142 1440 144
rect 1428 134 1440 142
rect 1458 142 1480 144
rect 1458 134 1470 142
rect 1488 134 1500 174
rect 1508 142 1520 174
rect 1528 142 1540 174
rect 1548 172 1610 174
rect 1548 162 1600 172
rect 1548 152 1590 162
rect 1548 142 1580 152
rect 1358 132 1380 134
rect 1388 132 1410 134
rect 1418 132 1440 134
rect 1448 132 1470 134
rect 1478 132 1500 134
rect 1358 124 1370 132
rect 1388 124 1400 132
rect 1418 124 1430 132
rect 1448 124 1460 132
rect 1478 124 1490 132
rect 1358 122 1380 124
rect 1388 122 1410 124
rect 1418 122 1440 124
rect 1448 122 1470 124
rect 1478 122 1500 124
rect 1368 114 1380 122
rect 1398 114 1410 122
rect 1428 114 1440 122
rect 1458 114 1470 122
rect 1488 114 1500 122
rect 1358 112 1380 114
rect 1388 112 1410 114
rect 1418 112 1440 114
rect 1448 112 1470 114
rect 1478 112 1500 114
rect 1358 104 1370 112
rect 1388 104 1400 112
rect 1418 104 1430 112
rect 1448 104 1460 112
rect 1478 104 1490 112
rect 1358 102 1380 104
rect 1388 102 1410 104
rect 1418 102 1440 104
rect 1448 102 1470 104
rect 1478 102 1500 104
rect 1368 94 1380 102
rect 1398 94 1410 102
rect 1428 94 1440 102
rect 1458 94 1470 102
rect 1488 94 1500 102
rect 1358 92 1380 94
rect 1388 92 1410 94
rect 1418 92 1440 94
rect 1448 92 1470 94
rect 1478 92 1500 94
rect 1358 84 1370 92
rect 1388 84 1400 92
rect 1418 84 1430 92
rect 1448 84 1460 92
rect 1478 84 1490 92
rect 1358 82 1380 84
rect 1388 82 1410 84
rect 1418 82 1440 84
rect 1448 82 1470 84
rect 1478 82 1500 84
rect 1368 74 1380 82
rect 1398 74 1410 82
rect 1428 74 1440 82
rect 1458 74 1470 82
rect 1488 74 1500 82
rect 1358 72 1380 74
rect 1388 72 1410 74
rect 1418 72 1440 74
rect 1448 72 1470 74
rect 1478 72 1500 74
rect 1358 64 1370 72
rect 1388 64 1400 72
rect 1418 64 1430 72
rect 1448 64 1460 72
rect 1478 64 1490 72
rect 1358 62 1380 64
rect 1388 62 1410 64
rect 1418 62 1440 64
rect 1448 62 1470 64
rect 1478 62 1500 64
rect 1368 54 1380 62
rect 1398 54 1410 62
rect 1428 54 1440 62
rect 1458 54 1470 62
rect 1488 54 1500 62
rect 1358 52 1380 54
rect 1388 52 1410 54
rect 1418 52 1440 54
rect 1448 52 1470 54
rect 1478 52 1500 54
rect 1358 44 1370 52
rect 1388 44 1400 52
rect 1418 44 1430 52
rect 1448 44 1460 52
rect 1478 44 1490 52
rect 1358 42 1380 44
rect 1388 42 1410 44
rect 1418 42 1440 44
rect 1448 42 1470 44
rect 1478 42 1500 44
rect 1368 34 1380 42
rect 1398 34 1410 42
rect 1428 34 1440 42
rect 1458 34 1470 42
rect 1488 34 1500 42
rect 1358 32 1380 34
rect 1388 32 1410 34
rect 1418 32 1440 34
rect 1448 32 1470 34
rect 1478 32 1500 34
rect 1358 24 1370 32
rect 1388 24 1400 32
rect 1418 24 1430 32
rect 1448 24 1460 32
rect 1478 24 1490 32
rect 1358 22 1380 24
rect 1388 22 1410 24
rect 1418 22 1440 24
rect 1448 22 1470 24
rect 1478 22 1500 24
rect 1368 14 1380 22
rect 1398 14 1410 22
rect 1428 14 1440 22
rect 1458 14 1470 22
rect 1488 14 1500 22
rect 1358 12 1380 14
rect 1388 12 1410 14
rect 1418 12 1440 14
rect 1448 12 1470 14
rect 1478 12 1500 14
rect 1358 4 1370 12
rect 1388 4 1400 12
rect 1418 4 1430 12
rect 1448 4 1460 12
rect 1478 4 1490 12
rect 1998 4 2000 502
rect 1346 0 2000 4
<< psubstratepcontact >>
rect 1584 1322 1992 1332
rect 1574 1312 1992 1322
rect 1564 1302 1992 1312
rect 1554 1292 1992 1302
rect 1544 1282 1992 1292
rect 1534 1272 1992 1282
rect 1524 1262 1992 1272
rect 1514 1252 1992 1262
rect 1504 1242 1992 1252
rect 1494 1232 1992 1242
rect 1484 1222 1992 1232
rect 1474 1212 1992 1222
rect 1464 1202 1992 1212
rect 1454 1192 1992 1202
rect 1444 1182 1992 1192
rect 1434 1172 1992 1182
rect 1424 1162 1992 1172
rect 1414 1152 1992 1162
rect 1404 1142 1992 1152
rect 1394 1132 1992 1142
rect 1384 1122 1992 1132
rect 1374 1112 1992 1122
rect 1364 1102 1992 1112
rect 1354 1092 1992 1102
rect 1344 1082 1992 1092
rect 1334 1072 1992 1082
rect 1324 1062 1992 1072
rect 1314 1054 1992 1062
rect 1314 1052 1572 1054
rect 1304 1044 1572 1052
rect 1304 1042 1562 1044
rect 1294 1034 1562 1042
rect 1294 1032 1552 1034
rect 1284 1024 1552 1032
rect 1284 1022 1542 1024
rect 1594 1022 1992 1054
rect 1274 1014 1542 1022
rect 1274 1012 1532 1014
rect 1584 1012 1992 1022
rect 1264 1004 1532 1012
rect 1264 1002 1522 1004
rect 1574 1002 1992 1012
rect 1254 994 1522 1002
rect 1254 992 1512 994
rect 1564 992 1992 1002
rect 1244 984 1512 992
rect 1244 982 1502 984
rect 1554 982 1992 992
rect 1234 974 1502 982
rect 1234 972 1492 974
rect 1544 972 1992 982
rect 1224 964 1492 972
rect 1224 962 1482 964
rect 1534 962 1992 972
rect 1214 954 1482 962
rect 1214 952 1472 954
rect 1524 952 1992 962
rect 1204 944 1472 952
rect 1204 942 1462 944
rect 1514 942 1992 952
rect 1194 934 1462 942
rect 1194 932 1452 934
rect 1504 932 1992 942
rect 1184 924 1452 932
rect 1184 922 1442 924
rect 1494 922 1992 932
rect 1174 914 1442 922
rect 1174 912 1432 914
rect 1484 912 1992 922
rect 1164 904 1432 912
rect 1164 902 1422 904
rect 1474 902 1992 912
rect 1154 894 1422 902
rect 1154 892 1412 894
rect 1464 892 1992 902
rect 1144 884 1412 892
rect 1454 884 1992 892
rect 1144 882 1402 884
rect 1454 882 1702 884
rect 1134 874 1402 882
rect 1444 874 1702 882
rect 1134 872 1392 874
rect 1444 872 1692 874
rect 1124 864 1392 872
rect 1434 864 1692 872
rect 1124 862 1382 864
rect 1434 862 1682 864
rect 1734 862 1992 884
rect 1114 854 1382 862
rect 1424 854 1682 862
rect 1114 852 1372 854
rect 1424 852 1672 854
rect 1724 852 1992 862
rect 1104 844 1372 852
rect 1414 844 1672 852
rect 1714 844 1992 852
rect 1104 842 1362 844
rect 1414 842 1662 844
rect 1714 842 1722 844
rect 1094 834 1362 842
rect 1404 834 1662 842
rect 1094 832 1352 834
rect 1404 832 1652 834
rect 1704 832 1722 842
rect 1734 834 1752 844
rect 1764 834 1782 844
rect 1794 834 1812 844
rect 1824 834 1842 844
rect 1854 834 1872 844
rect 1884 834 1902 844
rect 1914 834 1932 844
rect 1944 834 1962 844
rect 1974 834 1992 844
rect 1744 832 1752 834
rect 1774 832 1782 834
rect 1804 832 1812 834
rect 1834 832 1842 834
rect 1864 832 1872 834
rect 1894 832 1902 834
rect 1924 832 1932 834
rect 1954 832 1962 834
rect 1084 824 1352 832
rect 1394 824 1652 832
rect 1694 824 1732 832
rect 1744 824 1762 832
rect 1774 824 1792 832
rect 1804 824 1822 832
rect 1834 824 1852 832
rect 1864 824 1882 832
rect 1894 824 1912 832
rect 1924 824 1942 832
rect 1954 824 1972 832
rect 1084 822 1342 824
rect 1394 822 1642 824
rect 1694 822 1722 824
rect 1744 822 1752 824
rect 1774 822 1782 824
rect 1804 822 1812 824
rect 1834 822 1842 824
rect 1864 822 1872 824
rect 1894 822 1902 824
rect 1924 822 1932 824
rect 1954 822 1962 824
rect 1984 822 1992 834
rect 1074 814 1342 822
rect 1384 814 1642 822
rect 1684 814 1722 822
rect 1734 814 1752 822
rect 1764 814 1782 822
rect 1794 814 1812 822
rect 1824 814 1842 822
rect 1854 814 1872 822
rect 1884 814 1902 822
rect 1914 814 1932 822
rect 1944 814 1962 822
rect 1974 814 1992 822
rect 1074 812 1332 814
rect 1384 812 1632 814
rect 1684 812 1692 814
rect 1064 804 1332 812
rect 1374 804 1632 812
rect 1674 804 1692 812
rect 1704 812 1722 814
rect 1744 812 1752 814
rect 1774 812 1782 814
rect 1804 812 1812 814
rect 1834 812 1842 814
rect 1864 812 1872 814
rect 1894 812 1902 814
rect 1924 812 1932 814
rect 1954 812 1962 814
rect 1704 804 1732 812
rect 1744 804 1762 812
rect 1774 804 1792 812
rect 1804 804 1822 812
rect 1834 804 1852 812
rect 1864 804 1882 812
rect 1894 804 1912 812
rect 1924 804 1942 812
rect 1954 804 1972 812
rect 1064 802 1322 804
rect 1374 802 1622 804
rect 1674 802 1682 804
rect 1704 802 1722 804
rect 1744 802 1752 804
rect 1774 802 1782 804
rect 1804 802 1812 804
rect 1834 802 1842 804
rect 1864 802 1872 804
rect 1894 802 1902 804
rect 1924 802 1932 804
rect 1954 802 1962 804
rect 1984 802 1992 814
rect 1054 794 1322 802
rect 1364 794 1622 802
rect 1664 794 1682 802
rect 1694 794 1722 802
rect 1734 794 1752 802
rect 1764 794 1782 802
rect 1794 794 1812 802
rect 1824 794 1842 802
rect 1854 794 1872 802
rect 1884 794 1902 802
rect 1914 794 1932 802
rect 1944 794 1962 802
rect 1974 794 1992 802
rect 1054 792 1312 794
rect 1364 792 1612 794
rect 1664 792 1672 794
rect 1704 792 1722 794
rect 1744 792 1752 794
rect 1774 792 1782 794
rect 1804 792 1812 794
rect 1834 792 1842 794
rect 1864 792 1872 794
rect 1894 792 1902 794
rect 1924 792 1932 794
rect 1954 792 1962 794
rect 1044 784 1312 792
rect 1354 784 1612 792
rect 1654 784 1672 792
rect 1684 784 1692 792
rect 1704 784 1732 792
rect 1744 784 1762 792
rect 1774 784 1792 792
rect 1804 784 1822 792
rect 1834 784 1852 792
rect 1864 784 1882 792
rect 1894 784 1912 792
rect 1924 784 1942 792
rect 1954 784 1972 792
rect 1044 782 1302 784
rect 1354 782 1602 784
rect 1654 782 1662 784
rect 1704 782 1722 784
rect 1744 782 1752 784
rect 1774 782 1782 784
rect 1804 782 1812 784
rect 1834 782 1842 784
rect 1864 782 1872 784
rect 1894 782 1902 784
rect 1924 782 1932 784
rect 1954 782 1962 784
rect 1984 782 1992 794
rect 1034 774 1302 782
rect 1344 774 1602 782
rect 1644 774 1662 782
rect 1674 774 1682 782
rect 1034 772 1292 774
rect 1344 772 1592 774
rect 1644 772 1652 774
rect 1694 772 1722 782
rect 1734 774 1752 782
rect 1764 774 1782 782
rect 1794 774 1812 782
rect 1824 774 1842 782
rect 1854 774 1872 782
rect 1884 774 1902 782
rect 1914 774 1932 782
rect 1944 774 1962 782
rect 1974 774 1992 782
rect 1744 772 1752 774
rect 1774 772 1782 774
rect 1804 772 1812 774
rect 1834 772 1842 774
rect 1864 772 1872 774
rect 1894 772 1902 774
rect 1924 772 1932 774
rect 1954 772 1962 774
rect 1024 764 1292 772
rect 1334 764 1592 772
rect 1634 764 1652 772
rect 1664 764 1672 772
rect 1684 764 1732 772
rect 1744 764 1762 772
rect 1774 764 1792 772
rect 1804 764 1822 772
rect 1834 764 1852 772
rect 1864 764 1882 772
rect 1894 764 1912 772
rect 1924 764 1942 772
rect 1954 764 1972 772
rect 1024 762 1282 764
rect 1334 762 1582 764
rect 1634 762 1642 764
rect 1684 762 1692 764
rect 1014 754 1282 762
rect 1324 754 1582 762
rect 1624 754 1642 762
rect 1654 754 1662 762
rect 1674 754 1692 762
rect 1014 752 1272 754
rect 1324 752 1572 754
rect 1624 752 1632 754
rect 1674 752 1682 754
rect 1704 752 1722 764
rect 1744 762 1752 764
rect 1774 762 1782 764
rect 1804 762 1812 764
rect 1834 762 1842 764
rect 1864 762 1872 764
rect 1894 762 1902 764
rect 1924 762 1932 764
rect 1954 762 1962 764
rect 1984 762 1992 774
rect 1734 754 1752 762
rect 1764 754 1782 762
rect 1794 754 1812 762
rect 1824 754 1842 762
rect 1854 754 1872 762
rect 1884 754 1902 762
rect 1914 754 1932 762
rect 1944 754 1962 762
rect 1974 754 1992 762
rect 1744 752 1752 754
rect 1774 752 1782 754
rect 1804 752 1812 754
rect 1834 752 1842 754
rect 1864 752 1872 754
rect 1894 752 1902 754
rect 1924 752 1932 754
rect 1954 752 1962 754
rect 1004 744 1272 752
rect 1314 744 1572 752
rect 1614 744 1632 752
rect 1644 744 1652 752
rect 1664 744 1682 752
rect 1694 744 1732 752
rect 1744 744 1762 752
rect 1774 744 1792 752
rect 1804 744 1822 752
rect 1834 744 1852 752
rect 1864 744 1882 752
rect 1894 744 1912 752
rect 1924 744 1942 752
rect 1954 744 1972 752
rect 1004 742 1262 744
rect 1314 742 1562 744
rect 1614 742 1622 744
rect 1664 742 1672 744
rect 1694 742 1722 744
rect 1744 742 1752 744
rect 1774 742 1782 744
rect 1804 742 1812 744
rect 1834 742 1842 744
rect 1864 742 1872 744
rect 1894 742 1902 744
rect 1924 742 1932 744
rect 1954 742 1962 744
rect 1984 742 1992 754
rect 994 734 1262 742
rect 1304 734 1562 742
rect 1604 734 1622 742
rect 1634 734 1642 742
rect 1654 734 1672 742
rect 994 732 1252 734
rect 1304 732 1552 734
rect 1604 732 1612 734
rect 1654 732 1662 734
rect 1684 732 1722 742
rect 1734 734 1752 742
rect 1764 734 1782 742
rect 1794 734 1812 742
rect 1824 734 1842 742
rect 1854 734 1872 742
rect 1884 734 1902 742
rect 1914 734 1932 742
rect 1944 734 1962 742
rect 1974 734 1992 742
rect 1744 732 1752 734
rect 1774 732 1782 734
rect 1804 732 1812 734
rect 1834 732 1842 734
rect 1864 732 1872 734
rect 1894 732 1902 734
rect 1924 732 1932 734
rect 1954 732 1962 734
rect 984 724 1252 732
rect 1294 724 1552 732
rect 1594 724 1612 732
rect 1624 724 1632 732
rect 1644 724 1662 732
rect 1674 724 1732 732
rect 1744 724 1762 732
rect 1774 724 1792 732
rect 1804 724 1822 732
rect 1834 724 1852 732
rect 1864 724 1882 732
rect 1894 724 1912 732
rect 1924 724 1942 732
rect 1954 724 1972 732
rect 984 722 1242 724
rect 1294 722 1542 724
rect 1594 722 1602 724
rect 1644 722 1652 724
rect 1674 722 1722 724
rect 1744 722 1752 724
rect 1774 722 1782 724
rect 1804 722 1812 724
rect 1834 722 1842 724
rect 1864 722 1872 724
rect 1894 722 1902 724
rect 1924 722 1932 724
rect 1954 722 1962 724
rect 1984 722 1992 734
rect 974 714 1242 722
rect 1284 714 1542 722
rect 1584 714 1602 722
rect 1614 714 1622 722
rect 1634 714 1652 722
rect 974 712 1232 714
rect 1284 712 1532 714
rect 1584 712 1592 714
rect 1634 712 1642 714
rect 1664 712 1722 722
rect 1734 714 1752 722
rect 1764 714 1782 722
rect 1794 714 1812 722
rect 1824 714 1842 722
rect 1854 714 1872 722
rect 1884 714 1902 722
rect 1914 714 1932 722
rect 1944 714 1962 722
rect 1974 714 1992 722
rect 1744 712 1752 714
rect 1774 712 1782 714
rect 1804 712 1812 714
rect 1834 712 1842 714
rect 1864 712 1872 714
rect 1894 712 1902 714
rect 1924 712 1932 714
rect 1954 712 1962 714
rect 964 704 1232 712
rect 1274 704 1532 712
rect 1574 704 1592 712
rect 1604 704 1612 712
rect 1624 704 1642 712
rect 1654 704 1732 712
rect 1744 704 1762 712
rect 1774 704 1792 712
rect 1804 704 1822 712
rect 1834 704 1852 712
rect 1864 704 1882 712
rect 1894 704 1912 712
rect 1924 704 1942 712
rect 1954 704 1972 712
rect 964 702 1222 704
rect 1274 702 1522 704
rect 1574 702 1582 704
rect 1624 702 1632 704
rect 1654 702 1692 704
rect 954 694 1222 702
rect 1264 694 1522 702
rect 1564 694 1582 702
rect 1594 694 1602 702
rect 1614 694 1632 702
rect 954 692 1212 694
rect 1264 692 1512 694
rect 1564 692 1572 694
rect 944 684 1212 692
rect 1254 684 1512 692
rect 1554 684 1572 692
rect 1584 684 1592 692
rect 1604 684 1612 692
rect 1624 684 1632 694
rect 1644 694 1692 702
rect 1704 694 1722 704
rect 1744 702 1752 704
rect 1774 702 1782 704
rect 1804 702 1812 704
rect 1834 702 1842 704
rect 1864 702 1872 704
rect 1894 702 1902 704
rect 1924 702 1932 704
rect 1954 702 1962 704
rect 1984 702 1992 714
rect 1644 684 1682 694
rect 1694 684 1702 692
rect 1714 684 1722 694
rect 1734 694 1752 702
rect 1764 694 1782 702
rect 1794 694 1812 702
rect 1824 694 1842 702
rect 1854 694 1872 702
rect 1884 694 1902 702
rect 1914 694 1932 702
rect 1944 694 1962 702
rect 1974 694 1992 702
rect 1734 684 1742 694
rect 1754 684 1762 692
rect 1774 684 1782 694
rect 944 682 1202 684
rect 1254 682 1502 684
rect 1554 682 1562 684
rect 1644 682 1672 684
rect 934 674 1202 682
rect 1244 674 1502 682
rect 1544 674 1562 682
rect 1574 674 1582 682
rect 1594 674 1602 682
rect 1614 674 1622 682
rect 1634 674 1672 682
rect 1684 674 1692 682
rect 1704 674 1712 682
rect 1724 674 1732 682
rect 1744 674 1752 682
rect 1764 674 1772 682
rect 934 672 1192 674
rect 1244 672 1492 674
rect 1544 672 1552 674
rect 1634 672 1662 674
rect 924 664 1192 672
rect 1234 664 1492 672
rect 1534 664 1552 672
rect 1564 664 1572 672
rect 1584 664 1592 672
rect 1604 664 1612 672
rect 1624 664 1662 672
rect 1674 664 1682 672
rect 1694 664 1702 672
rect 1714 664 1722 672
rect 1734 664 1742 672
rect 1754 664 1762 672
rect 924 662 1182 664
rect 1234 662 1482 664
rect 1534 662 1542 664
rect 1624 662 1652 664
rect 914 654 1182 662
rect 1224 654 1482 662
rect 1524 654 1542 662
rect 1554 654 1562 662
rect 1574 654 1582 662
rect 1594 654 1602 662
rect 1614 654 1652 662
rect 1664 654 1672 662
rect 1684 654 1692 662
rect 1704 654 1712 662
rect 1724 654 1732 662
rect 1744 654 1752 662
rect 914 652 1172 654
rect 1224 652 1472 654
rect 1524 652 1532 654
rect 1614 652 1642 654
rect 904 644 1172 652
rect 1214 644 1472 652
rect 1514 644 1532 652
rect 1544 644 1552 652
rect 1564 644 1572 652
rect 1584 644 1592 652
rect 1604 644 1642 652
rect 1654 644 1662 652
rect 1674 644 1682 652
rect 1694 644 1702 652
rect 1714 644 1722 652
rect 1734 644 1742 652
rect 904 642 1162 644
rect 1214 642 1462 644
rect 1514 642 1522 644
rect 1604 642 1632 644
rect 894 634 1162 642
rect 1204 634 1462 642
rect 1504 634 1522 642
rect 1534 634 1542 642
rect 1554 634 1562 642
rect 1574 634 1582 642
rect 1594 634 1632 642
rect 1644 634 1652 642
rect 1664 634 1672 642
rect 1684 634 1692 642
rect 1704 634 1712 642
rect 1724 634 1732 642
rect 894 632 1152 634
rect 1204 632 1452 634
rect 1504 632 1512 634
rect 1594 632 1622 634
rect 884 624 1152 632
rect 1194 624 1452 632
rect 1494 624 1512 632
rect 1524 624 1532 632
rect 1544 624 1552 632
rect 1564 624 1572 632
rect 1584 624 1622 632
rect 1634 624 1642 632
rect 1654 624 1662 632
rect 1674 624 1682 632
rect 1694 624 1702 632
rect 1714 624 1722 632
rect 884 622 1142 624
rect 1194 622 1442 624
rect 1494 622 1502 624
rect 1584 622 1612 624
rect 874 614 1142 622
rect 1184 614 1442 622
rect 1484 614 1502 622
rect 1514 614 1522 622
rect 1534 614 1542 622
rect 1554 614 1562 622
rect 1574 614 1612 622
rect 1624 614 1632 622
rect 1644 614 1652 622
rect 1664 614 1672 622
rect 1684 614 1692 622
rect 1704 614 1712 622
rect 874 612 1132 614
rect 1184 612 1432 614
rect 1484 612 1492 614
rect 1574 612 1602 614
rect 864 604 1132 612
rect 1174 604 1432 612
rect 1474 604 1492 612
rect 1504 604 1512 612
rect 1524 604 1532 612
rect 1544 604 1552 612
rect 1564 604 1602 612
rect 1614 604 1622 612
rect 1634 604 1642 612
rect 1654 604 1662 612
rect 1674 604 1682 612
rect 1694 604 1702 612
rect 864 602 1122 604
rect 1174 602 1422 604
rect 1474 602 1482 604
rect 1564 602 1592 604
rect 854 594 1122 602
rect 1164 594 1422 602
rect 1464 594 1482 602
rect 1494 594 1502 602
rect 1514 594 1522 602
rect 1534 594 1542 602
rect 1554 594 1592 602
rect 1604 594 1612 602
rect 1624 594 1632 602
rect 1644 594 1652 602
rect 1664 594 1672 602
rect 1684 594 1692 602
rect 854 592 1112 594
rect 1164 592 1412 594
rect 1464 592 1472 594
rect 1554 592 1582 594
rect 844 584 1112 592
rect 1154 584 1412 592
rect 1454 584 1472 592
rect 1484 584 1492 592
rect 1504 584 1512 592
rect 1524 584 1532 592
rect 1544 584 1582 592
rect 1594 584 1602 592
rect 1614 584 1622 592
rect 1634 584 1642 592
rect 1654 584 1662 592
rect 1674 584 1682 592
rect 844 582 1102 584
rect 1154 582 1402 584
rect 1454 582 1462 584
rect 1544 582 1572 584
rect 834 574 1102 582
rect 1144 574 1402 582
rect 1444 574 1462 582
rect 1474 574 1482 582
rect 1494 574 1502 582
rect 1514 574 1522 582
rect 1534 574 1572 582
rect 1584 574 1592 582
rect 1604 574 1612 582
rect 1624 574 1632 582
rect 1644 574 1652 582
rect 1664 574 1672 582
rect 834 572 1092 574
rect 1144 572 1392 574
rect 1444 572 1452 574
rect 1534 572 1562 574
rect 824 564 1092 572
rect 1134 564 1392 572
rect 1434 564 1452 572
rect 1464 564 1472 572
rect 1484 564 1492 572
rect 1504 564 1512 572
rect 1524 564 1562 572
rect 1574 564 1582 572
rect 1594 564 1602 572
rect 1614 564 1622 572
rect 1634 564 1642 572
rect 1654 564 1662 572
rect 824 562 1082 564
rect 1134 562 1382 564
rect 1434 562 1442 564
rect 1524 562 1552 564
rect 814 554 1082 562
rect 1124 554 1382 562
rect 1424 554 1442 562
rect 1454 554 1462 562
rect 1474 554 1482 562
rect 1494 554 1502 562
rect 1514 554 1552 562
rect 1564 554 1572 562
rect 1584 554 1592 562
rect 1604 554 1612 562
rect 1624 554 1632 562
rect 1644 554 1652 562
rect 814 552 1072 554
rect 1124 552 1372 554
rect 1424 552 1432 554
rect 1514 552 1542 554
rect 804 544 1072 552
rect 1114 544 1372 552
rect 1414 544 1432 552
rect 1444 544 1452 552
rect 1464 544 1472 552
rect 1484 544 1492 552
rect 1504 544 1542 552
rect 1554 544 1562 552
rect 1574 544 1582 552
rect 1594 544 1602 552
rect 1614 544 1622 552
rect 1634 544 1642 552
rect 804 542 1062 544
rect 1114 542 1362 544
rect 1414 542 1422 544
rect 1504 542 1532 544
rect 794 534 1062 542
rect 1104 534 1362 542
rect 1404 534 1422 542
rect 1434 534 1442 542
rect 1454 534 1462 542
rect 1474 534 1482 542
rect 1494 534 1532 542
rect 1544 534 1552 542
rect 1564 534 1572 542
rect 1584 534 1592 542
rect 1604 534 1612 542
rect 1624 534 1632 542
rect 794 532 1052 534
rect 1104 532 1352 534
rect 1404 532 1412 534
rect 1494 532 1522 534
rect 784 524 1052 532
rect 1094 524 1352 532
rect 1394 524 1412 532
rect 1424 524 1432 532
rect 1444 524 1452 532
rect 1464 524 1472 532
rect 1484 524 1522 532
rect 1534 524 1542 532
rect 1554 524 1562 532
rect 1574 524 1582 532
rect 1594 524 1602 532
rect 1614 524 1622 532
rect 784 522 1042 524
rect 1094 522 1342 524
rect 1394 522 1402 524
rect 1484 522 1512 524
rect 774 514 1042 522
rect 1084 514 1342 522
rect 1384 514 1402 522
rect 1414 514 1422 522
rect 1434 514 1442 522
rect 1454 514 1462 522
rect 1474 514 1512 522
rect 1524 514 1532 522
rect 1544 514 1552 522
rect 1564 514 1572 522
rect 1584 514 1592 522
rect 1604 514 1612 522
rect 774 512 1032 514
rect 1084 512 1332 514
rect 1384 512 1392 514
rect 1474 512 1502 514
rect 764 504 1032 512
rect 1074 504 1332 512
rect 1374 504 1392 512
rect 1404 504 1412 512
rect 1424 504 1432 512
rect 1444 504 1452 512
rect 1464 504 1502 512
rect 1514 504 1522 512
rect 1534 504 1542 512
rect 1554 504 1562 512
rect 1574 504 1582 512
rect 1594 504 1602 512
rect 764 502 1022 504
rect 1074 502 1322 504
rect 1374 502 1382 504
rect 1464 502 1492 504
rect 754 494 1022 502
rect 1064 494 1322 502
rect 1364 494 1382 502
rect 1394 494 1402 502
rect 1414 494 1422 502
rect 1434 494 1442 502
rect 1454 494 1492 502
rect 1504 494 1512 502
rect 1524 494 1532 502
rect 1544 494 1552 502
rect 1564 494 1572 502
rect 1584 494 1592 502
rect 754 492 1012 494
rect 1064 492 1312 494
rect 1364 492 1372 494
rect 1454 492 1482 494
rect 744 484 1012 492
rect 1054 484 1312 492
rect 1354 484 1372 492
rect 1384 484 1392 492
rect 1404 484 1412 492
rect 1424 484 1432 492
rect 1444 484 1482 492
rect 1494 484 1502 492
rect 1514 484 1522 492
rect 1534 484 1542 492
rect 1554 484 1562 492
rect 1574 484 1582 492
rect 744 482 1002 484
rect 1054 482 1302 484
rect 1354 482 1362 484
rect 1444 482 1472 484
rect 734 474 1002 482
rect 1044 474 1302 482
rect 1344 474 1362 482
rect 1374 474 1382 482
rect 1394 474 1402 482
rect 1414 474 1422 482
rect 1434 474 1472 482
rect 1484 474 1492 482
rect 1504 474 1512 482
rect 1524 474 1532 482
rect 1544 474 1552 482
rect 1564 474 1572 482
rect 734 472 992 474
rect 1044 472 1292 474
rect 1344 472 1352 474
rect 1434 472 1462 474
rect 724 464 992 472
rect 1034 464 1292 472
rect 1334 464 1352 472
rect 1364 464 1372 472
rect 1384 464 1392 472
rect 1404 464 1412 472
rect 1424 464 1462 472
rect 1474 464 1482 472
rect 1494 464 1502 472
rect 1514 464 1522 472
rect 1534 464 1542 472
rect 1554 464 1562 472
rect 724 462 982 464
rect 1034 462 1282 464
rect 1334 462 1342 464
rect 1424 462 1452 464
rect 714 454 982 462
rect 1024 454 1282 462
rect 1324 454 1342 462
rect 1354 454 1362 462
rect 1374 454 1382 462
rect 1394 454 1402 462
rect 1414 454 1452 462
rect 1464 454 1472 462
rect 1484 454 1492 462
rect 1504 454 1512 462
rect 1524 454 1532 462
rect 1544 454 1552 462
rect 714 452 972 454
rect 1024 452 1272 454
rect 1324 452 1332 454
rect 1414 452 1442 454
rect 704 444 972 452
rect 1014 444 1272 452
rect 1314 444 1332 452
rect 1344 444 1352 452
rect 1364 444 1372 452
rect 1384 444 1392 452
rect 1404 444 1442 452
rect 1454 444 1462 452
rect 1474 444 1482 452
rect 1494 444 1502 452
rect 1514 444 1522 452
rect 1534 444 1542 452
rect 704 442 962 444
rect 1014 442 1262 444
rect 1314 442 1322 444
rect 1404 442 1432 444
rect 694 434 962 442
rect 1004 434 1262 442
rect 1304 434 1322 442
rect 1334 434 1342 442
rect 1354 434 1362 442
rect 1374 434 1382 442
rect 1394 434 1432 442
rect 1444 434 1452 442
rect 1464 434 1472 442
rect 1484 434 1492 442
rect 1504 434 1512 442
rect 1524 434 1532 442
rect 694 432 952 434
rect 1004 432 1252 434
rect 1304 432 1312 434
rect 1394 432 1422 434
rect 684 424 952 432
rect 994 424 1252 432
rect 1294 424 1312 432
rect 1324 424 1332 432
rect 1344 424 1352 432
rect 1364 424 1372 432
rect 1384 424 1422 432
rect 1434 424 1442 432
rect 1454 424 1462 432
rect 1474 424 1482 432
rect 1494 424 1502 432
rect 1514 424 1522 432
rect 684 422 942 424
rect 994 422 1242 424
rect 1294 422 1302 424
rect 1384 422 1412 424
rect 674 414 942 422
rect 984 414 1242 422
rect 1284 414 1302 422
rect 1314 414 1322 422
rect 1334 414 1342 422
rect 1354 414 1362 422
rect 1374 414 1412 422
rect 1424 414 1432 422
rect 1444 414 1452 422
rect 1464 414 1472 422
rect 1484 414 1492 422
rect 1504 414 1512 422
rect 674 412 932 414
rect 984 412 1232 414
rect 1284 412 1292 414
rect 1374 412 1402 414
rect 664 382 932 412
rect 974 404 1232 412
rect 1274 404 1292 412
rect 1304 404 1312 412
rect 1324 404 1332 412
rect 1344 404 1352 412
rect 1364 404 1402 412
rect 1414 404 1422 412
rect 1434 404 1442 412
rect 1454 404 1462 412
rect 1474 404 1482 412
rect 1494 404 1502 412
rect 974 402 1222 404
rect 1274 402 1282 404
rect 1364 402 1392 404
rect 964 394 1222 402
rect 1264 394 1282 402
rect 1294 394 1302 402
rect 1314 394 1322 402
rect 1334 394 1342 402
rect 1354 394 1392 402
rect 1404 394 1412 402
rect 1424 394 1432 402
rect 1444 394 1452 402
rect 1464 394 1472 402
rect 1484 394 1492 402
rect 964 392 1212 394
rect 1264 392 1272 394
rect 1354 392 1382 394
rect 954 384 1212 392
rect 1254 384 1272 392
rect 1284 384 1292 392
rect 1304 384 1312 392
rect 1324 384 1332 392
rect 1344 384 1382 392
rect 1394 384 1402 392
rect 1414 384 1422 392
rect 1434 384 1442 392
rect 1454 384 1462 392
rect 1474 384 1482 392
rect 954 382 1202 384
rect 1254 382 1262 384
rect 1344 382 1372 384
rect 664 374 1202 382
rect 1244 374 1262 382
rect 1274 374 1282 382
rect 1294 374 1302 382
rect 1314 374 1322 382
rect 1334 374 1372 382
rect 1384 374 1392 382
rect 1404 374 1412 382
rect 1424 374 1432 382
rect 1444 374 1452 382
rect 1464 374 1472 382
rect 664 364 1192 374
rect 1244 372 1252 374
rect 1334 372 1362 374
rect 1234 364 1252 372
rect 1264 364 1272 372
rect 1284 364 1292 372
rect 1304 364 1312 372
rect 1324 364 1362 372
rect 1374 364 1382 372
rect 1394 364 1402 372
rect 1414 364 1422 372
rect 1434 364 1442 372
rect 1454 364 1462 372
rect 664 354 1182 364
rect 1234 362 1242 364
rect 1324 362 1352 364
rect 1224 354 1242 362
rect 1254 354 1262 362
rect 1274 354 1282 362
rect 1294 354 1302 362
rect 1314 354 1352 362
rect 1364 354 1372 362
rect 1384 354 1392 362
rect 1404 354 1412 362
rect 1424 354 1432 362
rect 1444 354 1452 362
rect 664 344 1172 354
rect 1224 352 1232 354
rect 1314 352 1342 354
rect 1214 344 1232 352
rect 1244 344 1252 352
rect 1264 344 1272 352
rect 1284 344 1292 352
rect 1304 344 1342 352
rect 1354 344 1362 352
rect 1374 344 1382 352
rect 1394 344 1402 352
rect 1414 344 1422 352
rect 1434 344 1442 352
rect 664 334 1162 344
rect 1214 342 1222 344
rect 1304 342 1332 344
rect 1204 334 1222 342
rect 1234 334 1242 342
rect 1254 334 1262 342
rect 1274 334 1282 342
rect 1294 334 1332 342
rect 1344 334 1352 342
rect 1364 334 1372 342
rect 1384 334 1392 342
rect 1404 334 1412 342
rect 1424 334 1432 342
rect 664 324 1152 334
rect 1204 332 1212 334
rect 1294 332 1322 334
rect 1194 324 1212 332
rect 1224 324 1232 332
rect 1244 324 1252 332
rect 1264 324 1272 332
rect 1284 324 1322 332
rect 1334 324 1342 332
rect 1354 324 1362 332
rect 1374 324 1382 332
rect 1394 324 1402 332
rect 1414 324 1422 332
rect 664 314 1142 324
rect 1194 322 1202 324
rect 1284 322 1312 324
rect 1184 314 1202 322
rect 1214 314 1222 322
rect 1234 314 1242 322
rect 1254 314 1262 322
rect 1274 314 1312 322
rect 1324 314 1332 322
rect 1344 314 1352 322
rect 1364 314 1372 322
rect 1384 314 1392 322
rect 1404 314 1412 322
rect 664 304 1132 314
rect 1184 312 1192 314
rect 1274 312 1302 314
rect 1174 304 1192 312
rect 1204 304 1212 312
rect 1224 304 1232 312
rect 1244 304 1252 312
rect 1264 304 1302 312
rect 1314 304 1322 312
rect 1334 304 1342 312
rect 1354 304 1362 312
rect 1374 304 1382 312
rect 1394 304 1402 312
rect 664 294 1122 304
rect 1174 302 1182 304
rect 1264 302 1292 304
rect 1164 294 1182 302
rect 1194 294 1202 302
rect 1214 294 1222 302
rect 1234 294 1242 302
rect 1254 294 1292 302
rect 1304 294 1312 302
rect 1324 294 1332 302
rect 1344 294 1352 302
rect 1364 294 1372 302
rect 1384 294 1392 302
rect 664 274 1112 294
rect 1164 292 1172 294
rect 1254 292 1282 294
rect 1154 284 1172 292
rect 1184 284 1192 292
rect 1204 284 1212 292
rect 1224 284 1232 292
rect 1244 284 1282 292
rect 1294 284 1302 292
rect 1314 284 1322 292
rect 1334 284 1342 292
rect 1354 284 1362 292
rect 1374 284 1382 292
rect 1154 282 1162 284
rect 1244 282 1272 284
rect 1144 274 1162 282
rect 1174 274 1182 282
rect 1194 274 1202 282
rect 1214 274 1222 282
rect 1234 274 1272 282
rect 1284 274 1292 282
rect 1304 274 1312 282
rect 1324 274 1332 282
rect 1344 274 1352 282
rect 1364 274 1372 282
rect 664 242 1092 274
rect 1144 272 1152 274
rect 1234 272 1262 274
rect 1134 242 1152 272
rect 1164 244 1172 272
rect 1184 262 1192 272
rect 1204 264 1212 272
rect 1224 264 1262 272
rect 1224 262 1232 264
rect 1184 244 1202 262
rect 1214 244 1232 262
rect 1244 244 1262 264
rect 1274 262 1282 272
rect 1294 264 1302 272
rect 1314 262 1322 272
rect 1274 244 1292 262
rect 1304 244 1322 262
rect 1334 262 1342 272
rect 1354 264 1362 272
rect 1334 254 1352 262
rect 1334 244 1342 254
rect 1184 242 1192 244
rect 1214 242 1222 244
rect 1244 242 1252 244
rect 1274 242 1282 244
rect 1304 242 1312 244
rect 664 232 1162 242
rect 1174 234 1192 242
rect 1204 234 1222 242
rect 1234 234 1252 242
rect 1264 234 1282 242
rect 1294 234 1312 242
rect 1324 234 1332 242
rect 1184 232 1192 234
rect 1214 232 1222 234
rect 1244 232 1252 234
rect 1274 232 1282 234
rect 1304 232 1312 234
rect 664 224 1172 232
rect 1184 224 1202 232
rect 1214 224 1232 232
rect 1244 224 1262 232
rect 1274 224 1292 232
rect 1304 224 1322 232
rect 664 212 1162 224
rect 1184 222 1192 224
rect 1214 222 1222 224
rect 1244 222 1252 224
rect 1274 222 1282 224
rect 1304 222 1312 224
rect 1174 214 1192 222
rect 1204 214 1222 222
rect 1234 214 1252 222
rect 1264 214 1282 222
rect 1294 214 1312 222
rect 1184 212 1192 214
rect 1214 212 1222 214
rect 1244 212 1252 214
rect 1274 212 1282 214
rect 664 204 1172 212
rect 1184 204 1202 212
rect 1214 204 1232 212
rect 1244 204 1262 212
rect 1274 204 1292 212
rect 664 192 1162 204
rect 1184 202 1192 204
rect 1214 202 1222 204
rect 1244 202 1252 204
rect 1274 202 1282 204
rect 1304 202 1312 214
rect 1174 194 1192 202
rect 1204 194 1222 202
rect 1234 194 1252 202
rect 1264 194 1282 202
rect 1294 194 1312 202
rect 1184 192 1192 194
rect 1214 192 1222 194
rect 1244 192 1252 194
rect 1274 192 1282 194
rect 664 184 1172 192
rect 1184 184 1202 192
rect 1214 184 1232 192
rect 1244 184 1262 192
rect 1274 184 1292 192
rect 664 172 1162 184
rect 1184 182 1192 184
rect 1214 182 1222 184
rect 1244 182 1252 184
rect 1274 182 1282 184
rect 1304 182 1312 194
rect 1174 174 1192 182
rect 1204 174 1222 182
rect 1234 174 1252 182
rect 1264 174 1282 182
rect 1294 174 1312 182
rect 1184 172 1192 174
rect 1214 172 1222 174
rect 1244 172 1252 174
rect 1274 172 1282 174
rect 664 164 1172 172
rect 1184 164 1202 172
rect 1214 164 1232 172
rect 1244 164 1262 172
rect 1274 164 1292 172
rect 664 152 1162 164
rect 1184 162 1192 164
rect 1214 162 1222 164
rect 1244 162 1252 164
rect 1274 162 1282 164
rect 1304 162 1312 174
rect 1174 154 1192 162
rect 1204 154 1222 162
rect 1234 154 1252 162
rect 1264 154 1282 162
rect 1294 154 1312 162
rect 1184 152 1192 154
rect 1214 152 1222 154
rect 1244 152 1252 154
rect 1274 152 1282 154
rect 664 144 1172 152
rect 1184 144 1202 152
rect 1214 144 1232 152
rect 1244 144 1262 152
rect 1274 144 1292 152
rect 664 132 1162 144
rect 1184 142 1192 144
rect 1214 142 1222 144
rect 1244 142 1252 144
rect 1274 142 1282 144
rect 1304 142 1312 154
rect 1174 134 1192 142
rect 1204 134 1222 142
rect 1234 134 1252 142
rect 1264 134 1282 142
rect 1294 134 1312 142
rect 1184 132 1192 134
rect 1214 132 1222 134
rect 1244 132 1252 134
rect 1274 132 1282 134
rect 664 124 1172 132
rect 1184 124 1202 132
rect 1214 124 1232 132
rect 1244 124 1262 132
rect 1274 124 1292 132
rect 664 112 1162 124
rect 1184 122 1192 124
rect 1214 122 1222 124
rect 1244 122 1252 124
rect 1274 122 1282 124
rect 1304 122 1312 134
rect 1174 114 1192 122
rect 1204 114 1222 122
rect 1234 114 1252 122
rect 1264 114 1282 122
rect 1294 114 1312 122
rect 1184 112 1192 114
rect 1214 112 1222 114
rect 1244 112 1252 114
rect 1274 112 1282 114
rect 664 104 1172 112
rect 1184 104 1202 112
rect 1214 104 1232 112
rect 1244 104 1262 112
rect 1274 104 1292 112
rect 664 92 1162 104
rect 1184 102 1192 104
rect 1214 102 1222 104
rect 1244 102 1252 104
rect 1274 102 1282 104
rect 1304 102 1312 114
rect 1174 94 1192 102
rect 1204 94 1222 102
rect 1234 94 1252 102
rect 1264 94 1282 102
rect 1294 94 1312 102
rect 1184 92 1192 94
rect 1214 92 1222 94
rect 1244 92 1252 94
rect 1274 92 1282 94
rect 664 84 1172 92
rect 1184 84 1202 92
rect 1214 84 1232 92
rect 1244 84 1262 92
rect 1274 84 1292 92
rect 664 72 1162 84
rect 1184 82 1192 84
rect 1214 82 1222 84
rect 1244 82 1252 84
rect 1274 82 1282 84
rect 1304 82 1312 94
rect 1174 74 1192 82
rect 1204 74 1222 82
rect 1234 74 1252 82
rect 1264 74 1282 82
rect 1294 74 1312 82
rect 1184 72 1192 74
rect 1214 72 1222 74
rect 1244 72 1252 74
rect 1274 72 1282 74
rect 664 64 1172 72
rect 1184 64 1202 72
rect 1214 64 1232 72
rect 1244 64 1262 72
rect 1274 64 1292 72
rect 664 52 1162 64
rect 1184 62 1192 64
rect 1214 62 1222 64
rect 1244 62 1252 64
rect 1274 62 1282 64
rect 1304 62 1312 74
rect 1174 54 1192 62
rect 1204 54 1222 62
rect 1234 54 1252 62
rect 1264 54 1282 62
rect 1294 54 1312 62
rect 1184 52 1192 54
rect 1214 52 1222 54
rect 1244 52 1252 54
rect 1274 52 1282 54
rect 664 44 1172 52
rect 1184 44 1202 52
rect 1214 44 1232 52
rect 1244 44 1262 52
rect 1274 44 1292 52
rect 664 32 1162 44
rect 1184 42 1192 44
rect 1214 42 1222 44
rect 1244 42 1252 44
rect 1274 42 1282 44
rect 1304 42 1312 54
rect 1174 34 1192 42
rect 1204 34 1222 42
rect 1234 34 1252 42
rect 1264 34 1282 42
rect 1294 34 1312 42
rect 1184 32 1192 34
rect 1214 32 1222 34
rect 1244 32 1252 34
rect 1274 32 1282 34
rect 664 24 1172 32
rect 1184 24 1202 32
rect 1214 24 1232 32
rect 1244 24 1262 32
rect 1274 24 1292 32
rect 664 12 1162 24
rect 1184 22 1192 24
rect 1214 22 1222 24
rect 1244 22 1252 24
rect 1274 22 1282 24
rect 1304 22 1312 34
rect 1174 14 1192 22
rect 1204 14 1222 22
rect 1234 14 1252 22
rect 1264 14 1282 22
rect 1294 14 1312 22
rect 1184 12 1192 14
rect 1214 12 1222 14
rect 1244 12 1252 14
rect 1274 12 1282 14
rect 664 4 1172 12
rect 1184 4 1202 12
rect 1214 4 1232 12
rect 1244 4 1262 12
rect 1274 4 1292 12
rect 1304 4 1312 14
<< nsubstratencontact >>
rect 1820 632 1828 642
rect 1840 634 1858 642
rect 1870 634 1888 642
rect 1900 634 1918 642
rect 1930 634 1948 642
rect 1960 634 1978 642
rect 1990 634 1998 642
rect 1850 632 1858 634
rect 1880 632 1888 634
rect 1910 632 1918 634
rect 1940 632 1948 634
rect 1970 632 1978 634
rect 1810 624 1838 632
rect 1850 624 1868 632
rect 1880 624 1898 632
rect 1910 624 1928 632
rect 1940 624 1958 632
rect 1970 624 1988 632
rect 1810 622 1828 624
rect 1850 622 1858 624
rect 1880 622 1888 624
rect 1910 622 1918 624
rect 1940 622 1948 624
rect 1970 622 1978 624
rect 1800 614 1828 622
rect 1840 614 1858 622
rect 1870 614 1888 622
rect 1900 614 1918 622
rect 1930 614 1948 622
rect 1960 614 1978 622
rect 1990 614 1998 622
rect 1800 612 1808 614
rect 1790 604 1808 612
rect 1820 612 1828 614
rect 1850 612 1858 614
rect 1880 612 1888 614
rect 1910 612 1918 614
rect 1940 612 1948 614
rect 1970 612 1978 614
rect 1820 604 1838 612
rect 1850 604 1868 612
rect 1880 604 1898 612
rect 1910 604 1928 612
rect 1940 604 1958 612
rect 1970 604 1988 612
rect 1790 602 1798 604
rect 1820 602 1828 604
rect 1850 602 1858 604
rect 1880 602 1888 604
rect 1910 602 1918 604
rect 1940 602 1948 604
rect 1970 602 1978 604
rect 1780 594 1798 602
rect 1780 592 1788 594
rect 1810 592 1828 602
rect 1840 594 1858 602
rect 1870 594 1888 602
rect 1900 594 1918 602
rect 1930 594 1948 602
rect 1960 594 1978 602
rect 1990 594 1998 602
rect 1850 592 1858 594
rect 1880 592 1888 594
rect 1910 592 1918 594
rect 1940 592 1948 594
rect 1970 592 1978 594
rect 1770 584 1788 592
rect 1800 584 1838 592
rect 1770 582 1778 584
rect 1800 582 1808 584
rect 1760 574 1778 582
rect 1790 574 1808 582
rect 1760 572 1768 574
rect 1790 572 1798 574
rect 1820 572 1828 584
rect 1850 582 1868 592
rect 1880 584 1898 592
rect 1910 584 1928 592
rect 1940 584 1958 592
rect 1970 584 1988 592
rect 1880 582 1888 584
rect 1910 582 1918 584
rect 1940 582 1948 584
rect 1970 582 1978 584
rect 1840 574 1888 582
rect 1900 574 1918 582
rect 1930 574 1948 582
rect 1960 574 1978 582
rect 1990 574 1998 582
rect 1840 572 1868 574
rect 1750 564 1768 572
rect 1780 564 1798 572
rect 1810 564 1868 572
rect 1880 572 1888 574
rect 1910 572 1918 574
rect 1940 572 1948 574
rect 1970 572 1978 574
rect 1880 564 1898 572
rect 1910 564 1928 572
rect 1940 564 1958 572
rect 1970 564 1988 572
rect 1750 562 1758 564
rect 1780 562 1788 564
rect 1810 562 1858 564
rect 1880 562 1888 564
rect 1910 562 1918 564
rect 1940 562 1948 564
rect 1970 562 1978 564
rect 1740 554 1758 562
rect 1770 554 1788 562
rect 1800 554 1858 562
rect 1870 554 1888 562
rect 1900 554 1918 562
rect 1930 554 1948 562
rect 1960 554 1978 562
rect 1990 554 1998 562
rect 1740 552 1748 554
rect 1770 552 1778 554
rect 1800 552 1838 554
rect 1730 544 1748 552
rect 1760 544 1778 552
rect 1790 544 1838 552
rect 1850 552 1858 554
rect 1880 552 1888 554
rect 1910 552 1918 554
rect 1940 552 1948 554
rect 1970 552 1978 554
rect 1850 544 1868 552
rect 1880 544 1898 552
rect 1910 544 1928 552
rect 1940 544 1958 552
rect 1970 544 1988 552
rect 1730 542 1738 544
rect 1760 542 1768 544
rect 1790 542 1828 544
rect 1850 542 1858 544
rect 1880 542 1888 544
rect 1910 542 1918 544
rect 1940 542 1948 544
rect 1970 542 1978 544
rect 1720 534 1738 542
rect 1750 534 1768 542
rect 1780 534 1828 542
rect 1840 534 1858 542
rect 1870 534 1888 542
rect 1900 534 1918 542
rect 1930 534 1948 542
rect 1960 534 1978 542
rect 1990 534 1998 542
rect 1720 532 1728 534
rect 1750 532 1758 534
rect 1780 532 1808 534
rect 1710 524 1728 532
rect 1740 524 1758 532
rect 1770 531 1808 532
rect 1820 532 1828 534
rect 1850 532 1858 534
rect 1880 532 1888 534
rect 1910 532 1918 534
rect 1940 532 1948 534
rect 1970 532 1978 534
rect 1820 531 1838 532
rect 1770 524 1838 531
rect 1850 524 1868 532
rect 1880 524 1898 532
rect 1910 524 1928 532
rect 1940 524 1958 532
rect 1970 524 1988 532
rect 1710 522 1718 524
rect 1740 522 1748 524
rect 1770 523 1828 524
rect 1770 522 1808 523
rect 1700 514 1718 522
rect 1730 514 1748 522
rect 1760 514 1808 522
rect 1700 512 1708 514
rect 1730 512 1738 514
rect 1760 512 1798 514
rect 1820 512 1828 523
rect 1850 522 1858 524
rect 1880 522 1888 524
rect 1910 522 1918 524
rect 1940 522 1948 524
rect 1970 522 1978 524
rect 1840 514 1858 522
rect 1870 514 1888 522
rect 1900 514 1918 522
rect 1930 514 1948 522
rect 1960 514 1978 522
rect 1990 514 1998 522
rect 1850 512 1858 514
rect 1880 512 1888 514
rect 1910 512 1918 514
rect 1940 512 1948 514
rect 1970 512 1978 514
rect 1690 502 1708 512
rect 1720 502 1738 512
rect 1750 502 1798 512
rect 1810 502 1838 512
rect 1850 502 1868 512
rect 1880 502 1898 512
rect 1910 502 1928 512
rect 1940 502 1958 512
rect 1970 502 1988 512
rect 1680 494 1998 502
rect 1670 484 1678 492
rect 1690 484 1698 494
rect 1710 484 1718 494
rect 1730 484 1738 494
rect 1750 484 1788 494
rect 1800 484 1808 494
rect 1820 484 1828 494
rect 1840 484 1848 494
rect 1860 484 1868 494
rect 1750 482 1778 484
rect 1890 482 1998 494
rect 1660 474 1668 482
rect 1680 474 1688 482
rect 1700 474 1708 482
rect 1720 474 1728 482
rect 1740 474 1778 482
rect 1790 474 1798 482
rect 1810 474 1818 482
rect 1830 474 1838 482
rect 1850 474 1858 482
rect 1740 472 1768 474
rect 1880 472 1998 482
rect 1650 464 1658 472
rect 1670 464 1678 472
rect 1690 464 1698 472
rect 1710 464 1718 472
rect 1730 464 1768 472
rect 1780 464 1788 472
rect 1800 464 1808 472
rect 1820 464 1828 472
rect 1840 464 1848 472
rect 1730 462 1758 464
rect 1870 462 1998 472
rect 1640 454 1648 462
rect 1660 454 1668 462
rect 1680 454 1688 462
rect 1700 454 1708 462
rect 1720 454 1758 462
rect 1770 454 1778 462
rect 1790 454 1798 462
rect 1810 454 1818 462
rect 1830 454 1838 462
rect 1720 452 1748 454
rect 1860 452 1998 462
rect 1630 444 1638 452
rect 1650 444 1658 452
rect 1670 444 1678 452
rect 1690 444 1698 452
rect 1710 444 1748 452
rect 1760 444 1768 452
rect 1780 444 1788 452
rect 1800 444 1808 452
rect 1820 444 1828 452
rect 1710 442 1738 444
rect 1850 442 1998 452
rect 1620 434 1628 442
rect 1640 434 1648 442
rect 1660 434 1668 442
rect 1680 434 1688 442
rect 1700 434 1738 442
rect 1750 434 1758 442
rect 1770 434 1778 442
rect 1790 434 1798 442
rect 1810 434 1818 442
rect 1700 432 1728 434
rect 1840 432 1998 442
rect 1610 424 1618 432
rect 1630 424 1638 432
rect 1650 424 1658 432
rect 1670 424 1678 432
rect 1690 424 1728 432
rect 1740 424 1748 432
rect 1760 424 1768 432
rect 1780 424 1788 432
rect 1800 424 1808 432
rect 1690 422 1718 424
rect 1600 414 1608 422
rect 1620 414 1628 422
rect 1640 414 1648 422
rect 1660 414 1668 422
rect 1680 414 1718 422
rect 1730 414 1738 422
rect 1750 414 1758 422
rect 1770 414 1778 422
rect 1790 414 1798 422
rect 1830 414 1998 432
rect 1680 412 1708 414
rect 1590 404 1598 412
rect 1610 404 1618 412
rect 1630 404 1638 412
rect 1650 404 1658 412
rect 1670 404 1708 412
rect 1720 404 1728 412
rect 1740 404 1748 412
rect 1760 404 1768 412
rect 1780 404 1788 412
rect 1670 402 1698 404
rect 1840 402 1998 414
rect 1580 394 1588 402
rect 1600 394 1608 402
rect 1620 394 1628 402
rect 1640 394 1648 402
rect 1660 394 1698 402
rect 1710 394 1718 402
rect 1730 394 1738 402
rect 1750 394 1758 402
rect 1770 394 1778 402
rect 1660 392 1688 394
rect 1830 392 1998 402
rect 1570 384 1578 392
rect 1590 384 1598 392
rect 1610 384 1618 392
rect 1630 384 1638 392
rect 1650 384 1688 392
rect 1700 384 1708 392
rect 1720 384 1728 392
rect 1740 384 1748 392
rect 1760 384 1768 392
rect 1650 382 1678 384
rect 1820 382 1998 392
rect 1560 374 1568 382
rect 1580 374 1588 382
rect 1600 374 1608 382
rect 1620 374 1628 382
rect 1640 374 1678 382
rect 1690 374 1698 382
rect 1710 374 1718 382
rect 1730 374 1738 382
rect 1750 374 1758 382
rect 1640 372 1668 374
rect 1810 372 1998 382
rect 1550 364 1558 372
rect 1570 364 1578 372
rect 1590 364 1598 372
rect 1610 364 1618 372
rect 1630 364 1668 372
rect 1680 364 1688 372
rect 1700 364 1708 372
rect 1720 364 1728 372
rect 1740 364 1748 372
rect 1630 362 1658 364
rect 1800 362 1998 372
rect 1540 354 1548 362
rect 1560 354 1568 362
rect 1580 354 1588 362
rect 1600 354 1608 362
rect 1620 354 1658 362
rect 1670 354 1678 362
rect 1690 354 1698 362
rect 1710 354 1718 362
rect 1730 354 1738 362
rect 1620 352 1648 354
rect 1790 352 1998 362
rect 1530 344 1538 352
rect 1550 344 1558 352
rect 1570 344 1578 352
rect 1590 344 1598 352
rect 1610 344 1648 352
rect 1660 344 1668 352
rect 1680 344 1688 352
rect 1700 344 1708 352
rect 1720 344 1728 352
rect 1610 342 1638 344
rect 1780 342 1998 352
rect 1520 334 1528 342
rect 1540 334 1548 342
rect 1560 334 1568 342
rect 1580 334 1588 342
rect 1600 334 1638 342
rect 1650 334 1658 342
rect 1670 334 1678 342
rect 1690 334 1698 342
rect 1710 334 1718 342
rect 1600 332 1628 334
rect 1770 332 1998 342
rect 1510 324 1518 332
rect 1530 324 1538 332
rect 1550 324 1558 332
rect 1570 324 1578 332
rect 1590 324 1628 332
rect 1640 324 1648 332
rect 1660 324 1668 332
rect 1680 324 1688 332
rect 1700 324 1708 332
rect 1590 322 1618 324
rect 1760 322 1998 332
rect 1500 314 1508 322
rect 1520 314 1528 322
rect 1540 314 1548 322
rect 1560 314 1568 322
rect 1580 314 1618 322
rect 1630 314 1638 322
rect 1650 314 1658 322
rect 1670 314 1678 322
rect 1690 314 1698 322
rect 1580 312 1608 314
rect 1750 312 1998 322
rect 1490 304 1498 312
rect 1510 304 1518 312
rect 1530 304 1538 312
rect 1550 304 1558 312
rect 1570 304 1608 312
rect 1620 304 1628 312
rect 1640 304 1648 312
rect 1660 304 1668 312
rect 1680 304 1688 312
rect 1570 302 1598 304
rect 1740 302 1998 312
rect 1480 294 1488 302
rect 1500 294 1508 302
rect 1520 294 1528 302
rect 1540 294 1548 302
rect 1560 294 1598 302
rect 1610 294 1618 302
rect 1630 294 1638 302
rect 1650 294 1658 302
rect 1670 294 1678 302
rect 1560 292 1588 294
rect 1730 292 1998 302
rect 1470 284 1478 292
rect 1490 284 1498 292
rect 1510 284 1518 292
rect 1530 284 1538 292
rect 1550 284 1588 292
rect 1600 284 1608 292
rect 1620 284 1628 292
rect 1640 284 1648 292
rect 1660 284 1668 292
rect 1550 282 1578 284
rect 1720 282 1998 292
rect 1460 274 1468 282
rect 1480 274 1488 282
rect 1500 274 1508 282
rect 1520 274 1528 282
rect 1540 274 1578 282
rect 1590 274 1598 282
rect 1610 274 1618 282
rect 1630 274 1638 282
rect 1650 274 1658 282
rect 1540 272 1568 274
rect 1710 272 1998 282
rect 1450 264 1458 272
rect 1470 264 1478 272
rect 1490 264 1498 272
rect 1510 264 1518 272
rect 1530 264 1568 272
rect 1580 264 1588 272
rect 1600 264 1608 272
rect 1620 264 1628 272
rect 1640 264 1648 272
rect 1530 262 1558 264
rect 1700 262 1998 272
rect 1440 254 1448 262
rect 1460 254 1468 262
rect 1480 254 1488 262
rect 1500 254 1508 262
rect 1520 254 1558 262
rect 1570 254 1578 262
rect 1590 254 1598 262
rect 1610 254 1618 262
rect 1630 254 1638 262
rect 1520 252 1548 254
rect 1690 252 1998 262
rect 1430 244 1438 252
rect 1450 244 1458 252
rect 1470 244 1478 252
rect 1490 244 1498 252
rect 1510 244 1548 252
rect 1560 244 1568 252
rect 1580 244 1588 252
rect 1600 244 1608 252
rect 1620 244 1628 252
rect 1510 242 1538 244
rect 1680 242 1998 252
rect 1420 234 1428 242
rect 1440 234 1448 242
rect 1460 234 1468 242
rect 1480 234 1488 242
rect 1500 234 1538 242
rect 1550 234 1558 242
rect 1570 234 1578 242
rect 1590 234 1598 242
rect 1610 234 1618 242
rect 1500 232 1528 234
rect 1670 232 1998 242
rect 1410 224 1418 232
rect 1430 224 1438 232
rect 1450 224 1458 232
rect 1470 224 1478 232
rect 1490 224 1528 232
rect 1540 224 1548 232
rect 1560 224 1568 232
rect 1580 224 1588 232
rect 1600 224 1608 232
rect 1490 222 1518 224
rect 1660 222 1998 232
rect 1400 214 1408 222
rect 1420 214 1428 222
rect 1440 214 1448 222
rect 1460 214 1468 222
rect 1480 214 1518 222
rect 1530 214 1538 222
rect 1550 214 1558 222
rect 1570 214 1578 222
rect 1590 214 1598 222
rect 1480 212 1508 214
rect 1650 212 1998 222
rect 1390 204 1398 212
rect 1410 204 1418 212
rect 1430 204 1438 212
rect 1450 204 1458 212
rect 1470 204 1508 212
rect 1520 204 1528 212
rect 1540 204 1548 212
rect 1560 204 1568 212
rect 1580 204 1588 212
rect 1470 202 1498 204
rect 1640 202 1998 212
rect 1380 194 1388 202
rect 1400 194 1408 202
rect 1420 194 1428 202
rect 1440 194 1448 202
rect 1460 194 1498 202
rect 1510 194 1518 202
rect 1530 194 1538 202
rect 1550 194 1558 202
rect 1570 194 1578 202
rect 1460 192 1488 194
rect 1630 192 1998 202
rect 1370 182 1378 192
rect 1390 182 1398 192
rect 1410 182 1418 192
rect 1430 182 1438 192
rect 1450 182 1488 192
rect 1500 182 1508 192
rect 1520 182 1528 192
rect 1540 182 1548 192
rect 1560 182 1568 192
rect 1620 182 1998 192
rect 1360 174 1568 182
rect 1350 142 1358 172
rect 1370 144 1378 174
rect 1390 142 1398 174
rect 1350 134 1368 142
rect 1380 134 1398 142
rect 1410 142 1418 174
rect 1430 144 1468 174
rect 1410 134 1428 142
rect 1440 134 1458 144
rect 1480 142 1488 174
rect 1470 134 1488 142
rect 1500 142 1508 174
rect 1520 142 1528 174
rect 1540 142 1548 174
rect 1610 172 1998 182
rect 1600 162 1998 172
rect 1590 152 1998 162
rect 1580 142 1998 152
rect 1350 122 1358 134
rect 1380 132 1388 134
rect 1410 132 1418 134
rect 1440 132 1448 134
rect 1470 132 1478 134
rect 1500 132 1998 142
rect 1370 124 1388 132
rect 1400 124 1418 132
rect 1430 124 1448 132
rect 1460 124 1478 132
rect 1490 124 1998 132
rect 1380 122 1388 124
rect 1410 122 1418 124
rect 1440 122 1448 124
rect 1470 122 1478 124
rect 1350 114 1368 122
rect 1380 114 1398 122
rect 1410 114 1428 122
rect 1440 114 1458 122
rect 1470 114 1488 122
rect 1350 102 1358 114
rect 1380 112 1388 114
rect 1410 112 1418 114
rect 1440 112 1448 114
rect 1470 112 1478 114
rect 1500 112 1998 124
rect 1370 104 1388 112
rect 1400 104 1418 112
rect 1430 104 1448 112
rect 1460 104 1478 112
rect 1490 104 1998 112
rect 1380 102 1388 104
rect 1410 102 1418 104
rect 1440 102 1448 104
rect 1470 102 1478 104
rect 1350 94 1368 102
rect 1380 94 1398 102
rect 1410 94 1428 102
rect 1440 94 1458 102
rect 1470 94 1488 102
rect 1350 82 1358 94
rect 1380 92 1388 94
rect 1410 92 1418 94
rect 1440 92 1448 94
rect 1470 92 1478 94
rect 1500 92 1998 104
rect 1370 84 1388 92
rect 1400 84 1418 92
rect 1430 84 1448 92
rect 1460 84 1478 92
rect 1490 84 1998 92
rect 1380 82 1388 84
rect 1410 82 1418 84
rect 1440 82 1448 84
rect 1470 82 1478 84
rect 1350 74 1368 82
rect 1380 74 1398 82
rect 1410 74 1428 82
rect 1440 74 1458 82
rect 1470 74 1488 82
rect 1350 62 1358 74
rect 1380 72 1388 74
rect 1410 72 1418 74
rect 1440 72 1448 74
rect 1470 72 1478 74
rect 1500 72 1998 84
rect 1370 64 1388 72
rect 1400 64 1418 72
rect 1430 64 1448 72
rect 1460 64 1478 72
rect 1490 64 1998 72
rect 1380 62 1388 64
rect 1410 62 1418 64
rect 1440 62 1448 64
rect 1470 62 1478 64
rect 1350 54 1368 62
rect 1380 54 1398 62
rect 1410 54 1428 62
rect 1440 54 1458 62
rect 1470 54 1488 62
rect 1350 42 1358 54
rect 1380 52 1388 54
rect 1410 52 1418 54
rect 1440 52 1448 54
rect 1470 52 1478 54
rect 1500 52 1998 64
rect 1370 44 1388 52
rect 1400 44 1418 52
rect 1430 44 1448 52
rect 1460 44 1478 52
rect 1490 44 1998 52
rect 1380 42 1388 44
rect 1410 42 1418 44
rect 1440 42 1448 44
rect 1470 42 1478 44
rect 1350 34 1368 42
rect 1380 34 1398 42
rect 1410 34 1428 42
rect 1440 34 1458 42
rect 1470 34 1488 42
rect 1350 22 1358 34
rect 1380 32 1388 34
rect 1410 32 1418 34
rect 1440 32 1448 34
rect 1470 32 1478 34
rect 1500 32 1998 44
rect 1370 24 1388 32
rect 1400 24 1418 32
rect 1430 24 1448 32
rect 1460 24 1478 32
rect 1490 24 1998 32
rect 1380 22 1388 24
rect 1410 22 1418 24
rect 1440 22 1448 24
rect 1470 22 1478 24
rect 1350 14 1368 22
rect 1380 14 1398 22
rect 1410 14 1428 22
rect 1440 14 1458 22
rect 1470 14 1488 22
rect 1350 4 1358 14
rect 1380 12 1388 14
rect 1410 12 1418 14
rect 1440 12 1448 14
rect 1470 12 1478 14
rect 1500 12 1998 24
rect 1370 4 1388 12
rect 1400 4 1418 12
rect 1430 4 1448 12
rect 1460 4 1478 12
rect 1490 4 1998 12
<< metal1 >>
tri 1574 1332 1582 1340 se
rect 1582 1338 1722 1340
rect 1582 1332 2000 1338
tri 1566 1324 1574 1332 se
rect 1574 1324 1584 1332
tri 1564 1322 1566 1324 se
rect 1566 1322 1584 1324
tri 1556 1314 1564 1322 se
rect 1564 1314 1574 1322
tri 1554 1312 1556 1314 se
rect 1556 1312 1574 1314
tri 1546 1304 1554 1312 se
rect 1554 1304 1564 1312
tri 1544 1302 1546 1304 se
rect 1546 1302 1564 1304
tri 1536 1294 1544 1302 se
rect 1544 1294 1554 1302
tri 1534 1292 1536 1294 se
rect 1536 1292 1554 1294
tri 1526 1284 1534 1292 se
rect 1534 1284 1544 1292
tri 1524 1282 1526 1284 se
rect 1526 1282 1544 1284
tri 1516 1274 1524 1282 se
rect 1524 1274 1534 1282
tri 1514 1272 1516 1274 se
rect 1516 1272 1534 1274
tri 1506 1264 1514 1272 se
rect 1514 1264 1524 1272
tri 1504 1262 1506 1264 se
rect 1506 1262 1524 1264
tri 1496 1254 1504 1262 se
rect 1504 1254 1514 1262
tri 1494 1252 1496 1254 se
rect 1496 1252 1514 1254
tri 1486 1244 1494 1252 se
rect 1494 1244 1504 1252
tri 1484 1242 1486 1244 se
rect 1486 1242 1504 1244
tri 1476 1234 1484 1242 se
rect 1484 1234 1494 1242
tri 1474 1232 1476 1234 se
rect 1476 1232 1494 1234
tri 1466 1224 1474 1232 se
rect 1474 1224 1484 1232
tri 1464 1222 1466 1224 se
rect 1466 1222 1484 1224
tri 1456 1214 1464 1222 se
rect 1464 1214 1474 1222
tri 1454 1212 1456 1214 se
rect 1456 1212 1474 1214
tri 1446 1204 1454 1212 se
rect 1454 1204 1464 1212
tri 1444 1202 1446 1204 se
rect 1446 1202 1464 1204
tri 1436 1194 1444 1202 se
rect 1444 1194 1454 1202
tri 1434 1192 1436 1194 se
rect 1436 1192 1454 1194
tri 1426 1184 1434 1192 se
rect 1434 1184 1444 1192
tri 1424 1182 1426 1184 se
rect 1426 1182 1444 1184
tri 1416 1174 1424 1182 se
rect 1424 1174 1434 1182
tri 1414 1172 1416 1174 se
rect 1416 1172 1434 1174
tri 1406 1164 1414 1172 se
rect 1414 1164 1424 1172
tri 1404 1162 1406 1164 se
rect 1406 1162 1424 1164
tri 1396 1154 1404 1162 se
rect 1404 1154 1414 1162
tri 1394 1152 1396 1154 se
rect 1396 1152 1414 1154
tri 1386 1144 1394 1152 se
rect 1394 1144 1404 1152
tri 1384 1142 1386 1144 se
rect 1386 1142 1404 1144
tri 1376 1134 1384 1142 se
rect 1384 1134 1394 1142
tri 1374 1132 1376 1134 se
rect 1376 1132 1394 1134
tri 1366 1124 1374 1132 se
rect 1374 1124 1384 1132
tri 1364 1122 1366 1124 se
rect 1366 1122 1384 1124
tri 1356 1114 1364 1122 se
rect 1364 1114 1374 1122
tri 1354 1112 1356 1114 se
rect 1356 1112 1374 1114
tri 1346 1104 1354 1112 se
rect 1354 1104 1364 1112
tri 1344 1102 1346 1104 se
rect 1346 1102 1364 1104
tri 1336 1094 1344 1102 se
rect 1344 1094 1354 1102
tri 1334 1092 1336 1094 se
rect 1336 1092 1354 1094
tri 1326 1084 1334 1092 se
rect 1334 1084 1344 1092
tri 1324 1082 1326 1084 se
rect 1326 1082 1344 1084
tri 1316 1074 1324 1082 se
rect 1324 1074 1334 1082
tri 1314 1072 1316 1074 se
rect 1316 1072 1334 1074
tri 1306 1064 1314 1072 se
rect 1314 1064 1324 1072
tri 1304 1062 1306 1064 se
rect 1306 1062 1324 1064
tri 1296 1054 1304 1062 se
rect 1304 1054 1314 1062
tri 1294 1052 1296 1054 se
rect 1296 1052 1314 1054
tri 1286 1044 1294 1052 se
rect 1294 1044 1304 1052
rect 1572 1047 1594 1054
rect 1572 1044 1580 1047
tri 1580 1044 1583 1047 nw
tri 1583 1044 1586 1047 ne
rect 1586 1044 1594 1047
tri 1284 1042 1286 1044 se
rect 1286 1042 1304 1044
rect 1562 1042 1578 1044
tri 1578 1042 1580 1044 nw
tri 1586 1042 1588 1044 ne
rect 1588 1042 1594 1044
tri 1276 1034 1284 1042 se
rect 1284 1034 1294 1042
rect 1562 1039 1575 1042
tri 1575 1039 1578 1042 nw
tri 1588 1039 1591 1042 ne
rect 1562 1034 1570 1039
tri 1570 1034 1575 1039 nw
tri 1586 1034 1591 1039 se
rect 1591 1034 1594 1042
tri 1274 1032 1276 1034 se
rect 1276 1032 1294 1034
rect 1552 1032 1568 1034
tri 1568 1032 1570 1034 nw
tri 1584 1032 1586 1034 se
rect 1586 1032 1594 1034
tri 1266 1024 1274 1032 se
rect 1274 1024 1284 1032
rect 1552 1024 1560 1032
tri 1560 1024 1568 1032 nw
tri 1576 1024 1584 1032 se
rect 1584 1024 1594 1032
tri 1264 1022 1266 1024 se
rect 1266 1022 1284 1024
rect 1542 1022 1558 1024
tri 1558 1022 1560 1024 nw
tri 1574 1022 1576 1024 se
rect 1576 1022 1594 1024
tri 1256 1014 1264 1022 se
rect 1264 1014 1274 1022
rect 1542 1014 1550 1022
tri 1550 1014 1558 1022 nw
tri 1566 1014 1574 1022 se
rect 1574 1014 1584 1022
tri 1254 1012 1256 1014 se
rect 1256 1012 1274 1014
rect 1532 1012 1548 1014
tri 1548 1012 1550 1014 nw
tri 1564 1012 1566 1014 se
rect 1566 1012 1584 1014
tri 1250 1008 1254 1012 se
rect 1254 1008 1264 1012
tri 1246 1004 1250 1008 se
rect 1250 1004 1264 1008
rect 1532 1008 1544 1012
tri 1544 1008 1548 1012 nw
tri 1560 1008 1564 1012 se
rect 1564 1008 1574 1012
rect 1532 1004 1540 1008
tri 1540 1004 1544 1008 nw
tri 1556 1004 1560 1008 se
rect 1560 1004 1574 1008
tri 1244 1002 1246 1004 se
rect 1246 1002 1264 1004
rect 1522 1002 1538 1004
tri 1538 1002 1540 1004 nw
tri 1554 1002 1556 1004 se
rect 1556 1002 1574 1004
tri 1236 994 1244 1002 se
rect 1244 994 1254 1002
rect 1522 994 1530 1002
tri 1530 994 1538 1002 nw
tri 1546 994 1554 1002 se
rect 1554 994 1564 1002
tri 1234 992 1236 994 se
rect 1236 992 1254 994
rect 1512 992 1528 994
tri 1528 992 1530 994 nw
tri 1544 992 1546 994 se
rect 1546 992 1564 994
tri 1226 984 1234 992 se
rect 1234 984 1244 992
rect 1512 984 1520 992
tri 1520 984 1528 992 nw
tri 1536 984 1544 992 se
rect 1544 984 1554 992
tri 1224 982 1226 984 se
rect 1226 982 1244 984
rect 1502 982 1518 984
tri 1518 982 1520 984 nw
tri 1534 982 1536 984 se
rect 1536 982 1554 984
tri 1216 974 1224 982 se
rect 1224 974 1234 982
rect 1502 974 1510 982
tri 1510 974 1518 982 nw
tri 1526 974 1534 982 se
rect 1534 974 1544 982
tri 1214 972 1216 974 se
rect 1216 972 1234 974
rect 1492 972 1508 974
tri 1508 972 1510 974 nw
tri 1524 972 1526 974 se
rect 1526 972 1544 974
tri 1206 964 1214 972 se
rect 1214 964 1224 972
rect 1492 964 1500 972
tri 1500 964 1508 972 nw
tri 1516 964 1524 972 se
rect 1524 964 1534 972
tri 1204 962 1206 964 se
rect 1206 962 1224 964
rect 1482 962 1498 964
tri 1498 962 1500 964 nw
tri 1514 962 1516 964 se
rect 1516 962 1534 964
tri 1196 954 1204 962 se
rect 1204 954 1214 962
rect 1482 954 1490 962
tri 1490 954 1498 962 nw
tri 1506 954 1514 962 se
rect 1514 954 1524 962
tri 1194 952 1196 954 se
rect 1196 952 1214 954
rect 1472 952 1488 954
tri 1488 952 1490 954 nw
tri 1504 952 1506 954 se
rect 1506 952 1524 954
tri 1186 944 1194 952 se
rect 1194 944 1204 952
rect 1472 944 1480 952
tri 1480 944 1488 952 nw
tri 1496 944 1504 952 se
rect 1504 944 1514 952
tri 1184 942 1186 944 se
rect 1186 942 1204 944
rect 1462 942 1478 944
tri 1478 942 1480 944 nw
tri 1494 942 1496 944 se
rect 1496 942 1514 944
tri 1176 934 1184 942 se
rect 1184 934 1194 942
rect 1462 934 1470 942
tri 1470 934 1478 942 nw
tri 1486 934 1494 942 se
rect 1494 934 1504 942
tri 1174 932 1176 934 se
rect 1176 932 1194 934
rect 1452 932 1468 934
tri 1468 932 1470 934 nw
tri 1484 932 1486 934 se
rect 1486 932 1504 934
tri 1166 924 1174 932 se
rect 1174 924 1184 932
rect 1452 924 1460 932
tri 1460 924 1468 932 nw
tri 1476 924 1484 932 se
rect 1484 924 1494 932
tri 1164 922 1166 924 se
rect 1166 922 1184 924
rect 1442 922 1458 924
tri 1458 922 1460 924 nw
tri 1474 922 1476 924 se
rect 1476 922 1494 924
tri 1156 914 1164 922 se
rect 1164 914 1174 922
rect 1442 914 1450 922
tri 1450 914 1458 922 nw
tri 1466 914 1474 922 se
rect 1474 914 1484 922
tri 1154 912 1156 914 se
rect 1156 912 1174 914
rect 1432 912 1448 914
tri 1448 912 1450 914 nw
tri 1464 912 1466 914 se
rect 1466 912 1484 914
tri 1146 904 1154 912 se
rect 1154 904 1164 912
rect 1432 904 1440 912
tri 1440 904 1448 912 nw
tri 1456 904 1464 912 se
rect 1464 904 1474 912
tri 1144 902 1146 904 se
rect 1146 902 1164 904
rect 1422 902 1438 904
tri 1438 902 1440 904 nw
tri 1454 902 1456 904 se
rect 1456 902 1474 904
tri 1136 894 1144 902 se
rect 1144 894 1154 902
rect 1422 894 1430 902
tri 1430 894 1438 902 nw
tri 1446 894 1454 902 se
rect 1454 894 1464 902
tri 1134 892 1136 894 se
rect 1136 892 1154 894
rect 1412 892 1428 894
tri 1428 892 1430 894 nw
tri 1444 892 1446 894 se
rect 1446 892 1464 894
tri 1126 884 1134 892 se
rect 1134 884 1144 892
rect 1412 884 1420 892
tri 1420 884 1428 892 nw
tri 1436 884 1444 892 se
rect 1444 884 1454 892
tri 1124 882 1126 884 se
rect 1126 882 1144 884
rect 1402 882 1418 884
tri 1418 882 1420 884 nw
tri 1434 882 1436 884 se
rect 1436 882 1454 884
rect 1702 882 1720 884
tri 1720 882 1722 884 nw
tri 1722 882 1724 884 ne
rect 1724 882 1734 884
tri 1116 874 1124 882 se
rect 1124 874 1134 882
rect 1402 874 1410 882
tri 1410 874 1418 882 nw
tri 1426 874 1434 882 se
rect 1434 874 1444 882
rect 1702 876 1714 882
tri 1714 876 1720 882 nw
tri 1724 876 1730 882 ne
rect 1702 874 1712 876
tri 1712 874 1714 876 nw
tri 1728 874 1730 876 se
rect 1730 874 1734 882
tri 1114 872 1116 874 se
rect 1116 872 1134 874
rect 1392 872 1408 874
tri 1408 872 1410 874 nw
tri 1424 872 1426 874 se
rect 1426 872 1444 874
rect 1692 872 1710 874
tri 1710 872 1712 874 nw
tri 1726 872 1728 874 se
rect 1728 872 1734 874
tri 1106 864 1114 872 se
rect 1114 864 1124 872
rect 1392 864 1400 872
tri 1400 864 1408 872 nw
tri 1416 864 1424 872 se
rect 1424 864 1434 872
rect 1692 864 1702 872
tri 1702 864 1710 872 nw
tri 1718 864 1726 872 se
rect 1726 864 1734 872
tri 1104 862 1106 864 se
rect 1106 862 1124 864
rect 1382 862 1398 864
tri 1398 862 1400 864 nw
tri 1414 862 1416 864 se
rect 1416 862 1434 864
rect 1682 862 1700 864
tri 1700 862 1702 864 nw
tri 1716 862 1718 864 se
rect 1718 862 1734 864
tri 1096 854 1104 862 se
rect 1104 854 1114 862
rect 1382 854 1390 862
tri 1390 854 1398 862 nw
tri 1406 854 1414 862 se
rect 1414 854 1424 862
rect 1682 854 1692 862
tri 1692 854 1700 862 nw
tri 1708 854 1716 862 se
rect 1716 854 1724 862
tri 1094 852 1096 854 se
rect 1096 852 1114 854
rect 1372 852 1388 854
tri 1388 852 1390 854 nw
tri 1404 852 1406 854 se
rect 1406 852 1424 854
rect 1672 852 1690 854
tri 1690 852 1692 854 nw
tri 1706 852 1708 854 se
rect 1708 852 1724 854
tri 1086 844 1094 852 se
rect 1094 844 1104 852
rect 1372 844 1380 852
tri 1380 844 1388 852 nw
tri 1396 844 1404 852 se
rect 1404 844 1414 852
rect 1672 844 1682 852
tri 1682 844 1690 852 nw
tri 1698 844 1706 852 se
rect 1706 844 1714 852
tri 1084 842 1086 844 se
rect 1086 842 1104 844
rect 1362 842 1378 844
tri 1378 842 1380 844 nw
tri 1394 842 1396 844 se
rect 1396 842 1414 844
rect 1662 842 1680 844
tri 1680 842 1682 844 nw
tri 1696 842 1698 844 se
rect 1698 842 1714 844
rect 1722 842 1734 844
tri 1076 834 1084 842 se
rect 1084 834 1094 842
rect 1362 834 1370 842
tri 1370 834 1378 842 nw
tri 1386 834 1394 842 se
rect 1394 834 1404 842
rect 1662 834 1672 842
tri 1672 834 1680 842 nw
tri 1688 834 1696 842 se
rect 1696 834 1704 842
tri 1074 832 1076 834 se
rect 1076 832 1094 834
rect 1352 832 1368 834
tri 1368 832 1370 834 nw
tri 1384 832 1386 834 se
rect 1386 832 1404 834
rect 1652 832 1670 834
tri 1670 832 1672 834 nw
tri 1686 832 1688 834 se
rect 1688 832 1704 834
rect 1722 834 1724 842
rect 1732 834 1734 842
rect 1752 842 1764 844
rect 1752 834 1754 842
rect 1762 834 1764 842
rect 1782 842 1794 844
rect 1782 834 1784 842
rect 1792 834 1794 842
rect 1812 842 1824 844
rect 1812 834 1814 842
rect 1822 834 1824 842
rect 1842 842 1854 844
rect 1842 834 1844 842
rect 1852 834 1854 842
rect 1872 842 1884 844
rect 1872 834 1874 842
rect 1882 834 1884 842
rect 1902 842 1914 844
rect 1902 834 1904 842
rect 1912 834 1914 842
rect 1932 842 1944 844
rect 1932 834 1934 842
rect 1942 834 1944 842
rect 1962 842 1974 844
rect 1962 834 1964 842
rect 1972 834 1974 842
rect 1722 832 1744 834
rect 1752 832 1774 834
rect 1782 832 1804 834
rect 1812 832 1834 834
rect 1842 832 1864 834
rect 1872 832 1894 834
rect 1902 832 1924 834
rect 1932 832 1954 834
rect 1962 832 1984 834
tri 1066 824 1074 832 se
rect 1074 824 1084 832
rect 1352 824 1360 832
tri 1360 824 1368 832 nw
tri 1376 824 1384 832 se
rect 1384 824 1394 832
rect 1652 824 1662 832
tri 1662 824 1670 832 nw
tri 1678 824 1686 832 se
rect 1686 824 1694 832
rect 1732 824 1734 832
rect 1742 824 1744 832
rect 1762 824 1764 832
rect 1772 824 1774 832
rect 1792 824 1794 832
rect 1802 824 1804 832
rect 1822 824 1824 832
rect 1832 824 1834 832
rect 1852 824 1854 832
rect 1862 824 1864 832
rect 1882 824 1884 832
rect 1892 824 1894 832
rect 1912 824 1914 832
rect 1922 824 1924 832
rect 1942 824 1944 832
rect 1952 824 1954 832
rect 1972 824 1974 832
rect 1982 824 1984 832
tri 1064 822 1066 824 se
rect 1066 822 1084 824
rect 1342 822 1358 824
tri 1358 822 1360 824 nw
tri 1374 822 1376 824 se
rect 1376 822 1394 824
rect 1642 822 1660 824
tri 1660 822 1662 824 nw
tri 1676 822 1678 824 se
rect 1678 822 1694 824
rect 1722 822 1744 824
rect 1752 822 1774 824
rect 1782 822 1804 824
rect 1812 822 1834 824
rect 1842 822 1864 824
rect 1872 822 1894 824
rect 1902 822 1924 824
rect 1932 822 1954 824
rect 1962 822 1984 824
tri 1056 814 1064 822 se
rect 1064 814 1074 822
rect 1342 814 1350 822
tri 1350 814 1358 822 nw
tri 1366 814 1374 822 se
rect 1374 814 1384 822
rect 1642 814 1652 822
tri 1652 814 1660 822 nw
tri 1668 814 1676 822 se
rect 1676 814 1684 822
rect 1722 814 1724 822
rect 1732 814 1734 822
rect 1752 814 1754 822
rect 1762 814 1764 822
rect 1782 814 1784 822
rect 1792 814 1794 822
rect 1812 814 1814 822
rect 1822 814 1824 822
rect 1842 814 1844 822
rect 1852 814 1854 822
rect 1872 814 1874 822
rect 1882 814 1884 822
rect 1902 814 1904 822
rect 1912 814 1914 822
rect 1932 814 1934 822
rect 1942 814 1944 822
rect 1962 814 1964 822
rect 1972 814 1974 822
tri 1054 812 1056 814 se
rect 1056 812 1074 814
rect 1332 812 1348 814
tri 1348 812 1350 814 nw
tri 1364 812 1366 814 se
rect 1366 812 1384 814
rect 1632 812 1650 814
tri 1650 812 1652 814 nw
tri 1666 812 1668 814 se
rect 1668 812 1684 814
rect 1692 812 1704 814
rect 1722 812 1744 814
rect 1752 812 1774 814
rect 1782 812 1804 814
rect 1812 812 1834 814
rect 1842 812 1864 814
rect 1872 812 1894 814
rect 1902 812 1924 814
rect 1932 812 1954 814
rect 1962 812 1984 814
tri 1046 804 1054 812 se
rect 1054 804 1064 812
rect 1332 804 1340 812
tri 1340 804 1348 812 nw
tri 1356 804 1364 812 se
rect 1364 804 1374 812
rect 1632 804 1642 812
tri 1642 804 1650 812 nw
tri 1658 804 1666 812 se
rect 1666 804 1674 812
rect 1692 804 1694 812
rect 1702 804 1704 812
rect 1732 804 1734 812
rect 1742 804 1744 812
rect 1762 804 1764 812
rect 1772 804 1774 812
rect 1792 804 1794 812
rect 1802 804 1804 812
rect 1822 804 1824 812
rect 1832 804 1834 812
rect 1852 804 1854 812
rect 1862 804 1864 812
rect 1882 804 1884 812
rect 1892 804 1894 812
rect 1912 804 1914 812
rect 1922 804 1924 812
rect 1942 804 1944 812
rect 1952 804 1954 812
rect 1972 804 1974 812
rect 1982 804 1984 812
tri 1044 802 1046 804 se
rect 1046 802 1064 804
rect 1322 802 1338 804
tri 1338 802 1340 804 nw
tri 1354 802 1356 804 se
rect 1356 802 1374 804
rect 1622 802 1640 804
tri 1640 802 1642 804 nw
tri 1656 802 1658 804 se
rect 1658 802 1674 804
rect 1682 802 1704 804
rect 1722 802 1744 804
rect 1752 802 1774 804
rect 1782 802 1804 804
rect 1812 802 1834 804
rect 1842 802 1864 804
rect 1872 802 1894 804
rect 1902 802 1924 804
rect 1932 802 1954 804
rect 1962 802 1984 804
tri 1036 794 1044 802 se
rect 1044 794 1054 802
rect 1322 794 1330 802
tri 1330 794 1338 802 nw
tri 1346 794 1354 802 se
rect 1354 794 1364 802
rect 1622 794 1632 802
tri 1632 794 1640 802 nw
tri 1648 794 1656 802 se
rect 1656 794 1664 802
rect 1682 794 1684 802
rect 1692 794 1694 802
rect 1722 794 1724 802
rect 1732 794 1734 802
rect 1752 794 1754 802
rect 1762 794 1764 802
rect 1782 794 1784 802
rect 1792 794 1794 802
rect 1812 794 1814 802
rect 1822 794 1824 802
rect 1842 794 1844 802
rect 1852 794 1854 802
rect 1872 794 1874 802
rect 1882 794 1884 802
rect 1902 794 1904 802
rect 1912 794 1914 802
rect 1932 794 1934 802
rect 1942 794 1944 802
rect 1962 794 1964 802
rect 1972 794 1974 802
tri 1034 792 1036 794 se
rect 1036 792 1054 794
rect 1312 792 1328 794
tri 1328 792 1330 794 nw
tri 1344 792 1346 794 se
rect 1346 792 1364 794
rect 1612 792 1630 794
tri 1630 792 1632 794 nw
tri 1646 792 1648 794 se
rect 1648 792 1664 794
rect 1672 792 1704 794
rect 1722 792 1744 794
rect 1752 792 1774 794
rect 1782 792 1804 794
rect 1812 792 1834 794
rect 1842 792 1864 794
rect 1872 792 1894 794
rect 1902 792 1924 794
rect 1932 792 1954 794
rect 1962 792 1984 794
tri 1026 784 1034 792 se
rect 1034 784 1044 792
rect 1312 784 1320 792
tri 1320 784 1328 792 nw
tri 1336 784 1344 792 se
rect 1344 784 1354 792
rect 1612 784 1622 792
tri 1622 784 1630 792 nw
tri 1638 784 1646 792 se
rect 1646 784 1654 792
rect 1672 784 1674 792
rect 1682 784 1684 792
rect 1692 784 1694 792
rect 1702 784 1704 792
rect 1732 784 1734 792
rect 1742 784 1744 792
rect 1762 784 1764 792
rect 1772 784 1774 792
rect 1792 784 1794 792
rect 1802 784 1804 792
rect 1822 784 1824 792
rect 1832 784 1834 792
rect 1852 784 1854 792
rect 1862 784 1864 792
rect 1882 784 1884 792
rect 1892 784 1894 792
rect 1912 784 1914 792
rect 1922 784 1924 792
rect 1942 784 1944 792
rect 1952 784 1954 792
rect 1972 784 1974 792
rect 1982 784 1984 792
tri 1024 782 1026 784 se
rect 1026 782 1044 784
rect 1302 782 1318 784
tri 1318 782 1320 784 nw
tri 1334 782 1336 784 se
rect 1336 782 1354 784
rect 1602 782 1620 784
tri 1620 782 1622 784 nw
tri 1636 782 1638 784 se
rect 1638 782 1654 784
rect 1662 782 1704 784
rect 1722 782 1744 784
rect 1752 782 1774 784
rect 1782 782 1804 784
rect 1812 782 1834 784
rect 1842 782 1864 784
rect 1872 782 1894 784
rect 1902 782 1924 784
rect 1932 782 1954 784
rect 1962 782 1984 784
tri 1016 774 1024 782 se
rect 1024 774 1034 782
rect 1302 774 1310 782
tri 1310 774 1318 782 nw
tri 1326 774 1334 782 se
rect 1334 774 1344 782
rect 1602 774 1612 782
tri 1612 774 1620 782 nw
tri 1628 774 1636 782 se
rect 1636 774 1644 782
rect 1662 774 1664 782
rect 1672 774 1674 782
rect 1682 774 1684 782
rect 1692 774 1694 782
tri 1014 772 1016 774 se
rect 1016 772 1034 774
rect 1292 772 1308 774
tri 1308 772 1310 774 nw
tri 1324 772 1326 774 se
rect 1326 772 1344 774
rect 1592 772 1610 774
tri 1610 772 1612 774 nw
tri 1626 772 1628 774 se
rect 1628 772 1644 774
rect 1652 772 1694 774
rect 1722 774 1724 782
rect 1732 774 1734 782
rect 1752 774 1754 782
rect 1762 774 1764 782
rect 1782 774 1784 782
rect 1792 774 1794 782
rect 1812 774 1814 782
rect 1822 774 1824 782
rect 1842 774 1844 782
rect 1852 774 1854 782
rect 1872 774 1874 782
rect 1882 774 1884 782
rect 1902 774 1904 782
rect 1912 774 1914 782
rect 1932 774 1934 782
rect 1942 774 1944 782
rect 1962 774 1964 782
rect 1972 774 1974 782
rect 1722 772 1744 774
rect 1752 772 1774 774
rect 1782 772 1804 774
rect 1812 772 1834 774
rect 1842 772 1864 774
rect 1872 772 1894 774
rect 1902 772 1924 774
rect 1932 772 1954 774
rect 1962 772 1984 774
tri 1006 764 1014 772 se
rect 1014 764 1024 772
rect 1292 764 1300 772
tri 1300 764 1308 772 nw
tri 1316 764 1324 772 se
rect 1324 764 1334 772
rect 1592 764 1602 772
tri 1602 764 1610 772 nw
tri 1618 764 1626 772 se
rect 1626 764 1634 772
rect 1652 764 1654 772
rect 1662 764 1664 772
rect 1672 764 1674 772
rect 1682 764 1684 772
rect 1732 764 1734 772
rect 1742 764 1744 772
rect 1762 764 1764 772
rect 1772 764 1774 772
rect 1792 764 1794 772
rect 1802 764 1804 772
rect 1822 764 1824 772
rect 1832 764 1834 772
rect 1852 764 1854 772
rect 1862 764 1864 772
rect 1882 764 1884 772
rect 1892 764 1894 772
rect 1912 764 1914 772
rect 1922 764 1924 772
rect 1942 764 1944 772
rect 1952 764 1954 772
rect 1972 764 1974 772
rect 1982 764 1984 772
tri 1004 762 1006 764 se
rect 1006 762 1024 764
rect 1282 762 1298 764
tri 1298 762 1300 764 nw
tri 1314 762 1316 764 se
rect 1316 762 1334 764
rect 1582 762 1600 764
tri 1600 762 1602 764 nw
tri 1616 762 1618 764 se
rect 1618 762 1634 764
rect 1642 762 1684 764
rect 1692 762 1704 764
tri 996 754 1004 762 se
rect 1004 754 1014 762
rect 1282 754 1290 762
tri 1290 754 1298 762 nw
tri 1306 754 1314 762 se
rect 1314 754 1324 762
rect 1582 754 1592 762
tri 1592 754 1600 762 nw
tri 1608 754 1616 762 se
rect 1616 754 1624 762
rect 1642 754 1644 762
rect 1652 754 1654 762
rect 1662 754 1664 762
rect 1672 754 1674 762
rect 1692 754 1694 762
rect 1702 754 1704 762
tri 994 752 996 754 se
rect 996 752 1014 754
rect 1272 752 1288 754
tri 1288 752 1290 754 nw
tri 1304 752 1306 754 se
rect 1306 752 1324 754
rect 1572 752 1590 754
tri 1590 752 1592 754 nw
tri 1606 752 1608 754 se
rect 1608 752 1624 754
rect 1632 752 1674 754
rect 1682 752 1704 754
rect 1722 762 1744 764
rect 1752 762 1774 764
rect 1782 762 1804 764
rect 1812 762 1834 764
rect 1842 762 1864 764
rect 1872 762 1894 764
rect 1902 762 1924 764
rect 1932 762 1954 764
rect 1962 762 1984 764
rect 1722 754 1724 762
rect 1732 754 1734 762
rect 1752 754 1754 762
rect 1762 754 1764 762
rect 1782 754 1784 762
rect 1792 754 1794 762
rect 1812 754 1814 762
rect 1822 754 1824 762
rect 1842 754 1844 762
rect 1852 754 1854 762
rect 1872 754 1874 762
rect 1882 754 1884 762
rect 1902 754 1904 762
rect 1912 754 1914 762
rect 1932 754 1934 762
rect 1942 754 1944 762
rect 1962 754 1964 762
rect 1972 754 1974 762
rect 1722 752 1744 754
rect 1752 752 1774 754
rect 1782 752 1804 754
rect 1812 752 1834 754
rect 1842 752 1864 754
rect 1872 752 1894 754
rect 1902 752 1924 754
rect 1932 752 1954 754
rect 1962 752 1984 754
tri 986 744 994 752 se
rect 994 744 1004 752
rect 1272 744 1280 752
tri 1280 744 1288 752 nw
tri 1296 744 1304 752 se
rect 1304 744 1314 752
rect 1572 744 1582 752
tri 1582 744 1590 752 nw
tri 1598 744 1606 752 se
rect 1606 744 1614 752
rect 1632 744 1634 752
rect 1642 744 1644 752
rect 1652 744 1654 752
rect 1662 744 1664 752
rect 1682 744 1684 752
rect 1692 744 1694 752
rect 1732 744 1734 752
rect 1742 744 1744 752
rect 1762 744 1764 752
rect 1772 744 1774 752
rect 1792 744 1794 752
rect 1802 744 1804 752
rect 1822 744 1824 752
rect 1832 744 1834 752
rect 1852 744 1854 752
rect 1862 744 1864 752
rect 1882 744 1884 752
rect 1892 744 1894 752
rect 1912 744 1914 752
rect 1922 744 1924 752
rect 1942 744 1944 752
rect 1952 744 1954 752
rect 1972 744 1974 752
rect 1982 744 1984 752
tri 984 742 986 744 se
rect 986 742 1004 744
rect 1262 742 1278 744
tri 1278 742 1280 744 nw
tri 1294 742 1296 744 se
rect 1296 742 1314 744
rect 1562 742 1580 744
tri 1580 742 1582 744 nw
tri 1596 742 1598 744 se
rect 1598 742 1614 744
rect 1622 742 1664 744
rect 1672 742 1694 744
rect 1722 742 1744 744
rect 1752 742 1774 744
rect 1782 742 1804 744
rect 1812 742 1834 744
rect 1842 742 1864 744
rect 1872 742 1894 744
rect 1902 742 1924 744
rect 1932 742 1954 744
rect 1962 742 1984 744
tri 976 734 984 742 se
rect 984 734 994 742
rect 1262 734 1270 742
tri 1270 734 1278 742 nw
tri 1286 734 1294 742 se
rect 1294 734 1304 742
rect 1562 734 1572 742
tri 1572 734 1580 742 nw
tri 1588 734 1596 742 se
rect 1596 734 1604 742
rect 1622 734 1624 742
rect 1632 734 1634 742
rect 1642 734 1644 742
rect 1652 734 1654 742
rect 1672 734 1674 742
rect 1682 734 1684 742
tri 974 732 976 734 se
rect 976 732 994 734
rect 1252 732 1268 734
tri 1268 732 1270 734 nw
tri 1284 732 1286 734 se
rect 1286 732 1304 734
rect 1552 732 1570 734
tri 1570 732 1572 734 nw
tri 1586 732 1588 734 se
rect 1588 732 1604 734
rect 1612 732 1654 734
rect 1662 732 1684 734
rect 1722 734 1724 742
rect 1732 734 1734 742
rect 1752 734 1754 742
rect 1762 734 1764 742
rect 1782 734 1784 742
rect 1792 734 1794 742
rect 1812 734 1814 742
rect 1822 734 1824 742
rect 1842 734 1844 742
rect 1852 734 1854 742
rect 1872 734 1874 742
rect 1882 734 1884 742
rect 1902 734 1904 742
rect 1912 734 1914 742
rect 1932 734 1934 742
rect 1942 734 1944 742
rect 1962 734 1964 742
rect 1972 734 1974 742
rect 1722 732 1744 734
rect 1752 732 1774 734
rect 1782 732 1804 734
rect 1812 732 1834 734
rect 1842 732 1864 734
rect 1872 732 1894 734
rect 1902 732 1924 734
rect 1932 732 1954 734
rect 1962 732 1984 734
tri 966 724 974 732 se
rect 974 724 984 732
rect 1252 724 1260 732
tri 1260 724 1268 732 nw
tri 1276 724 1284 732 se
rect 1284 724 1294 732
rect 1552 724 1562 732
tri 1562 724 1570 732 nw
tri 1578 724 1586 732 se
rect 1586 724 1594 732
rect 1612 724 1614 732
rect 1622 724 1624 732
rect 1632 724 1634 732
rect 1642 724 1644 732
rect 1662 724 1664 732
rect 1672 724 1674 732
rect 1732 724 1734 732
rect 1742 724 1744 732
rect 1762 724 1764 732
rect 1772 724 1774 732
rect 1792 724 1794 732
rect 1802 724 1804 732
rect 1822 724 1824 732
rect 1832 724 1834 732
rect 1852 724 1854 732
rect 1862 724 1864 732
rect 1882 724 1884 732
rect 1892 724 1894 732
rect 1912 724 1914 732
rect 1922 724 1924 732
rect 1942 724 1944 732
rect 1952 724 1954 732
rect 1972 724 1974 732
rect 1982 724 1984 732
tri 964 722 966 724 se
rect 966 722 984 724
rect 1242 722 1258 724
tri 1258 722 1260 724 nw
tri 1274 722 1276 724 se
rect 1276 722 1294 724
rect 1542 722 1560 724
tri 1560 722 1562 724 nw
tri 1576 722 1578 724 se
rect 1578 722 1594 724
rect 1602 722 1644 724
rect 1652 722 1674 724
rect 1722 722 1744 724
rect 1752 722 1774 724
rect 1782 722 1804 724
rect 1812 722 1834 724
rect 1842 722 1864 724
rect 1872 722 1894 724
rect 1902 722 1924 724
rect 1932 722 1954 724
rect 1962 722 1984 724
tri 956 714 964 722 se
rect 964 714 974 722
rect 1242 714 1250 722
tri 1250 714 1258 722 nw
tri 1266 714 1274 722 se
rect 1274 714 1284 722
rect 1542 714 1552 722
tri 1552 714 1560 722 nw
tri 1568 714 1576 722 se
rect 1576 714 1584 722
rect 1602 714 1604 722
rect 1612 714 1614 722
rect 1622 714 1624 722
rect 1632 714 1634 722
rect 1652 714 1654 722
rect 1662 714 1664 722
tri 954 712 956 714 se
rect 956 712 974 714
rect 1232 712 1248 714
tri 1248 712 1250 714 nw
tri 1264 712 1266 714 se
rect 1266 712 1284 714
rect 1532 712 1550 714
tri 1550 712 1552 714 nw
tri 1566 712 1568 714 se
rect 1568 712 1584 714
rect 1592 712 1634 714
rect 1642 712 1664 714
rect 1722 714 1724 722
rect 1732 714 1734 722
rect 1752 714 1754 722
rect 1762 714 1764 722
rect 1782 714 1784 722
rect 1792 714 1794 722
rect 1812 714 1814 722
rect 1822 714 1824 722
rect 1842 714 1844 722
rect 1852 714 1854 722
rect 1872 714 1874 722
rect 1882 714 1884 722
rect 1902 714 1904 722
rect 1912 714 1914 722
rect 1932 714 1934 722
rect 1942 714 1944 722
rect 1962 714 1964 722
rect 1972 714 1974 722
rect 1722 712 1744 714
rect 1752 712 1774 714
rect 1782 712 1804 714
rect 1812 712 1834 714
rect 1842 712 1864 714
rect 1872 712 1894 714
rect 1902 712 1924 714
rect 1932 712 1954 714
rect 1962 712 1984 714
tri 946 704 954 712 se
rect 954 704 964 712
rect 1232 704 1240 712
tri 1240 704 1248 712 nw
tri 1256 704 1264 712 se
rect 1264 704 1274 712
rect 1532 704 1542 712
tri 1542 704 1550 712 nw
tri 1558 704 1566 712 se
rect 1566 704 1574 712
rect 1592 704 1594 712
rect 1602 704 1604 712
rect 1612 704 1614 712
rect 1622 704 1624 712
rect 1642 704 1644 712
rect 1652 704 1654 712
rect 1732 704 1734 712
rect 1742 704 1744 712
rect 1762 704 1764 712
rect 1772 704 1774 712
rect 1792 704 1794 712
rect 1802 704 1804 712
rect 1822 704 1824 712
rect 1832 704 1834 712
rect 1852 704 1854 712
rect 1862 704 1864 712
rect 1882 704 1884 712
rect 1892 704 1894 712
rect 1912 704 1914 712
rect 1922 704 1924 712
rect 1942 704 1944 712
rect 1952 704 1954 712
rect 1972 704 1974 712
rect 1982 704 1984 712
tri 944 702 946 704 se
rect 946 702 964 704
rect 1222 702 1238 704
tri 1238 702 1240 704 nw
tri 1254 702 1256 704 se
rect 1256 702 1274 704
rect 1522 702 1540 704
tri 1540 702 1542 704 nw
tri 1556 702 1558 704 se
rect 1558 702 1574 704
rect 1582 702 1624 704
rect 1632 702 1654 704
rect 1692 702 1704 704
tri 936 694 944 702 se
rect 944 694 954 702
rect 1222 694 1230 702
tri 1230 694 1238 702 nw
tri 1250 698 1254 702 se
rect 1254 698 1264 702
tri 1246 694 1250 698 se
rect 1250 694 1264 698
rect 1522 698 1536 702
tri 1536 698 1540 702 nw
tri 1552 698 1556 702 se
rect 1556 698 1564 702
rect 1522 694 1532 698
tri 1532 694 1536 698 nw
tri 1548 694 1552 698 se
rect 1552 694 1564 698
rect 1582 694 1584 702
rect 1592 694 1594 702
rect 1602 694 1604 702
rect 1612 694 1614 702
tri 934 692 936 694 se
rect 936 692 954 694
rect 1212 692 1228 694
tri 1228 692 1230 694 nw
tri 1244 692 1246 694 se
rect 1246 692 1264 694
rect 1512 692 1530 694
tri 1530 692 1532 694 nw
tri 1546 692 1548 694 se
rect 1548 692 1564 694
rect 1572 692 1624 694
tri 926 684 934 692 se
rect 934 684 944 692
rect 1212 690 1226 692
tri 1226 690 1228 692 nw
tri 1242 690 1244 692 se
rect 1244 690 1254 692
rect 1212 684 1220 690
tri 1220 684 1226 690 nw
tri 1236 684 1242 690 se
rect 1242 684 1254 690
rect 1512 684 1522 692
tri 1522 684 1530 692 nw
tri 1538 684 1546 692 se
rect 1546 684 1554 692
rect 1572 684 1574 692
rect 1582 684 1584 692
rect 1592 684 1594 692
rect 1602 684 1604 692
rect 1612 684 1614 692
rect 1622 684 1624 692
rect 1632 684 1634 702
rect 1642 684 1644 702
rect 1692 694 1694 702
rect 1702 694 1704 702
rect 1722 702 1744 704
rect 1752 702 1774 704
rect 1782 702 1804 704
rect 1812 702 1834 704
rect 1842 702 1864 704
rect 1872 702 1894 704
rect 1902 702 1924 704
rect 1932 702 1954 704
rect 1962 702 1984 704
rect 1682 692 1714 694
rect 1682 684 1684 692
rect 1692 684 1694 692
rect 1702 684 1704 692
rect 1712 684 1714 692
rect 1722 684 1724 702
rect 1732 684 1734 702
rect 1752 694 1754 702
rect 1762 694 1764 702
rect 1782 694 1784 702
rect 1792 694 1794 702
rect 1812 694 1814 702
rect 1822 694 1824 702
rect 1842 694 1844 702
rect 1852 694 1854 702
rect 1872 694 1874 702
rect 1882 694 1884 702
rect 1902 694 1904 702
rect 1912 694 1914 702
rect 1932 694 1934 702
rect 1942 694 1944 702
rect 1962 694 1964 702
rect 1972 694 1974 702
rect 1992 694 2000 1332
rect 1742 692 1774 694
rect 1742 684 1744 692
rect 1752 684 1754 692
rect 1762 684 1764 692
rect 1772 684 1774 692
rect 1782 688 2000 694
rect 1782 684 1786 688
tri 1786 684 1790 688 nw
tri 924 682 926 684 se
rect 926 682 944 684
rect 1202 682 1218 684
tri 1218 682 1220 684 nw
tri 1234 682 1236 684 se
rect 1236 682 1254 684
rect 1502 682 1520 684
tri 1520 682 1522 684 nw
tri 1536 682 1538 684 se
rect 1538 682 1554 684
rect 1562 682 1644 684
rect 1672 682 1784 684
tri 1784 682 1786 684 nw
tri 916 674 924 682 se
rect 924 674 934 682
rect 1202 674 1210 682
tri 1210 674 1218 682 nw
tri 1226 674 1234 682 se
rect 1234 674 1244 682
rect 1502 674 1512 682
tri 1512 674 1520 682 nw
tri 1528 674 1536 682 se
rect 1536 674 1544 682
rect 1562 674 1564 682
rect 1572 674 1574 682
rect 1582 674 1584 682
rect 1592 674 1594 682
rect 1602 674 1604 682
rect 1612 674 1614 682
rect 1622 674 1624 682
rect 1632 674 1634 682
rect 1672 674 1674 682
rect 1682 674 1684 682
rect 1692 674 1694 682
rect 1702 674 1704 682
rect 1712 674 1714 682
rect 1722 674 1724 682
rect 1732 674 1734 682
rect 1742 674 1744 682
rect 1752 674 1754 682
rect 1762 674 1764 682
rect 1772 674 1776 682
tri 1776 674 1784 682 nw
tri 914 672 916 674 se
rect 916 672 934 674
rect 1192 672 1208 674
tri 1208 672 1210 674 nw
tri 1224 672 1226 674 se
rect 1226 672 1244 674
rect 1492 672 1510 674
tri 1510 672 1512 674 nw
tri 1526 672 1528 674 se
rect 1528 672 1544 674
rect 1552 672 1634 674
rect 1662 672 1774 674
tri 1774 672 1776 674 nw
tri 906 664 914 672 se
rect 914 664 924 672
rect 1192 664 1200 672
tri 1200 664 1208 672 nw
tri 1216 664 1224 672 se
rect 1224 664 1234 672
rect 1492 664 1502 672
tri 1502 664 1510 672 nw
tri 1518 664 1526 672 se
rect 1526 664 1534 672
rect 1552 664 1554 672
rect 1562 664 1564 672
rect 1572 664 1574 672
rect 1582 664 1584 672
rect 1592 664 1594 672
rect 1602 664 1604 672
rect 1612 664 1614 672
rect 1622 664 1624 672
rect 1662 664 1664 672
rect 1672 664 1674 672
rect 1682 664 1684 672
rect 1692 664 1694 672
rect 1702 664 1704 672
rect 1712 664 1714 672
rect 1722 664 1724 672
rect 1732 664 1734 672
rect 1742 664 1744 672
rect 1752 664 1754 672
rect 1762 664 1766 672
tri 1766 664 1774 672 nw
tri 904 662 906 664 se
rect 906 662 924 664
rect 1182 662 1198 664
tri 1198 662 1200 664 nw
tri 1214 662 1216 664 se
rect 1216 662 1234 664
rect 1482 662 1500 664
tri 1500 662 1502 664 nw
tri 1516 662 1518 664 se
rect 1518 662 1534 664
rect 1542 662 1624 664
rect 1652 662 1764 664
tri 1764 662 1766 664 nw
tri 896 654 904 662 se
rect 904 654 914 662
rect 1182 654 1190 662
tri 1190 654 1198 662 nw
tri 1206 654 1214 662 se
rect 1214 654 1224 662
rect 1482 660 1498 662
tri 1498 660 1500 662 nw
tri 1514 660 1516 662 se
rect 1516 660 1524 662
rect 1482 654 1492 660
tri 1492 654 1498 660 nw
tri 1508 654 1514 660 se
rect 1514 654 1524 660
rect 1542 654 1544 662
rect 1552 654 1554 662
rect 1562 654 1564 662
rect 1572 654 1574 662
rect 1582 654 1584 662
rect 1592 654 1594 662
rect 1602 654 1604 662
rect 1612 654 1614 662
rect 1652 654 1654 662
rect 1662 654 1664 662
rect 1672 654 1674 662
rect 1682 654 1684 662
rect 1692 654 1694 662
rect 1702 654 1704 662
rect 1712 654 1714 662
rect 1722 654 1724 662
rect 1732 654 1734 662
rect 1742 654 1744 662
rect 1752 654 1756 662
tri 1756 654 1764 662 nw
tri 894 652 896 654 se
rect 896 652 914 654
rect 1172 652 1188 654
tri 1188 652 1190 654 nw
tri 1204 652 1206 654 se
rect 1206 652 1224 654
rect 1472 652 1490 654
tri 1490 652 1492 654 nw
tri 1506 652 1508 654 se
rect 1508 652 1524 654
rect 1532 652 1614 654
rect 1642 652 1754 654
tri 1754 652 1756 654 nw
tri 886 644 894 652 se
rect 894 644 904 652
rect 1172 644 1180 652
tri 1180 644 1188 652 nw
tri 1196 644 1204 652 se
rect 1204 644 1214 652
rect 1472 644 1482 652
tri 1482 644 1490 652 nw
tri 1498 644 1506 652 se
rect 1506 644 1514 652
rect 1532 644 1534 652
rect 1542 644 1544 652
rect 1552 644 1554 652
rect 1562 644 1564 652
rect 1572 644 1574 652
rect 1582 644 1584 652
rect 1592 644 1594 652
rect 1602 644 1604 652
rect 1642 644 1644 652
rect 1652 644 1654 652
rect 1662 644 1664 652
rect 1672 644 1674 652
rect 1682 644 1684 652
rect 1692 644 1694 652
rect 1702 644 1704 652
rect 1712 644 1714 652
rect 1722 644 1724 652
rect 1732 644 1734 652
rect 1742 644 1746 652
tri 1746 644 1754 652 nw
tri 1814 644 1822 652 se
rect 1822 644 2000 652
tri 884 642 886 644 se
rect 886 642 904 644
rect 1162 642 1178 644
tri 1178 642 1180 644 nw
tri 1194 642 1196 644 se
rect 1196 642 1214 644
rect 1462 642 1480 644
tri 1480 642 1482 644 nw
tri 1496 642 1498 644 se
rect 1498 642 1514 644
rect 1522 642 1604 644
rect 1632 642 1744 644
tri 1744 642 1746 644 nw
tri 1812 642 1814 644 se
rect 1814 642 2000 644
tri 876 634 884 642 se
rect 884 634 894 642
rect 1162 634 1170 642
tri 1170 634 1178 642 nw
tri 1186 634 1194 642 se
rect 1194 634 1204 642
rect 1462 634 1472 642
tri 1472 634 1480 642 nw
tri 1488 634 1496 642 se
rect 1496 634 1504 642
rect 1522 634 1524 642
rect 1532 634 1534 642
rect 1542 634 1544 642
rect 1552 634 1554 642
rect 1562 634 1564 642
rect 1572 634 1574 642
rect 1582 634 1584 642
rect 1592 634 1594 642
rect 1632 634 1634 642
rect 1642 634 1644 642
rect 1652 634 1654 642
rect 1662 634 1664 642
rect 1672 634 1674 642
rect 1682 634 1684 642
rect 1692 634 1694 642
rect 1702 634 1704 642
rect 1712 634 1714 642
rect 1722 634 1724 642
rect 1732 634 1736 642
tri 1736 634 1744 642 nw
tri 1804 634 1812 642 se
rect 1812 634 1820 642
tri 874 632 876 634 se
rect 876 632 894 634
rect 1152 632 1168 634
tri 1168 632 1170 634 nw
tri 1184 632 1186 634 se
rect 1186 632 1204 634
rect 1452 632 1470 634
tri 1470 632 1472 634 nw
tri 1486 632 1488 634 se
rect 1488 632 1504 634
rect 1512 632 1594 634
rect 1622 632 1734 634
tri 1734 632 1736 634 nw
tri 1802 632 1804 634 se
rect 1804 632 1820 634
rect 1828 634 1830 642
rect 1838 634 1840 642
rect 1858 634 1860 642
rect 1868 634 1870 642
rect 1888 634 1890 642
rect 1898 634 1900 642
rect 1918 634 1920 642
rect 1928 634 1930 642
rect 1948 634 1950 642
rect 1958 634 1960 642
rect 1978 634 1980 642
rect 1988 634 1990 642
rect 1998 634 2000 642
rect 1828 632 1850 634
rect 1858 632 1880 634
rect 1888 632 1910 634
rect 1918 632 1940 634
rect 1948 632 1970 634
rect 1978 632 2000 634
tri 866 624 874 632 se
rect 874 624 884 632
rect 1152 624 1160 632
tri 1160 624 1168 632 nw
tri 1176 624 1184 632 se
rect 1184 624 1194 632
rect 1452 624 1462 632
tri 1462 624 1470 632 nw
tri 1478 624 1486 632 se
rect 1486 624 1494 632
rect 1512 624 1514 632
rect 1522 624 1524 632
rect 1532 624 1534 632
rect 1542 624 1544 632
rect 1552 624 1554 632
rect 1562 624 1564 632
rect 1572 624 1574 632
rect 1582 624 1584 632
rect 1622 624 1624 632
rect 1632 624 1634 632
rect 1642 624 1644 632
rect 1652 624 1654 632
rect 1662 624 1664 632
rect 1672 624 1674 632
rect 1682 624 1684 632
rect 1692 624 1694 632
rect 1702 624 1704 632
rect 1712 624 1714 632
rect 1722 628 1730 632
tri 1730 628 1734 632 nw
tri 1798 628 1802 632 se
rect 1802 628 1810 632
rect 1722 624 1726 628
tri 1726 624 1730 628 nw
tri 1794 624 1798 628 se
rect 1798 624 1810 628
rect 1838 624 1840 632
rect 1848 624 1850 632
rect 1868 624 1870 632
rect 1878 624 1880 632
rect 1898 624 1900 632
rect 1908 624 1910 632
rect 1928 624 1930 632
rect 1938 624 1940 632
rect 1958 624 1960 632
rect 1968 624 1970 632
rect 1988 624 1990 632
rect 1998 624 2000 632
tri 864 622 866 624 se
rect 866 622 884 624
rect 1142 622 1158 624
tri 1158 622 1160 624 nw
tri 1174 622 1176 624 se
rect 1176 622 1194 624
rect 1442 622 1460 624
tri 1460 622 1462 624 nw
tri 1476 622 1478 624 se
rect 1478 622 1494 624
rect 1502 622 1584 624
rect 1612 622 1724 624
tri 1724 622 1726 624 nw
tri 1792 622 1794 624 se
rect 1794 622 1810 624
rect 1828 622 1850 624
rect 1858 622 1880 624
rect 1888 622 1910 624
rect 1918 622 1940 624
rect 1948 622 1970 624
rect 1978 622 2000 624
tri 856 614 864 622 se
rect 864 614 874 622
rect 1142 614 1150 622
tri 1150 614 1158 622 nw
tri 1166 614 1174 622 se
rect 1174 614 1184 622
rect 1442 614 1452 622
tri 1452 614 1460 622 nw
tri 1468 614 1476 622 se
rect 1476 614 1484 622
rect 1502 614 1504 622
rect 1512 614 1514 622
rect 1522 614 1524 622
rect 1532 614 1534 622
rect 1542 614 1544 622
rect 1552 614 1554 622
rect 1562 614 1564 622
rect 1572 614 1574 622
rect 1612 614 1614 622
rect 1622 614 1624 622
rect 1632 614 1634 622
rect 1642 614 1644 622
rect 1652 614 1654 622
rect 1662 614 1664 622
rect 1672 614 1674 622
rect 1682 614 1684 622
rect 1692 614 1694 622
rect 1702 614 1704 622
rect 1712 614 1716 622
tri 1716 614 1724 622 nw
tri 1784 614 1792 622 se
rect 1792 614 1800 622
rect 1828 614 1830 622
rect 1838 614 1840 622
rect 1858 614 1860 622
rect 1868 614 1870 622
rect 1888 614 1890 622
rect 1898 614 1900 622
rect 1918 614 1920 622
rect 1928 614 1930 622
rect 1948 614 1950 622
rect 1958 614 1960 622
rect 1978 614 1980 622
rect 1988 614 1990 622
rect 1998 614 2000 622
tri 854 612 856 614 se
rect 856 612 874 614
rect 1132 612 1148 614
tri 1148 612 1150 614 nw
tri 1164 612 1166 614 se
rect 1166 612 1184 614
rect 1432 612 1450 614
tri 1450 612 1452 614 nw
tri 1466 612 1468 614 se
rect 1468 612 1484 614
rect 1492 612 1574 614
rect 1602 612 1714 614
tri 1714 612 1716 614 nw
tri 1782 612 1784 614 se
rect 1784 612 1800 614
rect 1808 612 1820 614
rect 1828 612 1850 614
rect 1858 612 1880 614
rect 1888 612 1910 614
rect 1918 612 1940 614
rect 1948 612 1970 614
rect 1978 612 2000 614
tri 846 604 854 612 se
rect 854 604 864 612
rect 1132 604 1140 612
tri 1140 604 1148 612 nw
tri 1156 604 1164 612 se
rect 1164 604 1174 612
rect 1432 604 1442 612
tri 1442 604 1450 612 nw
tri 1458 604 1466 612 se
rect 1466 604 1474 612
rect 1492 604 1494 612
rect 1502 604 1504 612
rect 1512 604 1514 612
rect 1522 604 1524 612
rect 1532 604 1534 612
rect 1542 604 1544 612
rect 1552 604 1554 612
rect 1562 604 1564 612
rect 1602 604 1604 612
rect 1612 604 1614 612
rect 1622 604 1624 612
rect 1632 604 1634 612
rect 1642 604 1644 612
rect 1652 604 1654 612
rect 1662 604 1664 612
rect 1672 604 1674 612
rect 1682 604 1684 612
rect 1692 604 1694 612
rect 1702 604 1706 612
tri 1706 604 1714 612 nw
tri 1774 604 1782 612 se
rect 1782 604 1790 612
rect 1808 604 1810 612
rect 1818 604 1820 612
rect 1838 604 1840 612
rect 1848 604 1850 612
rect 1868 604 1870 612
rect 1878 604 1880 612
rect 1898 604 1900 612
rect 1908 604 1910 612
rect 1928 604 1930 612
rect 1938 604 1940 612
rect 1958 604 1960 612
rect 1968 604 1970 612
rect 1988 604 1990 612
rect 1998 604 2000 612
tri 844 602 846 604 se
rect 846 602 864 604
rect 1122 602 1138 604
tri 1138 602 1140 604 nw
tri 1154 602 1156 604 se
rect 1156 602 1174 604
rect 1422 602 1440 604
tri 1440 602 1442 604 nw
tri 1456 602 1458 604 se
rect 1458 602 1474 604
rect 1482 602 1564 604
rect 1592 602 1704 604
tri 1704 602 1706 604 nw
tri 1772 602 1774 604 se
rect 1774 602 1790 604
rect 1798 602 1820 604
rect 1828 602 1850 604
rect 1858 602 1880 604
rect 1888 602 1910 604
rect 1918 602 1940 604
rect 1948 602 1970 604
rect 1978 602 2000 604
tri 836 594 844 602 se
rect 844 594 854 602
rect 1122 594 1130 602
tri 1130 594 1138 602 nw
tri 1146 594 1154 602 se
rect 1154 594 1164 602
rect 1422 594 1432 602
tri 1432 594 1440 602 nw
tri 1448 594 1456 602 se
rect 1456 594 1464 602
rect 1482 594 1484 602
rect 1492 594 1494 602
rect 1502 594 1504 602
rect 1512 594 1514 602
rect 1522 594 1524 602
rect 1532 594 1534 602
rect 1542 594 1544 602
rect 1552 594 1554 602
rect 1592 594 1594 602
rect 1602 594 1604 602
rect 1612 594 1614 602
rect 1622 594 1624 602
rect 1632 594 1634 602
rect 1642 594 1644 602
rect 1652 594 1654 602
rect 1662 594 1664 602
rect 1672 594 1674 602
rect 1682 594 1684 602
rect 1692 594 1696 602
tri 1696 594 1704 602 nw
tri 1764 594 1772 602 se
rect 1772 594 1780 602
rect 1798 594 1800 602
rect 1808 594 1810 602
tri 834 592 836 594 se
rect 836 592 854 594
rect 1112 592 1128 594
tri 1128 592 1130 594 nw
tri 1144 592 1146 594 se
rect 1146 592 1164 594
rect 1412 592 1430 594
tri 1430 592 1432 594 nw
tri 1446 592 1448 594 se
rect 1448 592 1464 594
rect 1472 592 1554 594
rect 1582 592 1694 594
tri 1694 592 1696 594 nw
tri 1762 592 1764 594 se
rect 1764 592 1780 594
rect 1788 592 1810 594
rect 1828 594 1830 602
rect 1838 594 1840 602
rect 1858 594 1860 602
rect 1868 594 1870 602
rect 1888 594 1890 602
rect 1898 594 1900 602
rect 1918 594 1920 602
rect 1928 594 1930 602
rect 1948 594 1950 602
rect 1958 594 1960 602
rect 1978 594 1980 602
rect 1988 594 1990 602
rect 1998 594 2000 602
rect 1828 592 1850 594
rect 1858 592 1880 594
rect 1888 592 1910 594
rect 1918 592 1940 594
rect 1948 592 1970 594
rect 1978 592 2000 594
tri 826 584 834 592 se
rect 834 584 844 592
rect 1112 584 1120 592
tri 1120 584 1128 592 nw
tri 1136 584 1144 592 se
rect 1144 584 1154 592
rect 1412 584 1422 592
tri 1422 584 1430 592 nw
tri 1438 584 1446 592 se
rect 1446 584 1454 592
rect 1472 584 1474 592
rect 1482 584 1484 592
rect 1492 584 1494 592
rect 1502 584 1504 592
rect 1512 584 1514 592
rect 1522 584 1524 592
rect 1532 584 1534 592
rect 1542 584 1544 592
rect 1582 584 1584 592
rect 1592 584 1594 592
rect 1602 584 1604 592
rect 1612 584 1614 592
rect 1622 584 1624 592
rect 1632 584 1634 592
rect 1642 584 1644 592
rect 1652 584 1654 592
rect 1662 584 1664 592
rect 1672 584 1674 592
rect 1682 584 1686 592
tri 1686 584 1694 592 nw
tri 1754 584 1762 592 se
rect 1762 584 1770 592
rect 1788 584 1790 592
rect 1798 584 1800 592
rect 1838 584 1840 592
rect 1848 584 1850 592
tri 824 582 826 584 se
rect 826 582 844 584
rect 1102 582 1118 584
tri 1118 582 1120 584 nw
tri 1134 582 1136 584 se
rect 1136 582 1154 584
rect 1402 582 1420 584
tri 1420 582 1422 584 nw
tri 1436 582 1438 584 se
rect 1438 582 1454 584
rect 1462 582 1544 584
rect 1572 582 1684 584
tri 1684 582 1686 584 nw
tri 1752 582 1754 584 se
rect 1754 582 1770 584
rect 1778 582 1800 584
rect 1808 582 1820 584
tri 816 574 824 582 se
rect 824 574 834 582
rect 1102 574 1110 582
tri 1110 574 1118 582 nw
tri 1126 574 1134 582 se
rect 1134 574 1144 582
rect 1402 574 1412 582
tri 1412 574 1420 582 nw
tri 1428 574 1436 582 se
rect 1436 574 1444 582
rect 1462 574 1464 582
rect 1472 574 1474 582
rect 1482 574 1484 582
rect 1492 574 1494 582
rect 1502 574 1504 582
rect 1512 574 1514 582
rect 1522 574 1524 582
rect 1532 574 1534 582
rect 1572 574 1574 582
rect 1582 574 1584 582
rect 1592 574 1594 582
rect 1602 574 1604 582
rect 1612 574 1614 582
rect 1622 574 1624 582
rect 1632 574 1634 582
rect 1642 574 1644 582
rect 1652 574 1654 582
rect 1662 574 1664 582
rect 1672 574 1676 582
tri 1676 574 1684 582 nw
tri 1744 574 1752 582 se
rect 1752 574 1760 582
rect 1778 574 1780 582
rect 1788 574 1790 582
rect 1808 574 1810 582
rect 1818 574 1820 582
tri 814 572 816 574 se
rect 816 572 834 574
rect 1092 572 1108 574
tri 1108 572 1110 574 nw
tri 1124 572 1126 574 se
rect 1126 572 1144 574
rect 1392 572 1410 574
tri 1410 572 1412 574 nw
tri 1426 572 1428 574 se
rect 1428 572 1444 574
rect 1452 572 1534 574
rect 1562 572 1674 574
tri 1674 572 1676 574 nw
tri 1742 572 1744 574 se
rect 1744 572 1760 574
rect 1768 572 1790 574
rect 1798 572 1820 574
rect 1828 582 1850 584
rect 1868 584 1870 592
rect 1878 584 1880 592
rect 1898 584 1900 592
rect 1908 584 1910 592
rect 1928 584 1930 592
rect 1938 584 1940 592
rect 1958 584 1960 592
rect 1968 584 1970 592
rect 1988 584 1990 592
rect 1998 584 2000 592
rect 1868 582 1880 584
rect 1888 582 1910 584
rect 1918 582 1940 584
rect 1948 582 1970 584
rect 1978 582 2000 584
rect 1828 574 1830 582
rect 1838 574 1840 582
rect 1888 574 1890 582
rect 1898 574 1900 582
rect 1918 574 1920 582
rect 1928 574 1930 582
rect 1948 574 1950 582
rect 1958 574 1960 582
rect 1978 574 1980 582
rect 1988 574 1990 582
rect 1998 574 2000 582
rect 1828 572 1840 574
rect 1868 572 1880 574
rect 1888 572 1910 574
rect 1918 572 1940 574
rect 1948 572 1970 574
rect 1978 572 2000 574
tri 806 564 814 572 se
rect 814 564 824 572
rect 1092 564 1100 572
tri 1100 564 1108 572 nw
tri 1116 564 1124 572 se
rect 1124 564 1134 572
rect 1392 564 1402 572
tri 1402 564 1410 572 nw
tri 1418 564 1426 572 se
rect 1426 564 1434 572
rect 1452 564 1454 572
rect 1462 564 1464 572
rect 1472 564 1474 572
rect 1482 564 1484 572
rect 1492 564 1494 572
rect 1502 564 1504 572
rect 1512 564 1514 572
rect 1522 564 1524 572
rect 1562 564 1564 572
rect 1572 564 1574 572
rect 1582 564 1584 572
rect 1592 564 1594 572
rect 1602 564 1604 572
rect 1612 564 1614 572
rect 1622 564 1624 572
rect 1632 564 1634 572
rect 1642 564 1644 572
rect 1652 564 1654 572
rect 1662 564 1666 572
tri 1666 564 1674 572 nw
tri 1734 564 1742 572 se
rect 1742 564 1750 572
rect 1768 564 1770 572
rect 1778 564 1780 572
rect 1798 564 1800 572
rect 1808 564 1810 572
rect 1868 564 1870 572
rect 1878 564 1880 572
rect 1898 564 1900 572
rect 1908 564 1910 572
rect 1928 564 1930 572
rect 1938 564 1940 572
rect 1958 564 1960 572
rect 1968 564 1970 572
rect 1988 564 1990 572
rect 1998 564 2000 572
tri 804 562 806 564 se
rect 806 562 824 564
rect 1082 562 1098 564
tri 1098 562 1100 564 nw
tri 1114 562 1116 564 se
rect 1116 562 1134 564
rect 1382 562 1400 564
tri 1400 562 1402 564 nw
tri 1416 562 1418 564 se
rect 1418 562 1434 564
rect 1442 562 1524 564
rect 1552 562 1664 564
tri 1664 562 1666 564 nw
tri 1732 562 1734 564 se
rect 1734 562 1750 564
rect 1758 562 1780 564
rect 1788 562 1810 564
rect 1858 562 1880 564
rect 1888 562 1910 564
rect 1918 562 1940 564
rect 1948 562 1970 564
rect 1978 562 2000 564
tri 796 554 804 562 se
rect 804 554 814 562
rect 1082 554 1090 562
tri 1090 554 1098 562 nw
tri 1106 554 1114 562 se
rect 1114 554 1124 562
rect 1382 554 1392 562
tri 1392 554 1400 562 nw
tri 1408 554 1416 562 se
rect 1416 554 1424 562
rect 1442 554 1444 562
rect 1452 554 1454 562
rect 1462 554 1464 562
rect 1472 554 1474 562
rect 1482 554 1484 562
rect 1492 554 1494 562
rect 1502 554 1504 562
rect 1512 554 1514 562
rect 1552 554 1554 562
rect 1562 554 1564 562
rect 1572 554 1574 562
rect 1582 554 1584 562
rect 1592 554 1594 562
rect 1602 554 1604 562
rect 1612 554 1614 562
rect 1622 554 1624 562
rect 1632 554 1634 562
rect 1642 554 1644 562
rect 1652 560 1662 562
tri 1662 560 1664 562 nw
tri 1730 560 1732 562 se
rect 1732 560 1740 562
rect 1652 554 1656 560
tri 1656 554 1662 560 nw
tri 1724 554 1730 560 se
rect 1730 554 1740 560
rect 1758 554 1760 562
rect 1768 554 1770 562
rect 1788 554 1790 562
rect 1798 554 1800 562
rect 1858 554 1860 562
rect 1868 554 1870 562
rect 1888 554 1890 562
rect 1898 554 1900 562
rect 1918 554 1920 562
rect 1928 554 1930 562
rect 1948 554 1950 562
rect 1958 554 1960 562
rect 1978 554 1980 562
rect 1988 554 1990 562
rect 1998 554 2000 562
tri 794 552 796 554 se
rect 796 552 814 554
rect 1072 552 1088 554
tri 1088 552 1090 554 nw
tri 1104 552 1106 554 se
rect 1106 552 1124 554
rect 1372 552 1390 554
tri 1390 552 1392 554 nw
tri 1406 552 1408 554 se
rect 1408 552 1424 554
rect 1432 552 1514 554
rect 1542 552 1654 554
tri 1654 552 1656 554 nw
tri 1722 552 1724 554 se
rect 1724 552 1740 554
rect 1748 552 1770 554
rect 1778 552 1800 554
rect 1838 552 1850 554
rect 1858 552 1880 554
rect 1888 552 1910 554
rect 1918 552 1940 554
rect 1948 552 1970 554
rect 1978 552 2000 554
tri 786 544 794 552 se
rect 794 544 804 552
rect 1072 544 1080 552
tri 1080 544 1088 552 nw
tri 1096 544 1104 552 se
rect 1104 544 1114 552
rect 1372 544 1382 552
tri 1382 544 1390 552 nw
tri 1398 544 1406 552 se
rect 1406 544 1414 552
rect 1432 544 1434 552
rect 1442 544 1444 552
rect 1452 544 1454 552
rect 1462 544 1464 552
rect 1472 544 1474 552
rect 1482 544 1484 552
rect 1492 544 1494 552
rect 1502 544 1504 552
rect 1542 544 1544 552
rect 1552 544 1554 552
rect 1562 544 1564 552
rect 1572 544 1574 552
rect 1582 544 1584 552
rect 1592 544 1594 552
rect 1602 544 1604 552
rect 1612 544 1614 552
rect 1622 544 1624 552
rect 1632 544 1634 552
rect 1642 544 1646 552
tri 1646 544 1654 552 nw
tri 1714 544 1722 552 se
rect 1722 544 1730 552
rect 1748 544 1750 552
rect 1758 544 1760 552
rect 1778 544 1780 552
rect 1788 544 1790 552
rect 1838 544 1840 552
rect 1848 544 1850 552
rect 1868 544 1870 552
rect 1878 544 1880 552
rect 1898 544 1900 552
rect 1908 544 1910 552
rect 1928 544 1930 552
rect 1938 544 1940 552
rect 1958 544 1960 552
rect 1968 544 1970 552
rect 1988 544 1990 552
rect 1998 544 2000 552
tri 784 542 786 544 se
rect 786 542 804 544
rect 1062 542 1078 544
tri 1078 542 1080 544 nw
tri 1094 542 1096 544 se
rect 1096 542 1114 544
rect 1362 542 1380 544
tri 1380 542 1382 544 nw
tri 1396 542 1398 544 se
rect 1398 542 1414 544
rect 1422 542 1504 544
rect 1532 542 1644 544
tri 1644 542 1646 544 nw
tri 1712 542 1714 544 se
rect 1714 542 1730 544
rect 1738 542 1760 544
rect 1768 542 1790 544
rect 1828 542 1850 544
rect 1858 542 1880 544
rect 1888 542 1910 544
rect 1918 542 1940 544
rect 1948 542 1970 544
rect 1978 542 2000 544
tri 776 534 784 542 se
rect 784 534 794 542
rect 1062 534 1070 542
tri 1070 534 1078 542 nw
tri 1086 534 1094 542 se
rect 1094 534 1104 542
rect 1362 534 1372 542
tri 1372 534 1380 542 nw
tri 1388 534 1396 542 se
rect 1396 534 1404 542
rect 1422 534 1424 542
rect 1432 534 1434 542
rect 1442 534 1444 542
rect 1452 534 1454 542
rect 1462 534 1464 542
rect 1472 534 1474 542
rect 1482 534 1484 542
rect 1492 534 1494 542
rect 1532 534 1534 542
rect 1542 534 1544 542
rect 1552 534 1554 542
rect 1562 534 1564 542
rect 1572 534 1574 542
rect 1582 534 1584 542
rect 1592 534 1594 542
rect 1602 534 1604 542
rect 1612 534 1614 542
rect 1622 534 1624 542
rect 1632 534 1636 542
tri 1636 534 1644 542 nw
tri 1704 534 1712 542 se
rect 1712 534 1720 542
rect 1738 534 1740 542
rect 1748 534 1750 542
rect 1768 534 1770 542
rect 1778 534 1780 542
rect 1828 534 1830 542
rect 1838 534 1840 542
rect 1858 534 1860 542
rect 1868 534 1870 542
rect 1888 534 1890 542
rect 1898 534 1900 542
rect 1918 534 1920 542
rect 1928 534 1930 542
rect 1948 534 1950 542
rect 1958 534 1960 542
rect 1978 534 1980 542
rect 1988 534 1990 542
rect 1998 534 2000 542
tri 774 532 776 534 se
rect 776 532 794 534
rect 1052 532 1068 534
tri 1068 532 1070 534 nw
tri 1084 532 1086 534 se
rect 1086 532 1104 534
rect 1352 532 1370 534
tri 1370 532 1372 534 nw
tri 1386 532 1388 534 se
rect 1388 532 1404 534
rect 1412 532 1494 534
rect 1522 532 1634 534
tri 1634 532 1636 534 nw
tri 1702 532 1704 534 se
rect 1704 532 1720 534
rect 1728 532 1750 534
rect 1758 532 1780 534
tri 766 524 774 532 se
rect 774 524 784 532
rect 1052 524 1060 532
tri 1060 524 1068 532 nw
tri 1076 524 1084 532 se
rect 1084 524 1094 532
rect 1352 524 1362 532
tri 1362 524 1370 532 nw
tri 1378 524 1386 532 se
rect 1386 524 1394 532
rect 1412 524 1414 532
rect 1422 524 1424 532
rect 1432 524 1434 532
rect 1442 524 1444 532
rect 1452 524 1454 532
rect 1462 524 1464 532
rect 1472 524 1474 532
rect 1482 524 1484 532
rect 1522 524 1524 532
rect 1532 524 1534 532
rect 1542 524 1544 532
rect 1552 524 1554 532
rect 1562 524 1564 532
rect 1572 524 1574 532
rect 1582 524 1584 532
rect 1592 524 1594 532
rect 1602 524 1604 532
rect 1612 524 1614 532
rect 1622 524 1626 532
tri 1626 524 1634 532 nw
tri 1694 524 1702 532 se
rect 1702 524 1710 532
rect 1728 524 1730 532
rect 1738 524 1740 532
rect 1758 524 1760 532
rect 1768 524 1770 532
rect 1808 531 1820 534
rect 1828 532 1850 534
rect 1858 532 1880 534
rect 1888 532 1910 534
rect 1918 532 1940 534
rect 1948 532 1970 534
rect 1978 532 2000 534
rect 1838 524 1840 532
rect 1848 524 1850 532
rect 1868 524 1870 532
rect 1878 524 1880 532
rect 1898 524 1900 532
rect 1908 524 1910 532
rect 1928 524 1930 532
rect 1938 524 1940 532
rect 1958 524 1960 532
rect 1968 524 1970 532
rect 1988 524 1990 532
rect 1998 524 2000 532
tri 765 523 766 524 se
rect 766 523 784 524
tri 764 522 765 523 se
rect 765 522 784 523
rect 1042 523 1059 524
tri 1059 523 1060 524 nw
tri 1075 523 1076 524 se
rect 1076 523 1094 524
rect 1042 522 1058 523
tri 1058 522 1059 523 nw
tri 1074 522 1075 523 se
rect 1075 522 1094 523
rect 1342 523 1361 524
tri 1361 523 1362 524 nw
tri 1377 523 1378 524 se
rect 1378 523 1394 524
rect 1342 522 1360 523
tri 1360 522 1361 523 nw
tri 1376 522 1377 523 se
rect 1377 522 1394 523
rect 1402 522 1484 524
rect 1512 523 1625 524
tri 1625 523 1626 524 nw
tri 1693 523 1694 524 se
rect 1694 523 1710 524
rect 1512 522 1624 523
tri 1624 522 1625 523 nw
tri 1692 522 1693 523 se
rect 1693 522 1710 523
rect 1718 522 1740 524
rect 1748 522 1770 524
rect 1808 522 1820 523
tri 756 514 764 522 se
rect 764 514 774 522
rect 1042 514 1050 522
tri 1050 514 1058 522 nw
tri 1066 514 1074 522 se
rect 1074 514 1084 522
rect 1342 514 1352 522
tri 1352 514 1360 522 nw
tri 1368 514 1376 522 se
rect 1376 514 1384 522
rect 1402 514 1404 522
rect 1412 514 1414 522
rect 1422 514 1424 522
rect 1432 514 1434 522
rect 1442 514 1444 522
rect 1452 514 1454 522
rect 1462 514 1464 522
rect 1472 514 1474 522
rect 1512 514 1514 522
rect 1522 514 1524 522
rect 1532 514 1534 522
rect 1542 514 1544 522
rect 1552 514 1554 522
rect 1562 514 1564 522
rect 1572 514 1574 522
rect 1582 514 1584 522
rect 1592 514 1594 522
rect 1602 514 1604 522
rect 1612 514 1616 522
tri 1616 514 1624 522 nw
tri 1684 514 1692 522 se
rect 1692 514 1700 522
rect 1718 514 1720 522
rect 1728 514 1730 522
rect 1748 514 1750 522
rect 1758 514 1760 522
rect 1808 514 1810 522
rect 1818 514 1820 522
tri 754 512 756 514 se
rect 756 512 774 514
rect 1032 512 1048 514
tri 1048 512 1050 514 nw
tri 1064 512 1066 514 se
rect 1066 512 1084 514
rect 1332 512 1350 514
tri 1350 512 1352 514 nw
tri 1366 512 1368 514 se
rect 1368 512 1384 514
rect 1392 512 1474 514
rect 1502 512 1614 514
tri 1614 512 1616 514 nw
tri 1682 512 1684 514 se
rect 1684 512 1700 514
rect 1708 512 1730 514
rect 1738 512 1760 514
rect 1798 512 1820 514
rect 1828 522 1850 524
rect 1858 522 1880 524
rect 1888 522 1910 524
rect 1918 522 1940 524
rect 1948 522 1970 524
rect 1978 522 2000 524
rect 1828 514 1830 522
rect 1838 514 1840 522
rect 1858 514 1860 522
rect 1868 514 1870 522
rect 1888 514 1890 522
rect 1898 514 1900 522
rect 1918 514 1920 522
rect 1928 514 1930 522
rect 1948 514 1950 522
rect 1958 514 1960 522
rect 1978 514 1980 522
rect 1988 514 1990 522
rect 1998 514 2000 522
rect 1828 512 1850 514
rect 1858 512 1880 514
rect 1888 512 1910 514
rect 1918 512 1940 514
rect 1948 512 1970 514
rect 1978 512 2000 514
tri 746 504 754 512 se
rect 754 504 764 512
rect 1032 504 1040 512
tri 1040 504 1048 512 nw
tri 1056 504 1064 512 se
rect 1064 504 1074 512
rect 1332 504 1342 512
tri 1342 504 1350 512 nw
tri 1358 504 1366 512 se
rect 1366 504 1374 512
rect 1392 504 1394 512
rect 1402 504 1404 512
rect 1412 504 1414 512
rect 1422 504 1424 512
rect 1432 504 1434 512
rect 1442 504 1444 512
rect 1452 504 1454 512
rect 1462 504 1464 512
rect 1502 504 1504 512
rect 1512 504 1514 512
rect 1522 504 1524 512
rect 1532 504 1534 512
rect 1542 504 1544 512
rect 1552 504 1554 512
rect 1562 504 1564 512
rect 1572 504 1574 512
rect 1582 504 1584 512
rect 1592 504 1594 512
rect 1602 504 1606 512
tri 1606 504 1614 512 nw
tri 1674 504 1682 512 se
rect 1682 504 1690 512
tri 744 502 746 504 se
rect 746 502 764 504
rect 1022 502 1038 504
tri 1038 502 1040 504 nw
tri 1054 502 1056 504 se
rect 1056 502 1074 504
rect 1322 502 1340 504
tri 1340 502 1342 504 nw
tri 1356 502 1358 504 se
rect 1358 502 1374 504
rect 1382 502 1464 504
rect 1492 502 1604 504
tri 1604 502 1606 504 nw
tri 1672 502 1674 504 se
rect 1674 502 1690 504
rect 1708 504 1710 512
rect 1718 504 1720 512
rect 1708 502 1720 504
rect 1738 504 1740 512
rect 1748 504 1750 512
rect 1738 502 1750 504
rect 1798 504 1800 512
rect 1808 504 1810 512
rect 1798 502 1810 504
rect 1838 504 1840 512
rect 1848 504 1850 512
rect 1838 502 1850 504
rect 1868 504 1870 512
rect 1878 504 1880 512
rect 1868 502 1880 504
rect 1898 504 1900 512
rect 1908 504 1910 512
rect 1898 502 1910 504
rect 1928 504 1930 512
rect 1938 504 1940 512
rect 1928 502 1940 504
rect 1958 504 1960 512
rect 1968 504 1970 512
rect 1958 502 1970 504
rect 1988 504 1990 512
rect 1998 504 2000 512
rect 1988 502 2000 504
tri 736 494 744 502 se
rect 744 494 754 502
rect 1022 494 1030 502
tri 1030 494 1038 502 nw
tri 1046 494 1054 502 se
rect 1054 494 1064 502
rect 1322 494 1332 502
tri 1332 494 1340 502 nw
tri 1348 494 1356 502 se
rect 1356 494 1364 502
rect 1382 494 1384 502
rect 1392 494 1394 502
rect 1402 494 1404 502
rect 1412 494 1414 502
rect 1422 494 1424 502
rect 1432 494 1434 502
rect 1442 494 1444 502
rect 1452 494 1454 502
rect 1492 494 1494 502
rect 1502 494 1504 502
rect 1512 494 1514 502
rect 1522 494 1524 502
rect 1532 494 1534 502
rect 1542 494 1544 502
rect 1552 494 1554 502
rect 1562 494 1564 502
rect 1572 494 1574 502
rect 1582 494 1584 502
rect 1592 494 1596 502
tri 1596 494 1604 502 nw
tri 1664 494 1672 502 se
rect 1672 494 1680 502
tri 734 492 736 494 se
rect 736 492 754 494
rect 1012 492 1028 494
tri 1028 492 1030 494 nw
tri 1044 492 1046 494 se
rect 1046 492 1064 494
rect 1312 492 1330 494
tri 1330 492 1332 494 nw
tri 1346 492 1348 494 se
rect 1348 492 1364 494
rect 1372 492 1454 494
rect 1482 492 1594 494
tri 1594 492 1596 494 nw
tri 1662 492 1664 494 se
rect 1664 492 1690 494
tri 726 484 734 492 se
rect 734 484 744 492
rect 1012 484 1020 492
tri 1020 484 1028 492 nw
tri 1036 484 1044 492 se
rect 1044 484 1054 492
rect 1312 484 1322 492
tri 1322 484 1330 492 nw
tri 1338 484 1346 492 se
rect 1346 484 1354 492
rect 1372 484 1374 492
rect 1382 484 1384 492
rect 1392 484 1394 492
rect 1402 484 1404 492
rect 1412 484 1414 492
rect 1422 484 1424 492
rect 1432 484 1434 492
rect 1442 484 1444 492
rect 1482 484 1484 492
rect 1492 484 1494 492
rect 1502 484 1504 492
rect 1512 484 1514 492
rect 1522 484 1524 492
rect 1532 484 1534 492
rect 1542 484 1544 492
rect 1552 484 1554 492
rect 1562 484 1564 492
rect 1572 484 1574 492
rect 1582 484 1586 492
tri 1586 484 1594 492 nw
tri 1654 484 1662 492 se
rect 1662 484 1670 492
rect 1678 484 1680 492
rect 1688 484 1690 492
rect 1698 492 1710 494
rect 1698 484 1700 492
rect 1708 484 1710 492
rect 1718 492 1730 494
rect 1718 484 1720 492
rect 1728 484 1730 492
rect 1738 492 1750 494
rect 1738 484 1740 492
rect 1748 484 1750 492
rect 1788 492 1800 494
rect 1788 484 1790 492
rect 1798 484 1800 492
rect 1808 492 1820 494
rect 1808 484 1810 492
rect 1818 484 1820 492
rect 1828 492 1840 494
rect 1828 484 1830 492
rect 1838 484 1840 492
rect 1848 492 1860 494
rect 1848 484 1850 492
rect 1858 484 1860 492
rect 1868 492 1890 494
rect 1868 484 1870 492
rect 1878 484 1890 492
tri 724 482 726 484 se
rect 726 482 744 484
rect 1002 482 1018 484
tri 1018 482 1020 484 nw
tri 1034 482 1036 484 se
rect 1036 482 1054 484
rect 1302 482 1320 484
tri 1320 482 1322 484 nw
tri 1336 482 1338 484 se
rect 1338 482 1354 484
rect 1362 482 1444 484
rect 1472 482 1584 484
tri 1584 482 1586 484 nw
tri 1652 482 1654 484 se
rect 1654 482 1750 484
rect 1778 482 1890 484
tri 716 474 724 482 se
rect 724 474 734 482
rect 1002 474 1010 482
tri 1010 474 1018 482 nw
tri 1026 474 1034 482 se
rect 1034 474 1044 482
rect 1302 474 1312 482
tri 1312 474 1320 482 nw
tri 1328 474 1336 482 se
rect 1336 474 1344 482
rect 1362 474 1364 482
rect 1372 474 1374 482
rect 1382 474 1384 482
rect 1392 474 1394 482
rect 1402 474 1404 482
rect 1412 474 1414 482
rect 1422 474 1424 482
rect 1432 474 1434 482
rect 1472 474 1474 482
rect 1482 474 1484 482
rect 1492 474 1494 482
rect 1502 474 1504 482
rect 1512 474 1514 482
rect 1522 474 1524 482
rect 1532 474 1534 482
rect 1542 474 1544 482
rect 1552 474 1554 482
rect 1562 474 1564 482
rect 1572 474 1576 482
tri 1576 474 1584 482 nw
tri 1644 474 1652 482 se
rect 1652 474 1660 482
rect 1668 474 1670 482
rect 1678 474 1680 482
rect 1688 474 1690 482
rect 1698 474 1700 482
rect 1708 474 1710 482
rect 1718 474 1720 482
rect 1728 474 1730 482
rect 1738 474 1740 482
rect 1778 474 1780 482
rect 1788 474 1790 482
rect 1798 474 1800 482
rect 1808 474 1810 482
rect 1818 474 1820 482
rect 1828 474 1830 482
rect 1838 474 1840 482
rect 1848 474 1850 482
rect 1858 474 1860 482
rect 1868 474 1880 482
tri 714 472 716 474 se
rect 716 472 734 474
rect 992 472 1008 474
tri 1008 472 1010 474 nw
tri 1024 472 1026 474 se
rect 1026 472 1044 474
rect 1292 472 1310 474
tri 1310 472 1312 474 nw
tri 1326 472 1328 474 se
rect 1328 472 1344 474
rect 1352 472 1434 474
rect 1462 472 1574 474
tri 1574 472 1576 474 nw
tri 1642 472 1644 474 se
rect 1644 472 1740 474
rect 1768 472 1880 474
tri 706 464 714 472 se
rect 714 464 724 472
rect 992 464 1000 472
tri 1000 464 1008 472 nw
tri 1016 464 1024 472 se
rect 1024 464 1034 472
rect 1292 464 1302 472
tri 1302 464 1310 472 nw
tri 1318 464 1326 472 se
rect 1326 464 1334 472
rect 1352 464 1354 472
rect 1362 464 1364 472
rect 1372 464 1374 472
rect 1382 464 1384 472
rect 1392 464 1394 472
rect 1402 464 1404 472
rect 1412 464 1414 472
rect 1422 464 1424 472
rect 1462 464 1464 472
rect 1472 464 1474 472
rect 1482 464 1484 472
rect 1492 464 1494 472
rect 1502 464 1504 472
rect 1512 464 1514 472
rect 1522 464 1524 472
rect 1532 464 1534 472
rect 1542 464 1544 472
rect 1552 464 1554 472
rect 1562 464 1566 472
tri 1566 464 1574 472 nw
tri 1634 464 1642 472 se
rect 1642 464 1650 472
rect 1658 464 1660 472
rect 1668 464 1670 472
rect 1678 464 1680 472
rect 1688 464 1690 472
rect 1698 464 1700 472
rect 1708 464 1710 472
rect 1718 464 1720 472
rect 1728 464 1730 472
rect 1768 464 1770 472
rect 1778 464 1780 472
rect 1788 464 1790 472
rect 1798 464 1800 472
rect 1808 464 1810 472
rect 1818 464 1820 472
rect 1828 464 1830 472
rect 1838 464 1840 472
rect 1848 464 1850 472
rect 1858 464 1870 472
tri 704 462 706 464 se
rect 706 462 724 464
rect 982 462 998 464
tri 998 462 1000 464 nw
tri 1014 462 1016 464 se
rect 1016 462 1034 464
rect 1282 462 1300 464
tri 1300 462 1302 464 nw
tri 1316 462 1318 464 se
rect 1318 462 1334 464
rect 1342 462 1424 464
rect 1452 462 1564 464
tri 1564 462 1566 464 nw
tri 1632 462 1634 464 se
rect 1634 462 1730 464
rect 1758 462 1870 464
tri 696 454 704 462 se
rect 704 454 714 462
rect 982 454 990 462
tri 990 454 998 462 nw
tri 1006 454 1014 462 se
rect 1014 454 1024 462
rect 1282 454 1292 462
tri 1292 454 1300 462 nw
tri 1308 454 1316 462 se
rect 1316 454 1324 462
rect 1342 454 1344 462
rect 1352 454 1354 462
rect 1362 454 1364 462
rect 1372 454 1374 462
rect 1382 454 1384 462
rect 1392 454 1394 462
rect 1402 454 1404 462
rect 1412 454 1414 462
rect 1452 454 1454 462
rect 1462 454 1464 462
rect 1472 454 1474 462
rect 1482 454 1484 462
rect 1492 454 1494 462
rect 1502 454 1504 462
rect 1512 454 1514 462
rect 1522 454 1524 462
rect 1532 454 1534 462
rect 1542 454 1544 462
rect 1552 454 1556 462
tri 1556 454 1564 462 nw
tri 1624 454 1632 462 se
rect 1632 454 1640 462
rect 1648 454 1650 462
rect 1658 454 1660 462
rect 1668 454 1670 462
rect 1678 454 1680 462
rect 1688 454 1690 462
rect 1698 454 1700 462
rect 1708 454 1710 462
rect 1718 454 1720 462
rect 1758 454 1760 462
rect 1768 454 1770 462
rect 1778 454 1780 462
rect 1788 454 1790 462
rect 1798 454 1800 462
rect 1808 454 1810 462
rect 1818 454 1820 462
rect 1828 454 1830 462
rect 1838 454 1840 462
rect 1848 454 1860 462
tri 694 452 696 454 se
rect 696 452 714 454
rect 972 452 988 454
tri 988 452 990 454 nw
tri 1004 452 1006 454 se
rect 1006 452 1024 454
rect 1272 452 1290 454
tri 1290 452 1292 454 nw
tri 1306 452 1308 454 se
rect 1308 452 1324 454
rect 1332 452 1414 454
rect 1442 452 1554 454
tri 1554 452 1556 454 nw
tri 1622 452 1624 454 se
rect 1624 452 1720 454
rect 1748 452 1860 454
tri 686 444 694 452 se
rect 694 444 704 452
rect 972 444 980 452
tri 980 444 988 452 nw
tri 996 444 1004 452 se
rect 1004 444 1014 452
rect 1272 444 1282 452
tri 1282 444 1290 452 nw
tri 1298 444 1306 452 se
rect 1306 444 1314 452
rect 1332 444 1334 452
rect 1342 444 1344 452
rect 1352 444 1354 452
rect 1362 444 1364 452
rect 1372 444 1374 452
rect 1382 444 1384 452
rect 1392 444 1394 452
rect 1402 444 1404 452
rect 1442 444 1444 452
rect 1452 444 1454 452
rect 1462 444 1464 452
rect 1472 444 1474 452
rect 1482 444 1484 452
rect 1492 444 1494 452
rect 1502 444 1504 452
rect 1512 444 1514 452
rect 1522 444 1524 452
rect 1532 444 1534 452
rect 1542 444 1546 452
tri 1546 444 1554 452 nw
tri 1614 444 1622 452 se
rect 1622 444 1630 452
rect 1638 444 1640 452
rect 1648 444 1650 452
rect 1658 444 1660 452
rect 1668 444 1670 452
rect 1678 444 1680 452
rect 1688 444 1690 452
rect 1698 444 1700 452
rect 1708 444 1710 452
rect 1748 444 1750 452
rect 1758 444 1760 452
rect 1768 444 1770 452
rect 1778 444 1780 452
rect 1788 444 1790 452
rect 1798 444 1800 452
rect 1808 444 1810 452
rect 1818 444 1820 452
rect 1828 444 1830 452
rect 1838 444 1850 452
tri 684 442 686 444 se
rect 686 442 704 444
rect 962 442 978 444
tri 978 442 980 444 nw
tri 994 442 996 444 se
rect 996 442 1014 444
rect 1262 442 1280 444
tri 1280 442 1282 444 nw
tri 1296 442 1298 444 se
rect 1298 442 1314 444
rect 1322 442 1404 444
rect 1432 442 1544 444
tri 1544 442 1546 444 nw
tri 1612 442 1614 444 se
rect 1614 442 1710 444
rect 1738 442 1850 444
tri 676 434 684 442 se
rect 684 434 694 442
rect 962 434 970 442
tri 970 434 978 442 nw
tri 986 434 994 442 se
rect 994 434 1004 442
rect 1262 434 1272 442
tri 1272 434 1280 442 nw
tri 1288 434 1296 442 se
rect 1296 434 1304 442
rect 1322 434 1324 442
rect 1332 434 1334 442
rect 1342 434 1344 442
rect 1352 434 1354 442
rect 1362 434 1364 442
rect 1372 434 1374 442
rect 1382 434 1384 442
rect 1392 434 1394 442
rect 1432 434 1434 442
rect 1442 434 1444 442
rect 1452 434 1454 442
rect 1462 434 1464 442
rect 1472 434 1474 442
rect 1482 434 1484 442
rect 1492 434 1494 442
rect 1502 434 1504 442
rect 1512 434 1514 442
rect 1522 434 1524 442
rect 1532 434 1536 442
tri 1536 434 1544 442 nw
tri 1604 434 1612 442 se
rect 1612 434 1620 442
rect 1628 434 1630 442
rect 1638 434 1640 442
rect 1648 434 1650 442
rect 1658 434 1660 442
rect 1668 434 1670 442
rect 1678 434 1680 442
rect 1688 434 1690 442
rect 1698 434 1700 442
rect 1738 434 1740 442
rect 1748 434 1750 442
rect 1758 434 1760 442
rect 1768 434 1770 442
rect 1778 434 1780 442
rect 1788 434 1790 442
rect 1798 434 1800 442
rect 1808 434 1810 442
rect 1818 434 1820 442
rect 1828 434 1840 442
tri 674 432 676 434 se
rect 676 432 694 434
rect 952 432 968 434
tri 968 432 970 434 nw
tri 984 432 986 434 se
rect 986 432 1004 434
rect 1252 432 1270 434
tri 1270 432 1272 434 nw
tri 1286 432 1288 434 se
rect 1288 432 1304 434
rect 1312 432 1394 434
rect 1422 432 1534 434
tri 1534 432 1536 434 nw
tri 1602 432 1604 434 se
rect 1604 432 1700 434
rect 1728 432 1840 434
tri 666 424 674 432 se
rect 674 424 684 432
rect 952 424 960 432
tri 960 424 968 432 nw
tri 976 424 984 432 se
rect 984 424 994 432
rect 1252 424 1262 432
tri 1262 424 1270 432 nw
tri 1278 424 1286 432 se
rect 1286 424 1294 432
rect 1312 424 1314 432
rect 1322 424 1324 432
rect 1332 424 1334 432
rect 1342 424 1344 432
rect 1352 424 1354 432
rect 1362 424 1364 432
rect 1372 424 1374 432
rect 1382 424 1384 432
rect 1422 424 1424 432
rect 1432 424 1434 432
rect 1442 424 1444 432
rect 1452 424 1454 432
rect 1462 424 1464 432
rect 1472 424 1474 432
rect 1482 424 1484 432
rect 1492 424 1494 432
rect 1502 424 1504 432
rect 1512 424 1514 432
rect 1522 424 1526 432
tri 1526 424 1534 432 nw
tri 1594 424 1602 432 se
rect 1602 424 1610 432
rect 1618 424 1620 432
rect 1628 424 1630 432
rect 1638 424 1640 432
rect 1648 424 1650 432
rect 1658 424 1660 432
rect 1668 424 1670 432
rect 1678 424 1680 432
rect 1688 424 1690 432
rect 1728 424 1730 432
rect 1738 424 1740 432
rect 1748 424 1750 432
rect 1758 424 1760 432
rect 1768 424 1770 432
rect 1778 424 1780 432
rect 1788 424 1790 432
rect 1798 424 1800 432
rect 1808 424 1810 432
rect 1818 424 1830 432
tri 664 422 666 424 se
rect 666 422 684 424
rect 942 422 958 424
tri 958 422 960 424 nw
tri 974 422 976 424 se
rect 976 422 994 424
rect 1242 422 1260 424
tri 1260 422 1262 424 nw
tri 1276 422 1278 424 se
rect 1278 422 1294 424
rect 1302 422 1384 424
rect 1412 422 1524 424
tri 1524 422 1526 424 nw
tri 1592 422 1594 424 se
rect 1594 422 1690 424
rect 1718 422 1830 424
tri 662 420 664 422 se
rect 664 420 674 422
rect 662 412 674 420
rect 942 420 956 422
tri 956 420 958 422 nw
tri 972 420 974 422 se
rect 974 420 984 422
rect 942 414 950 420
tri 950 414 956 420 nw
tri 966 414 972 420 se
rect 972 414 984 420
rect 1242 414 1252 422
tri 1252 414 1260 422 nw
tri 1268 414 1276 422 se
rect 1276 414 1284 422
rect 1302 414 1304 422
rect 1312 414 1314 422
rect 1322 414 1324 422
rect 1332 414 1334 422
rect 1342 414 1344 422
rect 1352 414 1354 422
rect 1362 414 1364 422
rect 1372 414 1374 422
rect 1412 414 1414 422
rect 1422 414 1424 422
rect 1432 414 1434 422
rect 1442 414 1444 422
rect 1452 414 1454 422
rect 1462 414 1464 422
rect 1472 414 1474 422
rect 1482 414 1484 422
rect 1492 414 1494 422
rect 1502 414 1504 422
rect 1512 416 1518 422
tri 1518 416 1524 422 nw
tri 1586 416 1592 422 se
rect 1592 416 1600 422
rect 1512 414 1516 416
tri 1516 414 1518 416 nw
tri 1584 414 1586 416 se
rect 1586 414 1600 416
rect 1608 414 1610 422
rect 1618 414 1620 422
rect 1628 414 1630 422
rect 1638 414 1640 422
rect 1648 414 1650 422
rect 1658 414 1660 422
rect 1668 414 1670 422
rect 1678 414 1680 422
rect 1718 414 1720 422
rect 1728 414 1730 422
rect 1738 414 1740 422
rect 1748 414 1750 422
rect 1758 414 1760 422
rect 1768 414 1770 422
rect 1778 414 1780 422
rect 1788 414 1790 422
rect 1798 414 1800 422
rect 1808 415 1830 422
rect 1808 414 1822 415
tri 1822 414 1823 415 nw
tri 1823 414 1824 415 ne
rect 1824 414 1830 415
rect 932 412 948 414
tri 948 412 950 414 nw
tri 964 412 966 414 se
rect 966 412 984 414
rect 1232 412 1250 414
tri 1250 412 1252 414 nw
tri 1266 412 1268 414 se
rect 1268 412 1284 414
rect 1292 412 1374 414
rect 1402 412 1514 414
tri 1514 412 1516 414 nw
tri 1582 412 1584 414 se
rect 1584 412 1680 414
rect 1708 412 1820 414
tri 1820 412 1822 414 nw
tri 1824 412 1826 414 ne
rect 1826 412 1840 414
rect 662 4 664 412
rect 932 404 940 412
tri 940 404 948 412 nw
tri 956 404 964 412 se
rect 964 404 974 412
rect 1232 404 1242 412
tri 1242 404 1250 412 nw
tri 1258 404 1266 412 se
rect 1266 404 1274 412
rect 1292 404 1294 412
rect 1302 404 1304 412
rect 1312 404 1314 412
rect 1322 404 1324 412
rect 1332 404 1334 412
rect 1342 404 1344 412
rect 1352 404 1354 412
rect 1362 404 1364 412
rect 1402 404 1404 412
rect 1412 404 1414 412
rect 1422 404 1424 412
rect 1432 404 1434 412
rect 1442 404 1444 412
rect 1452 404 1454 412
rect 1462 404 1464 412
rect 1472 404 1474 412
rect 1482 404 1484 412
rect 1492 404 1494 412
rect 1502 404 1506 412
tri 1506 404 1514 412 nw
tri 1574 404 1582 412 se
rect 1582 404 1590 412
rect 1598 404 1600 412
rect 1608 404 1610 412
rect 1618 404 1620 412
rect 1628 404 1630 412
rect 1638 404 1640 412
rect 1648 404 1650 412
rect 1658 404 1660 412
rect 1668 404 1670 412
rect 1708 404 1710 412
rect 1718 404 1720 412
rect 1728 404 1730 412
rect 1738 404 1740 412
rect 1748 404 1750 412
rect 1758 404 1760 412
rect 1768 404 1770 412
rect 1778 404 1780 412
rect 1788 404 1790 412
rect 1798 407 1815 412
tri 1815 407 1820 412 nw
tri 1826 407 1831 412 ne
rect 1798 404 1812 407
tri 1812 404 1815 407 nw
tri 1828 404 1831 407 se
rect 1831 404 1840 412
rect 932 402 938 404
tri 938 402 940 404 nw
tri 954 402 956 404 se
rect 956 402 974 404
rect 1222 402 1240 404
tri 1240 402 1242 404 nw
tri 1256 402 1258 404 se
rect 1258 402 1274 404
rect 1282 402 1364 404
rect 1392 402 1504 404
tri 1504 402 1506 404 nw
tri 1572 402 1574 404 se
rect 1574 402 1670 404
rect 1698 402 1810 404
tri 1810 402 1812 404 nw
tri 1826 402 1828 404 se
rect 1828 402 1840 404
rect 932 394 933 402
tri 933 397 938 402 nw
tri 949 397 954 402 se
rect 954 397 964 402
tri 933 394 936 397 sw
tri 946 394 949 397 se
rect 949 394 964 397
rect 1222 394 1232 402
tri 1232 394 1240 402 nw
tri 1250 396 1256 402 se
rect 1256 396 1264 402
tri 1248 394 1250 396 se
rect 1250 394 1264 396
rect 1282 394 1284 402
rect 1292 394 1294 402
rect 1302 394 1304 402
rect 1312 394 1314 402
rect 1322 394 1324 402
rect 1332 394 1334 402
rect 1342 394 1344 402
rect 1352 394 1354 402
rect 1392 394 1394 402
rect 1402 394 1404 402
rect 1412 394 1414 402
rect 1422 394 1424 402
rect 1432 394 1434 402
rect 1442 394 1444 402
rect 1452 394 1454 402
rect 1462 394 1464 402
rect 1472 394 1474 402
rect 1482 394 1484 402
rect 1492 396 1498 402
tri 1498 396 1504 402 nw
tri 1566 396 1572 402 se
rect 1572 396 1580 402
rect 1492 394 1496 396
tri 1496 394 1498 396 nw
tri 1564 394 1566 396 se
rect 1566 394 1580 396
rect 1588 394 1590 402
rect 1598 394 1600 402
rect 1608 394 1610 402
rect 1618 394 1620 402
rect 1628 394 1630 402
rect 1638 394 1640 402
rect 1648 394 1650 402
rect 1658 394 1660 402
rect 1698 394 1700 402
rect 1708 394 1710 402
rect 1718 394 1720 402
rect 1728 394 1730 402
rect 1738 394 1740 402
rect 1748 394 1750 402
rect 1758 394 1760 402
rect 1768 394 1770 402
rect 1778 394 1780 402
rect 1788 394 1802 402
tri 1802 394 1810 402 nw
tri 1818 394 1826 402 se
rect 1826 394 1830 402
rect 932 392 936 394
tri 936 392 938 394 sw
tri 944 392 946 394 se
rect 946 392 964 394
rect 1212 392 1230 394
tri 1230 392 1232 394 nw
tri 1246 392 1248 394 se
rect 1248 392 1264 394
rect 1272 392 1354 394
rect 1382 392 1494 394
tri 1494 392 1496 394 nw
tri 1562 392 1564 394 se
rect 1564 392 1660 394
rect 1688 392 1800 394
tri 1800 392 1802 394 nw
tri 1816 392 1818 394 se
rect 1818 392 1830 394
rect 932 389 938 392
tri 938 389 941 392 sw
tri 941 389 944 392 se
rect 944 389 954 392
rect 932 382 954 389
rect 1212 388 1226 392
tri 1226 388 1230 392 nw
tri 1242 388 1246 392 se
rect 1246 388 1254 392
rect 1212 384 1222 388
tri 1222 384 1226 388 nw
tri 1238 384 1242 388 se
rect 1242 384 1254 388
rect 1272 384 1274 392
rect 1282 384 1284 392
rect 1292 384 1294 392
rect 1302 384 1304 392
rect 1312 384 1314 392
rect 1322 384 1324 392
rect 1332 384 1334 392
rect 1342 384 1344 392
rect 1382 384 1384 392
rect 1392 384 1394 392
rect 1402 384 1404 392
rect 1412 384 1414 392
rect 1422 384 1424 392
rect 1432 384 1434 392
rect 1442 384 1444 392
rect 1452 384 1454 392
rect 1462 384 1464 392
rect 1472 384 1474 392
rect 1482 384 1486 392
tri 1486 384 1494 392 nw
tri 1554 384 1562 392 se
rect 1562 384 1570 392
rect 1578 384 1580 392
rect 1588 384 1590 392
rect 1598 384 1600 392
rect 1608 384 1610 392
rect 1618 384 1620 392
rect 1628 384 1630 392
rect 1638 384 1640 392
rect 1648 384 1650 392
rect 1688 384 1690 392
rect 1698 384 1700 392
rect 1708 384 1710 392
rect 1718 384 1720 392
rect 1728 384 1730 392
rect 1738 384 1740 392
rect 1748 384 1750 392
rect 1758 384 1760 392
rect 1768 384 1770 392
rect 1778 384 1792 392
tri 1792 384 1800 392 nw
tri 1808 384 1816 392 se
rect 1816 384 1820 392
rect 1202 382 1220 384
tri 1220 382 1222 384 nw
tri 1236 382 1238 384 se
rect 1238 382 1254 384
rect 1262 382 1344 384
rect 1372 382 1484 384
tri 1484 382 1486 384 nw
tri 1552 382 1554 384 se
rect 1554 382 1650 384
rect 1678 382 1790 384
tri 1790 382 1792 384 nw
tri 1806 382 1808 384 se
rect 1808 382 1820 384
rect 1202 374 1212 382
tri 1212 374 1220 382 nw
tri 1228 374 1236 382 se
rect 1236 374 1244 382
rect 1262 374 1264 382
rect 1272 374 1274 382
rect 1282 374 1284 382
rect 1292 374 1294 382
rect 1302 374 1304 382
rect 1312 374 1314 382
rect 1322 374 1324 382
rect 1332 374 1334 382
rect 1372 374 1374 382
rect 1382 374 1384 382
rect 1392 374 1394 382
rect 1402 374 1404 382
rect 1412 374 1414 382
rect 1422 374 1424 382
rect 1432 374 1434 382
rect 1442 374 1444 382
rect 1452 374 1454 382
rect 1462 374 1464 382
rect 1472 374 1476 382
tri 1476 374 1484 382 nw
tri 1544 374 1552 382 se
rect 1552 374 1560 382
rect 1568 374 1570 382
rect 1578 374 1580 382
rect 1588 374 1590 382
rect 1598 374 1600 382
rect 1608 374 1610 382
rect 1618 374 1620 382
rect 1628 374 1630 382
rect 1638 374 1640 382
rect 1678 374 1680 382
rect 1688 374 1690 382
rect 1698 374 1700 382
rect 1708 374 1710 382
rect 1718 374 1720 382
rect 1728 374 1730 382
rect 1738 374 1740 382
rect 1748 374 1750 382
rect 1758 374 1760 382
rect 1768 374 1782 382
tri 1782 374 1790 382 nw
tri 1798 374 1806 382 se
rect 1806 374 1810 382
rect 1192 372 1210 374
tri 1210 372 1212 374 nw
tri 1226 372 1228 374 se
rect 1228 372 1244 374
rect 1252 372 1334 374
rect 1362 372 1474 374
tri 1474 372 1476 374 nw
tri 1542 372 1544 374 se
rect 1544 372 1640 374
rect 1668 372 1780 374
tri 1780 372 1782 374 nw
tri 1796 372 1798 374 se
rect 1798 372 1810 374
rect 1192 364 1202 372
tri 1202 364 1210 372 nw
tri 1218 364 1226 372 se
rect 1226 364 1234 372
rect 1252 364 1254 372
rect 1262 364 1264 372
rect 1272 364 1274 372
rect 1282 364 1284 372
rect 1292 364 1294 372
rect 1302 364 1304 372
rect 1312 364 1314 372
rect 1322 364 1324 372
rect 1362 364 1364 372
rect 1372 364 1374 372
rect 1382 364 1384 372
rect 1392 364 1394 372
rect 1402 364 1404 372
rect 1412 364 1414 372
rect 1422 364 1424 372
rect 1432 364 1434 372
rect 1442 364 1444 372
rect 1452 364 1454 372
rect 1462 364 1466 372
tri 1466 364 1474 372 nw
tri 1534 364 1542 372 se
rect 1542 364 1550 372
rect 1558 364 1560 372
rect 1568 364 1570 372
rect 1578 364 1580 372
rect 1588 364 1590 372
rect 1598 364 1600 372
rect 1608 364 1610 372
rect 1618 364 1620 372
rect 1628 364 1630 372
rect 1668 364 1670 372
rect 1678 364 1680 372
rect 1688 364 1690 372
rect 1698 364 1700 372
rect 1708 364 1710 372
rect 1718 364 1720 372
rect 1728 364 1730 372
rect 1738 364 1740 372
rect 1748 364 1750 372
rect 1758 364 1772 372
tri 1772 364 1780 372 nw
tri 1788 364 1796 372 se
rect 1796 364 1800 372
rect 1182 362 1200 364
tri 1200 362 1202 364 nw
tri 1216 362 1218 364 se
rect 1218 362 1234 364
rect 1242 362 1324 364
rect 1352 362 1464 364
tri 1464 362 1466 364 nw
tri 1532 362 1534 364 se
rect 1534 362 1630 364
rect 1658 362 1770 364
tri 1770 362 1772 364 nw
tri 1786 362 1788 364 se
rect 1788 362 1800 364
rect 1182 354 1192 362
tri 1192 354 1200 362 nw
tri 1208 354 1216 362 se
rect 1216 354 1224 362
rect 1242 354 1244 362
rect 1252 354 1254 362
rect 1262 354 1264 362
rect 1272 354 1274 362
rect 1282 354 1284 362
rect 1292 354 1294 362
rect 1302 354 1304 362
rect 1312 354 1314 362
rect 1352 354 1354 362
rect 1362 354 1364 362
rect 1372 354 1374 362
rect 1382 354 1384 362
rect 1392 354 1394 362
rect 1402 354 1404 362
rect 1412 354 1414 362
rect 1422 354 1424 362
rect 1432 354 1434 362
rect 1442 354 1444 362
rect 1452 354 1456 362
tri 1456 354 1464 362 nw
tri 1524 354 1532 362 se
rect 1532 354 1540 362
rect 1548 354 1550 362
rect 1558 354 1560 362
rect 1568 354 1570 362
rect 1578 354 1580 362
rect 1588 354 1590 362
rect 1598 354 1600 362
rect 1608 354 1610 362
rect 1618 354 1620 362
rect 1658 354 1660 362
rect 1668 354 1670 362
rect 1678 354 1680 362
rect 1688 354 1690 362
rect 1698 354 1700 362
rect 1708 354 1710 362
rect 1718 354 1720 362
rect 1728 354 1730 362
rect 1738 354 1740 362
rect 1748 354 1762 362
tri 1762 354 1770 362 nw
tri 1778 354 1786 362 se
rect 1786 354 1790 362
rect 1172 352 1190 354
tri 1190 352 1192 354 nw
tri 1206 352 1208 354 se
rect 1208 352 1224 354
rect 1232 352 1314 354
rect 1342 352 1454 354
tri 1454 352 1456 354 nw
tri 1522 352 1524 354 se
rect 1524 352 1620 354
rect 1648 352 1760 354
tri 1760 352 1762 354 nw
tri 1776 352 1778 354 se
rect 1778 352 1790 354
rect 1172 344 1182 352
tri 1182 344 1190 352 nw
tri 1198 344 1206 352 se
rect 1206 344 1214 352
rect 1232 344 1234 352
rect 1242 344 1244 352
rect 1252 344 1254 352
rect 1262 344 1264 352
rect 1272 344 1274 352
rect 1282 344 1284 352
rect 1292 344 1294 352
rect 1302 344 1304 352
rect 1342 344 1344 352
rect 1352 344 1354 352
rect 1362 344 1364 352
rect 1372 344 1374 352
rect 1382 344 1384 352
rect 1392 344 1394 352
rect 1402 344 1404 352
rect 1412 344 1414 352
rect 1422 344 1424 352
rect 1432 344 1434 352
rect 1442 344 1446 352
tri 1446 344 1454 352 nw
tri 1514 344 1522 352 se
rect 1522 344 1530 352
rect 1538 344 1540 352
rect 1548 344 1550 352
rect 1558 344 1560 352
rect 1568 344 1570 352
rect 1578 344 1580 352
rect 1588 344 1590 352
rect 1598 344 1600 352
rect 1608 344 1610 352
rect 1648 344 1650 352
rect 1658 344 1660 352
rect 1668 344 1670 352
rect 1678 344 1680 352
rect 1688 344 1690 352
rect 1698 344 1700 352
rect 1708 344 1710 352
rect 1718 344 1720 352
rect 1728 344 1730 352
rect 1738 344 1752 352
tri 1752 344 1760 352 nw
tri 1768 344 1776 352 se
rect 1776 344 1780 352
rect 1162 342 1180 344
tri 1180 342 1182 344 nw
tri 1196 342 1198 344 se
rect 1198 342 1214 344
rect 1222 342 1304 344
rect 1332 342 1444 344
tri 1444 342 1446 344 nw
tri 1512 342 1514 344 se
rect 1514 342 1610 344
rect 1638 342 1750 344
tri 1750 342 1752 344 nw
tri 1766 342 1768 344 se
rect 1768 342 1780 344
rect 1162 334 1172 342
tri 1172 334 1180 342 nw
tri 1188 334 1196 342 se
rect 1196 334 1204 342
rect 1222 334 1224 342
rect 1232 334 1234 342
rect 1242 334 1244 342
rect 1252 334 1254 342
rect 1262 334 1264 342
rect 1272 334 1274 342
rect 1282 334 1284 342
rect 1292 334 1294 342
rect 1332 334 1334 342
rect 1342 334 1344 342
rect 1352 334 1354 342
rect 1362 334 1364 342
rect 1372 334 1374 342
rect 1382 334 1384 342
rect 1392 334 1394 342
rect 1402 334 1404 342
rect 1412 334 1414 342
rect 1422 334 1424 342
rect 1432 334 1436 342
tri 1436 334 1444 342 nw
tri 1504 334 1512 342 se
rect 1512 334 1520 342
rect 1528 334 1530 342
rect 1538 334 1540 342
rect 1548 334 1550 342
rect 1558 334 1560 342
rect 1568 334 1570 342
rect 1578 334 1580 342
rect 1588 334 1590 342
rect 1598 334 1600 342
rect 1638 334 1640 342
rect 1648 334 1650 342
rect 1658 334 1660 342
rect 1668 334 1670 342
rect 1678 334 1680 342
rect 1688 334 1690 342
rect 1698 334 1700 342
rect 1708 334 1710 342
rect 1718 334 1720 342
rect 1728 334 1742 342
tri 1742 334 1750 342 nw
tri 1758 334 1766 342 se
rect 1766 334 1770 342
rect 1152 332 1170 334
tri 1170 332 1172 334 nw
tri 1186 332 1188 334 se
rect 1188 332 1204 334
rect 1212 332 1294 334
rect 1322 332 1434 334
tri 1434 332 1436 334 nw
tri 1502 332 1504 334 se
rect 1504 332 1600 334
rect 1628 332 1740 334
tri 1740 332 1742 334 nw
tri 1756 332 1758 334 se
rect 1758 332 1770 334
rect 1152 324 1162 332
tri 1162 324 1170 332 nw
tri 1178 324 1186 332 se
rect 1186 324 1194 332
rect 1212 324 1214 332
rect 1222 324 1224 332
rect 1232 324 1234 332
rect 1242 324 1244 332
rect 1252 324 1254 332
rect 1262 324 1264 332
rect 1272 324 1274 332
rect 1282 324 1284 332
rect 1322 324 1324 332
rect 1332 324 1334 332
rect 1342 324 1344 332
rect 1352 324 1354 332
rect 1362 324 1364 332
rect 1372 324 1374 332
rect 1382 324 1384 332
rect 1392 324 1394 332
rect 1402 324 1404 332
rect 1412 324 1414 332
rect 1422 328 1430 332
tri 1430 328 1434 332 nw
tri 1498 328 1502 332 se
rect 1502 328 1510 332
rect 1422 324 1426 328
tri 1426 324 1430 328 nw
tri 1494 324 1498 328 se
rect 1498 324 1510 328
rect 1518 324 1520 332
rect 1528 324 1530 332
rect 1538 324 1540 332
rect 1548 324 1550 332
rect 1558 324 1560 332
rect 1568 324 1570 332
rect 1578 324 1580 332
rect 1588 324 1590 332
rect 1628 324 1630 332
rect 1638 324 1640 332
rect 1648 324 1650 332
rect 1658 324 1660 332
rect 1668 324 1670 332
rect 1678 324 1680 332
rect 1688 324 1690 332
rect 1698 324 1700 332
rect 1708 324 1710 332
rect 1718 324 1732 332
tri 1732 324 1740 332 nw
tri 1748 324 1756 332 se
rect 1756 324 1760 332
rect 1142 322 1160 324
tri 1160 322 1162 324 nw
tri 1176 322 1178 324 se
rect 1178 322 1194 324
rect 1202 322 1284 324
rect 1312 322 1424 324
tri 1424 322 1426 324 nw
tri 1492 322 1494 324 se
rect 1494 322 1590 324
rect 1618 322 1730 324
tri 1730 322 1732 324 nw
tri 1746 322 1748 324 se
rect 1748 322 1760 324
rect 1142 314 1152 322
tri 1152 314 1160 322 nw
tri 1168 314 1176 322 se
rect 1176 314 1184 322
rect 1202 314 1204 322
rect 1212 314 1214 322
rect 1222 314 1224 322
rect 1232 314 1234 322
rect 1242 314 1244 322
rect 1252 314 1254 322
rect 1262 314 1264 322
rect 1272 314 1274 322
rect 1312 314 1314 322
rect 1322 314 1324 322
rect 1332 314 1334 322
rect 1342 314 1344 322
rect 1352 314 1354 322
rect 1362 314 1364 322
rect 1372 314 1374 322
rect 1382 314 1384 322
rect 1392 314 1394 322
rect 1402 314 1404 322
rect 1412 314 1416 322
tri 1416 314 1424 322 nw
tri 1484 314 1492 322 se
rect 1492 314 1500 322
rect 1508 314 1510 322
rect 1518 314 1520 322
rect 1528 314 1530 322
rect 1538 314 1540 322
rect 1548 314 1550 322
rect 1558 314 1560 322
rect 1568 314 1570 322
rect 1578 314 1580 322
rect 1618 314 1620 322
rect 1628 314 1630 322
rect 1638 314 1640 322
rect 1648 314 1650 322
rect 1658 314 1660 322
rect 1668 314 1670 322
rect 1678 314 1680 322
rect 1688 314 1690 322
rect 1698 314 1700 322
rect 1708 314 1722 322
tri 1722 314 1730 322 nw
tri 1738 314 1746 322 se
rect 1746 314 1750 322
rect 1132 312 1150 314
tri 1150 312 1152 314 nw
tri 1166 312 1168 314 se
rect 1168 312 1184 314
rect 1192 312 1274 314
rect 1302 312 1414 314
tri 1414 312 1416 314 nw
tri 1482 312 1484 314 se
rect 1484 312 1580 314
rect 1608 312 1720 314
tri 1720 312 1722 314 nw
tri 1736 312 1738 314 se
rect 1738 312 1750 314
rect 1132 304 1142 312
tri 1142 304 1150 312 nw
tri 1158 304 1166 312 se
rect 1166 304 1174 312
rect 1192 304 1194 312
rect 1202 304 1204 312
rect 1212 304 1214 312
rect 1222 304 1224 312
rect 1232 304 1234 312
rect 1242 304 1244 312
rect 1252 304 1254 312
rect 1262 304 1264 312
rect 1302 304 1304 312
rect 1312 304 1314 312
rect 1322 304 1324 312
rect 1332 304 1334 312
rect 1342 304 1344 312
rect 1352 304 1354 312
rect 1362 304 1364 312
rect 1372 304 1374 312
rect 1382 304 1384 312
rect 1392 304 1394 312
rect 1402 304 1406 312
tri 1406 304 1414 312 nw
tri 1474 304 1482 312 se
rect 1482 304 1490 312
rect 1498 304 1500 312
rect 1508 304 1510 312
rect 1518 304 1520 312
rect 1528 304 1530 312
rect 1538 304 1540 312
rect 1548 304 1550 312
rect 1558 304 1560 312
rect 1568 304 1570 312
rect 1608 304 1610 312
rect 1618 304 1620 312
rect 1628 304 1630 312
rect 1638 304 1640 312
rect 1648 304 1650 312
rect 1658 304 1660 312
rect 1668 304 1670 312
rect 1678 304 1680 312
rect 1688 304 1690 312
rect 1698 304 1712 312
tri 1712 304 1720 312 nw
tri 1728 304 1736 312 se
rect 1736 304 1740 312
rect 1122 302 1140 304
tri 1140 302 1142 304 nw
tri 1156 302 1158 304 se
rect 1158 302 1174 304
rect 1182 302 1264 304
rect 1292 302 1404 304
tri 1404 302 1406 304 nw
tri 1472 302 1474 304 se
rect 1474 302 1570 304
rect 1598 302 1710 304
tri 1710 302 1712 304 nw
tri 1726 302 1728 304 se
rect 1728 302 1740 304
rect 1122 294 1132 302
tri 1132 294 1140 302 nw
tri 1148 294 1156 302 se
rect 1156 294 1164 302
rect 1182 294 1184 302
rect 1192 294 1194 302
rect 1202 294 1204 302
rect 1212 294 1214 302
rect 1222 294 1224 302
rect 1232 294 1234 302
rect 1242 294 1244 302
rect 1252 294 1254 302
rect 1292 294 1294 302
rect 1302 294 1304 302
rect 1312 294 1314 302
rect 1322 294 1324 302
rect 1332 294 1334 302
rect 1342 294 1344 302
rect 1352 294 1354 302
rect 1362 294 1364 302
rect 1372 294 1374 302
rect 1382 294 1384 302
rect 1392 294 1396 302
tri 1396 294 1404 302 nw
tri 1464 294 1472 302 se
rect 1472 294 1480 302
rect 1488 294 1490 302
rect 1498 294 1500 302
rect 1508 294 1510 302
rect 1518 294 1520 302
rect 1528 294 1530 302
rect 1538 294 1540 302
rect 1548 294 1550 302
rect 1558 294 1560 302
rect 1598 294 1600 302
rect 1608 294 1610 302
rect 1618 294 1620 302
rect 1628 294 1630 302
rect 1638 294 1640 302
rect 1648 294 1650 302
rect 1658 294 1660 302
rect 1668 294 1670 302
rect 1678 294 1680 302
rect 1688 294 1702 302
tri 1702 294 1710 302 nw
tri 1718 294 1726 302 se
rect 1726 294 1730 302
rect 1112 292 1130 294
tri 1130 292 1132 294 nw
tri 1146 292 1148 294 se
rect 1148 292 1164 294
rect 1172 292 1254 294
rect 1282 292 1394 294
tri 1394 292 1396 294 nw
tri 1462 292 1464 294 se
rect 1464 292 1560 294
rect 1588 292 1700 294
tri 1700 292 1702 294 nw
tri 1716 292 1718 294 se
rect 1718 292 1730 294
rect 1112 284 1122 292
tri 1122 284 1130 292 nw
tri 1138 284 1146 292 se
rect 1146 284 1154 292
rect 1172 284 1174 292
rect 1182 284 1184 292
rect 1192 284 1194 292
rect 1202 284 1204 292
rect 1212 284 1214 292
rect 1222 284 1224 292
rect 1232 284 1234 292
rect 1242 284 1244 292
rect 1282 284 1284 292
rect 1292 284 1294 292
rect 1302 284 1304 292
rect 1312 284 1314 292
rect 1322 284 1324 292
rect 1332 284 1334 292
rect 1342 284 1344 292
rect 1352 284 1354 292
rect 1362 284 1364 292
rect 1372 284 1374 292
rect 1382 284 1386 292
tri 1386 284 1394 292 nw
tri 1454 284 1462 292 se
rect 1462 284 1470 292
rect 1478 284 1480 292
rect 1488 284 1490 292
rect 1498 284 1500 292
rect 1508 284 1510 292
rect 1518 284 1520 292
rect 1528 284 1530 292
rect 1538 284 1540 292
rect 1548 284 1550 292
rect 1588 284 1590 292
rect 1598 284 1600 292
rect 1608 284 1610 292
rect 1618 284 1620 292
rect 1628 284 1630 292
rect 1638 284 1640 292
rect 1648 284 1650 292
rect 1658 284 1660 292
rect 1668 284 1670 292
rect 1678 284 1692 292
tri 1692 284 1700 292 nw
tri 1708 284 1716 292 se
rect 1716 284 1720 292
rect 1112 282 1120 284
tri 1120 282 1122 284 nw
tri 1136 282 1138 284 se
rect 1138 282 1154 284
rect 1162 282 1244 284
rect 1272 282 1384 284
tri 1384 282 1386 284 nw
tri 1452 282 1454 284 se
rect 1454 282 1550 284
rect 1578 282 1690 284
tri 1690 282 1692 284 nw
tri 1706 282 1708 284 se
rect 1708 282 1720 284
tri 1112 274 1120 282 nw
tri 1128 274 1136 282 se
rect 1136 274 1144 282
rect 1162 274 1164 282
rect 1172 274 1174 282
rect 1182 274 1184 282
rect 1192 274 1194 282
rect 1202 274 1204 282
rect 1212 274 1214 282
rect 1222 274 1224 282
rect 1232 274 1234 282
rect 1272 274 1274 282
rect 1282 274 1284 282
rect 1292 274 1294 282
rect 1302 274 1304 282
rect 1312 274 1314 282
rect 1322 274 1324 282
rect 1332 274 1334 282
rect 1342 274 1344 282
rect 1352 274 1354 282
rect 1362 274 1364 282
rect 1372 274 1376 282
tri 1376 274 1384 282 nw
tri 1444 274 1452 282 se
rect 1452 274 1460 282
rect 1468 274 1470 282
rect 1478 274 1480 282
rect 1488 274 1490 282
rect 1498 274 1500 282
rect 1508 274 1510 282
rect 1518 274 1520 282
rect 1528 274 1530 282
rect 1538 274 1540 282
rect 1578 274 1580 282
rect 1588 274 1590 282
rect 1598 274 1600 282
rect 1608 274 1610 282
rect 1618 274 1620 282
rect 1628 274 1630 282
rect 1638 274 1640 282
rect 1648 274 1650 282
rect 1658 274 1660 282
rect 1668 274 1682 282
tri 1682 274 1690 282 nw
tri 1698 274 1706 282 se
rect 1706 274 1710 282
rect 1092 272 1110 274
tri 1110 272 1112 274 nw
tri 1126 272 1128 274 se
rect 1128 272 1144 274
rect 1152 272 1234 274
rect 1262 272 1374 274
tri 1374 272 1376 274 nw
tri 1442 272 1444 274 se
rect 1444 272 1540 274
rect 1568 272 1680 274
tri 1680 272 1682 274 nw
tri 1696 272 1698 274 se
rect 1698 272 1710 274
rect 1092 264 1102 272
tri 1102 264 1110 272 nw
tri 1118 264 1126 272 se
rect 1126 264 1134 272
rect 1092 262 1100 264
tri 1100 262 1102 264 nw
tri 1116 262 1118 264 se
rect 1118 262 1134 264
rect 1092 254 1094 262
tri 1094 256 1100 262 nw
tri 1110 256 1116 262 se
rect 1116 256 1134 262
tri 1094 254 1096 256 sw
tri 1108 254 1110 256 se
rect 1110 254 1134 256
rect 1092 252 1096 254
tri 1096 252 1098 254 sw
tri 1106 252 1108 254 se
rect 1108 252 1134 254
rect 1092 248 1098 252
tri 1098 248 1102 252 sw
tri 1102 248 1106 252 se
rect 1106 248 1134 252
rect 1092 242 1134 248
rect 1152 244 1154 272
rect 1162 244 1164 272
rect 1172 244 1174 272
rect 1182 244 1184 272
rect 1192 264 1194 272
rect 1202 264 1204 272
rect 1212 264 1214 272
rect 1222 264 1224 272
rect 1192 262 1224 264
rect 1232 262 1244 264
rect 1202 244 1204 262
rect 1212 244 1214 262
rect 1232 244 1234 262
rect 1242 244 1244 262
rect 1262 244 1264 272
rect 1272 244 1274 272
rect 1282 264 1284 272
rect 1292 264 1294 272
rect 1302 264 1304 272
rect 1312 264 1314 272
rect 1282 262 1314 264
rect 1292 244 1294 262
rect 1302 244 1304 262
rect 1322 244 1324 272
rect 1332 244 1334 272
rect 1342 264 1344 272
rect 1352 264 1354 272
rect 1362 264 1366 272
tri 1366 264 1374 272 nw
tri 1434 264 1442 272 se
rect 1442 264 1450 272
rect 1458 264 1460 272
rect 1468 264 1470 272
rect 1478 264 1480 272
rect 1488 264 1490 272
rect 1498 264 1500 272
rect 1508 264 1510 272
rect 1518 264 1520 272
rect 1528 264 1530 272
rect 1568 264 1570 272
rect 1578 264 1580 272
rect 1588 264 1590 272
rect 1598 264 1600 272
rect 1608 264 1610 272
rect 1618 264 1620 272
rect 1628 264 1630 272
rect 1638 264 1640 272
rect 1648 264 1650 272
rect 1658 264 1672 272
tri 1672 264 1680 272 nw
tri 1688 264 1696 272 se
rect 1696 264 1700 272
rect 1342 262 1364 264
tri 1364 262 1366 264 nw
tri 1432 262 1434 264 se
rect 1434 262 1530 264
rect 1558 262 1670 264
tri 1670 262 1672 264 nw
tri 1686 262 1688 264 se
rect 1688 262 1700 264
rect 1352 254 1356 262
tri 1356 254 1364 262 nw
tri 1424 254 1432 262 se
rect 1432 254 1440 262
rect 1448 254 1450 262
rect 1458 254 1460 262
rect 1468 254 1470 262
rect 1478 254 1480 262
rect 1488 254 1490 262
rect 1498 254 1500 262
rect 1508 254 1510 262
rect 1518 254 1520 262
rect 1558 254 1560 262
rect 1568 254 1570 262
rect 1578 254 1580 262
rect 1588 254 1590 262
rect 1598 254 1600 262
rect 1608 254 1610 262
rect 1618 254 1620 262
rect 1628 254 1630 262
rect 1638 254 1640 262
rect 1648 254 1662 262
tri 1662 254 1670 262 nw
tri 1678 254 1686 262 se
rect 1686 254 1690 262
rect 1342 252 1354 254
tri 1354 252 1356 254 nw
tri 1422 252 1424 254 se
rect 1424 252 1520 254
rect 1548 252 1660 254
tri 1660 252 1662 254 nw
tri 1676 252 1678 254 se
rect 1678 252 1690 254
rect 1342 244 1346 252
tri 1346 244 1354 252 nw
tri 1414 244 1422 252 se
rect 1422 244 1430 252
rect 1438 244 1440 252
rect 1448 244 1450 252
rect 1458 244 1460 252
rect 1468 244 1470 252
rect 1478 244 1480 252
rect 1488 244 1490 252
rect 1498 244 1500 252
rect 1508 244 1510 252
rect 1548 244 1550 252
rect 1558 244 1560 252
rect 1568 244 1570 252
rect 1578 244 1580 252
rect 1588 244 1590 252
rect 1598 244 1600 252
rect 1608 244 1610 252
rect 1618 244 1620 252
rect 1628 244 1630 252
rect 1638 244 1652 252
tri 1652 244 1660 252 nw
tri 1668 244 1676 252 se
rect 1676 244 1680 252
rect 1152 242 1184 244
rect 1192 242 1214 244
rect 1222 242 1244 244
rect 1252 242 1274 244
rect 1282 242 1304 244
rect 1312 242 1344 244
tri 1344 242 1346 244 nw
tri 1412 242 1414 244 se
rect 1414 242 1510 244
rect 1538 242 1650 244
tri 1650 242 1652 244 nw
tri 1666 242 1668 244 se
rect 1668 242 1680 244
rect 1162 234 1164 242
rect 1172 234 1174 242
rect 1192 234 1194 242
rect 1202 234 1204 242
rect 1222 234 1224 242
rect 1232 234 1234 242
rect 1252 234 1254 242
rect 1262 234 1264 242
rect 1282 234 1284 242
rect 1292 234 1294 242
rect 1312 234 1314 242
rect 1322 234 1324 242
rect 1332 234 1336 242
tri 1336 234 1344 242 nw
tri 1404 234 1412 242 se
rect 1412 234 1420 242
rect 1428 234 1430 242
rect 1438 234 1440 242
rect 1448 234 1450 242
rect 1458 234 1460 242
rect 1468 234 1470 242
rect 1478 234 1480 242
rect 1488 234 1490 242
rect 1498 234 1500 242
rect 1538 234 1540 242
rect 1548 234 1550 242
rect 1558 234 1560 242
rect 1568 234 1570 242
rect 1578 234 1580 242
rect 1588 234 1590 242
rect 1598 234 1600 242
rect 1608 234 1610 242
rect 1618 234 1620 242
rect 1628 234 1642 242
tri 1642 234 1650 242 nw
tri 1658 234 1666 242 se
rect 1666 234 1670 242
rect 1162 232 1184 234
rect 1192 232 1214 234
rect 1222 232 1244 234
rect 1252 232 1274 234
rect 1282 232 1304 234
rect 1312 232 1334 234
tri 1334 232 1336 234 nw
tri 1402 232 1404 234 se
rect 1404 232 1500 234
rect 1528 232 1640 234
tri 1640 232 1642 234 nw
tri 1656 232 1658 234 se
rect 1658 232 1670 234
rect 1172 224 1174 232
rect 1182 224 1184 232
rect 1202 224 1204 232
rect 1212 224 1214 232
rect 1232 224 1234 232
rect 1242 224 1244 232
rect 1262 224 1264 232
rect 1272 224 1274 232
rect 1292 224 1294 232
rect 1302 224 1304 232
rect 1322 224 1326 232
tri 1326 224 1334 232 nw
tri 1394 224 1402 232 se
rect 1402 224 1410 232
rect 1418 224 1420 232
rect 1428 224 1430 232
rect 1438 224 1440 232
rect 1448 224 1450 232
rect 1458 224 1460 232
rect 1468 224 1470 232
rect 1478 224 1480 232
rect 1488 224 1490 232
rect 1528 224 1530 232
rect 1538 224 1540 232
rect 1548 224 1550 232
rect 1558 224 1560 232
rect 1568 224 1570 232
rect 1578 224 1580 232
rect 1588 224 1590 232
rect 1598 224 1600 232
rect 1608 224 1610 232
rect 1618 224 1632 232
tri 1632 224 1640 232 nw
tri 1648 224 1656 232 se
rect 1656 224 1660 232
rect 1162 222 1184 224
rect 1192 222 1214 224
rect 1222 222 1244 224
rect 1252 222 1274 224
rect 1282 222 1304 224
rect 1312 222 1324 224
tri 1324 222 1326 224 nw
tri 1392 222 1394 224 se
rect 1394 222 1490 224
rect 1518 222 1630 224
tri 1630 222 1632 224 nw
tri 1646 222 1648 224 se
rect 1648 222 1660 224
rect 1162 214 1164 222
rect 1172 214 1174 222
rect 1192 214 1194 222
rect 1202 214 1204 222
rect 1222 214 1224 222
rect 1232 214 1234 222
rect 1252 214 1254 222
rect 1262 214 1264 222
rect 1282 214 1284 222
rect 1292 214 1294 222
rect 1312 214 1316 222
tri 1316 214 1324 222 nw
tri 1384 214 1392 222 se
rect 1392 214 1400 222
rect 1408 214 1410 222
rect 1418 214 1420 222
rect 1428 214 1430 222
rect 1438 214 1440 222
rect 1448 214 1450 222
rect 1458 214 1460 222
rect 1468 214 1470 222
rect 1478 214 1480 222
rect 1518 214 1520 222
rect 1528 214 1530 222
rect 1538 214 1540 222
rect 1548 214 1550 222
rect 1558 214 1560 222
rect 1568 214 1570 222
rect 1578 214 1580 222
rect 1588 214 1590 222
rect 1598 214 1600 222
rect 1608 214 1622 222
tri 1622 214 1630 222 nw
tri 1638 214 1646 222 se
rect 1646 214 1650 222
rect 1162 212 1184 214
rect 1192 212 1214 214
rect 1222 212 1244 214
rect 1252 212 1274 214
rect 1282 212 1304 214
rect 1172 204 1174 212
rect 1182 204 1184 212
rect 1202 204 1204 212
rect 1212 204 1214 212
rect 1232 204 1234 212
rect 1242 204 1244 212
rect 1262 204 1264 212
rect 1272 204 1274 212
rect 1292 204 1294 212
rect 1302 204 1304 212
rect 1162 202 1184 204
rect 1192 202 1214 204
rect 1222 202 1244 204
rect 1252 202 1274 204
rect 1282 202 1304 204
rect 1312 212 1314 214
tri 1314 212 1316 214 nw
tri 1382 212 1384 214 se
rect 1384 212 1480 214
rect 1508 212 1620 214
tri 1620 212 1622 214 nw
tri 1636 212 1638 214 se
rect 1638 212 1650 214
tri 1312 210 1314 212 nw
tri 1380 210 1382 212 se
rect 1382 210 1390 212
tri 1374 204 1380 210 se
rect 1380 204 1390 210
rect 1398 204 1400 212
rect 1408 204 1410 212
rect 1418 204 1420 212
rect 1428 204 1430 212
rect 1438 204 1440 212
rect 1448 204 1450 212
rect 1458 204 1460 212
rect 1468 204 1470 212
rect 1508 204 1510 212
rect 1518 204 1520 212
rect 1528 204 1530 212
rect 1538 204 1540 212
rect 1548 204 1550 212
rect 1558 204 1560 212
rect 1568 204 1570 212
rect 1578 204 1580 212
rect 1588 204 1590 212
rect 1598 204 1612 212
tri 1612 204 1620 212 nw
tri 1628 204 1636 212 se
rect 1636 204 1640 212
tri 1372 202 1374 204 se
rect 1374 202 1470 204
rect 1498 202 1610 204
tri 1610 202 1612 204 nw
tri 1626 202 1628 204 se
rect 1628 202 1640 204
rect 1162 194 1164 202
rect 1172 194 1174 202
rect 1192 194 1194 202
rect 1202 194 1204 202
rect 1222 194 1224 202
rect 1232 194 1234 202
rect 1252 194 1254 202
rect 1262 194 1264 202
rect 1282 194 1284 202
rect 1292 194 1294 202
tri 1364 194 1372 202 se
rect 1372 194 1380 202
rect 1388 194 1390 202
rect 1398 194 1400 202
rect 1408 194 1410 202
rect 1418 194 1420 202
rect 1428 194 1430 202
rect 1438 194 1440 202
rect 1448 194 1450 202
rect 1458 194 1460 202
rect 1498 194 1500 202
rect 1508 194 1510 202
rect 1518 194 1520 202
rect 1528 194 1530 202
rect 1538 194 1540 202
rect 1548 194 1550 202
rect 1558 194 1560 202
rect 1568 194 1570 202
rect 1578 194 1580 202
rect 1588 194 1602 202
tri 1602 194 1610 202 nw
tri 1618 194 1626 202 se
rect 1626 194 1630 202
rect 1162 192 1184 194
rect 1192 192 1214 194
rect 1222 192 1244 194
rect 1252 192 1274 194
rect 1282 192 1304 194
rect 1172 184 1174 192
rect 1182 184 1184 192
rect 1202 184 1204 192
rect 1212 184 1214 192
rect 1232 184 1234 192
rect 1242 184 1244 192
rect 1262 184 1264 192
rect 1272 184 1274 192
rect 1292 184 1294 192
rect 1302 184 1304 192
rect 1162 182 1184 184
rect 1192 182 1214 184
rect 1222 182 1244 184
rect 1252 182 1274 184
rect 1282 182 1304 184
tri 1362 192 1364 194 se
rect 1364 192 1460 194
rect 1488 192 1600 194
tri 1600 192 1602 194 nw
tri 1616 192 1618 194 se
rect 1618 192 1630 194
tri 1354 184 1362 192 se
rect 1362 184 1370 192
tri 1352 182 1354 184 se
rect 1354 182 1370 184
rect 1378 184 1380 192
rect 1388 184 1390 192
rect 1378 182 1390 184
rect 1398 184 1400 192
rect 1408 184 1410 192
rect 1398 182 1410 184
rect 1418 184 1420 192
rect 1428 184 1430 192
rect 1418 182 1430 184
rect 1438 184 1440 192
rect 1448 184 1450 192
rect 1438 182 1450 184
rect 1488 184 1490 192
rect 1498 184 1500 192
rect 1488 182 1500 184
rect 1508 184 1510 192
rect 1518 184 1520 192
rect 1508 182 1520 184
rect 1528 184 1530 192
rect 1538 184 1540 192
rect 1528 182 1540 184
rect 1548 184 1550 192
rect 1558 184 1560 192
rect 1548 182 1560 184
rect 1568 184 1570 192
rect 1578 184 1592 192
tri 1592 184 1600 192 nw
tri 1608 184 1616 192 se
rect 1616 184 1620 192
rect 1568 182 1590 184
tri 1590 182 1592 184 nw
tri 1606 182 1608 184 se
rect 1608 182 1620 184
rect 1162 174 1164 182
rect 1172 174 1174 182
rect 1192 174 1194 182
rect 1202 174 1204 182
rect 1222 174 1224 182
rect 1232 174 1234 182
rect 1252 174 1254 182
rect 1262 174 1264 182
rect 1282 174 1284 182
rect 1292 174 1294 182
rect 1162 172 1184 174
rect 1192 172 1214 174
rect 1222 172 1244 174
rect 1252 172 1274 174
rect 1282 172 1304 174
rect 1172 164 1174 172
rect 1182 164 1184 172
rect 1202 164 1204 172
rect 1212 164 1214 172
rect 1232 164 1234 172
rect 1242 164 1244 172
rect 1262 164 1264 172
rect 1272 164 1274 172
rect 1292 164 1294 172
rect 1302 164 1304 172
rect 1162 162 1184 164
rect 1192 162 1214 164
rect 1222 162 1244 164
rect 1252 162 1274 164
rect 1282 162 1304 164
rect 1162 154 1164 162
rect 1172 154 1174 162
rect 1192 154 1194 162
rect 1202 154 1204 162
rect 1222 154 1224 162
rect 1232 154 1234 162
rect 1252 154 1254 162
rect 1262 154 1264 162
rect 1282 154 1284 162
rect 1292 154 1294 162
rect 1162 152 1184 154
rect 1192 152 1214 154
rect 1222 152 1244 154
rect 1252 152 1274 154
rect 1282 152 1304 154
rect 1172 144 1174 152
rect 1182 144 1184 152
rect 1202 144 1204 152
rect 1212 144 1214 152
rect 1232 144 1234 152
rect 1242 144 1244 152
rect 1262 144 1264 152
rect 1272 144 1274 152
rect 1292 144 1294 152
rect 1302 144 1304 152
rect 1162 142 1184 144
rect 1192 142 1214 144
rect 1222 142 1244 144
rect 1252 142 1274 144
rect 1282 142 1304 144
rect 1162 134 1164 142
rect 1172 134 1174 142
rect 1192 134 1194 142
rect 1202 134 1204 142
rect 1222 134 1224 142
rect 1232 134 1234 142
rect 1252 134 1254 142
rect 1262 134 1264 142
rect 1282 134 1284 142
rect 1292 134 1294 142
rect 1162 132 1184 134
rect 1192 132 1214 134
rect 1222 132 1244 134
rect 1252 132 1274 134
rect 1282 132 1304 134
rect 1172 124 1174 132
rect 1182 124 1184 132
rect 1202 124 1204 132
rect 1212 124 1214 132
rect 1232 124 1234 132
rect 1242 124 1244 132
rect 1262 124 1264 132
rect 1272 124 1274 132
rect 1292 124 1294 132
rect 1302 124 1304 132
rect 1162 122 1184 124
rect 1192 122 1214 124
rect 1222 122 1244 124
rect 1252 122 1274 124
rect 1282 122 1304 124
rect 1162 114 1164 122
rect 1172 114 1174 122
rect 1192 114 1194 122
rect 1202 114 1204 122
rect 1222 114 1224 122
rect 1232 114 1234 122
rect 1252 114 1254 122
rect 1262 114 1264 122
rect 1282 114 1284 122
rect 1292 114 1294 122
rect 1162 112 1184 114
rect 1192 112 1214 114
rect 1222 112 1244 114
rect 1252 112 1274 114
rect 1282 112 1304 114
rect 1172 104 1174 112
rect 1182 104 1184 112
rect 1202 104 1204 112
rect 1212 104 1214 112
rect 1232 104 1234 112
rect 1242 104 1244 112
rect 1262 104 1264 112
rect 1272 104 1274 112
rect 1292 104 1294 112
rect 1302 104 1304 112
rect 1162 102 1184 104
rect 1192 102 1214 104
rect 1222 102 1244 104
rect 1252 102 1274 104
rect 1282 102 1304 104
rect 1162 94 1164 102
rect 1172 94 1174 102
rect 1192 94 1194 102
rect 1202 94 1204 102
rect 1222 94 1224 102
rect 1232 94 1234 102
rect 1252 94 1254 102
rect 1262 94 1264 102
rect 1282 94 1284 102
rect 1292 94 1294 102
rect 1162 92 1184 94
rect 1192 92 1214 94
rect 1222 92 1244 94
rect 1252 92 1274 94
rect 1282 92 1304 94
rect 1172 84 1174 92
rect 1182 84 1184 92
rect 1202 84 1204 92
rect 1212 84 1214 92
rect 1232 84 1234 92
rect 1242 84 1244 92
rect 1262 84 1264 92
rect 1272 84 1274 92
rect 1292 84 1294 92
rect 1302 84 1304 92
rect 1162 82 1184 84
rect 1192 82 1214 84
rect 1222 82 1244 84
rect 1252 82 1274 84
rect 1282 82 1304 84
rect 1162 74 1164 82
rect 1172 74 1174 82
rect 1192 74 1194 82
rect 1202 74 1204 82
rect 1222 74 1224 82
rect 1232 74 1234 82
rect 1252 74 1254 82
rect 1262 74 1264 82
rect 1282 74 1284 82
rect 1292 74 1294 82
rect 1162 72 1184 74
rect 1192 72 1214 74
rect 1222 72 1244 74
rect 1252 72 1274 74
rect 1282 72 1304 74
rect 1172 64 1174 72
rect 1182 64 1184 72
rect 1202 64 1204 72
rect 1212 64 1214 72
rect 1232 64 1234 72
rect 1242 64 1244 72
rect 1262 64 1264 72
rect 1272 64 1274 72
rect 1292 64 1294 72
rect 1302 64 1304 72
rect 1162 62 1184 64
rect 1192 62 1214 64
rect 1222 62 1244 64
rect 1252 62 1274 64
rect 1282 62 1304 64
rect 1162 54 1164 62
rect 1172 54 1174 62
rect 1192 54 1194 62
rect 1202 54 1204 62
rect 1222 54 1224 62
rect 1232 54 1234 62
rect 1252 54 1254 62
rect 1262 54 1264 62
rect 1282 54 1284 62
rect 1292 54 1294 62
rect 1162 52 1184 54
rect 1192 52 1214 54
rect 1222 52 1244 54
rect 1252 52 1274 54
rect 1282 52 1304 54
rect 1172 44 1174 52
rect 1182 44 1184 52
rect 1202 44 1204 52
rect 1212 44 1214 52
rect 1232 44 1234 52
rect 1242 44 1244 52
rect 1262 44 1264 52
rect 1272 44 1274 52
rect 1292 44 1294 52
rect 1302 44 1304 52
rect 1162 42 1184 44
rect 1192 42 1214 44
rect 1222 42 1244 44
rect 1252 42 1274 44
rect 1282 42 1304 44
rect 1162 34 1164 42
rect 1172 34 1174 42
rect 1192 34 1194 42
rect 1202 34 1204 42
rect 1222 34 1224 42
rect 1232 34 1234 42
rect 1252 34 1254 42
rect 1262 34 1264 42
rect 1282 34 1284 42
rect 1292 34 1294 42
rect 1162 32 1184 34
rect 1192 32 1214 34
rect 1222 32 1244 34
rect 1252 32 1274 34
rect 1282 32 1304 34
rect 1172 24 1174 32
rect 1182 24 1184 32
rect 1202 24 1204 32
rect 1212 24 1214 32
rect 1232 24 1234 32
rect 1242 24 1244 32
rect 1262 24 1264 32
rect 1272 24 1274 32
rect 1292 24 1294 32
rect 1302 24 1304 32
rect 1162 22 1184 24
rect 1192 22 1214 24
rect 1222 22 1244 24
rect 1252 22 1274 24
rect 1282 22 1304 24
rect 1162 14 1164 22
rect 1172 14 1174 22
rect 1192 14 1194 22
rect 1202 14 1204 22
rect 1222 14 1224 22
rect 1232 14 1234 22
rect 1252 14 1254 22
rect 1262 14 1264 22
rect 1282 14 1284 22
rect 1292 14 1294 22
rect 1162 12 1184 14
rect 1192 12 1214 14
rect 1222 12 1244 14
rect 1252 12 1274 14
rect 1282 12 1304 14
rect 1172 4 1174 12
rect 1182 4 1184 12
rect 1202 4 1204 12
rect 1212 4 1214 12
rect 1232 4 1234 12
rect 1242 4 1244 12
rect 1262 4 1264 12
rect 1272 4 1274 12
rect 1292 4 1294 12
rect 1302 4 1304 12
rect 662 0 1312 4
tri 1348 178 1352 182 se
rect 1352 178 1360 182
rect 1348 174 1360 178
rect 1568 178 1586 182
tri 1586 178 1590 182 nw
tri 1602 178 1606 182 se
rect 1606 178 1610 182
rect 1568 174 1582 178
tri 1582 174 1586 178 nw
tri 1598 174 1602 178 se
rect 1602 174 1610 178
rect 1348 172 1370 174
rect 1348 4 1350 172
rect 1358 144 1360 172
rect 1368 144 1370 172
rect 1378 172 1390 174
rect 1378 144 1380 172
rect 1388 144 1390 172
rect 1358 142 1390 144
rect 1398 172 1410 174
rect 1368 134 1370 142
rect 1378 134 1380 142
rect 1398 134 1400 172
rect 1408 134 1410 172
rect 1418 172 1430 174
rect 1418 144 1420 172
rect 1428 144 1430 172
rect 1468 172 1480 174
rect 1468 144 1470 172
rect 1478 144 1480 172
rect 1418 142 1440 144
rect 1428 134 1430 142
rect 1438 134 1440 142
rect 1458 142 1480 144
rect 1488 172 1500 174
rect 1458 134 1460 142
rect 1468 134 1470 142
rect 1488 134 1490 172
rect 1498 134 1500 172
rect 1508 172 1520 174
rect 1508 144 1510 172
rect 1518 144 1520 172
rect 1508 142 1520 144
rect 1528 172 1540 174
rect 1528 144 1530 172
rect 1538 144 1540 172
rect 1528 142 1540 144
rect 1548 172 1580 174
tri 1580 172 1582 174 nw
tri 1596 172 1598 174 se
rect 1598 172 1610 174
rect 1548 164 1550 172
rect 1558 164 1572 172
tri 1572 164 1580 172 nw
tri 1588 164 1596 172 se
rect 1596 164 1600 172
rect 1548 162 1570 164
tri 1570 162 1572 164 nw
tri 1586 162 1588 164 se
rect 1588 162 1600 164
rect 1548 154 1567 162
tri 1567 159 1570 162 nw
tri 1583 159 1586 162 se
rect 1586 159 1590 162
tri 1567 154 1572 159 sw
tri 1578 154 1583 159 se
rect 1583 154 1590 159
rect 1548 152 1572 154
tri 1572 152 1574 154 sw
tri 1576 152 1578 154 se
rect 1578 152 1590 154
rect 1548 151 1574 152
tri 1574 151 1575 152 sw
tri 1575 151 1576 152 se
rect 1576 151 1580 152
rect 1548 142 1580 151
rect 1358 132 1380 134
rect 1388 132 1410 134
rect 1418 132 1440 134
rect 1448 132 1470 134
rect 1478 132 1500 134
rect 1358 124 1360 132
rect 1368 124 1370 132
rect 1388 124 1390 132
rect 1398 124 1400 132
rect 1418 124 1420 132
rect 1428 124 1430 132
rect 1448 124 1450 132
rect 1458 124 1460 132
rect 1478 124 1480 132
rect 1488 124 1490 132
rect 1358 122 1380 124
rect 1388 122 1410 124
rect 1418 122 1440 124
rect 1448 122 1470 124
rect 1478 122 1500 124
rect 1368 114 1370 122
rect 1378 114 1380 122
rect 1398 114 1400 122
rect 1408 114 1410 122
rect 1428 114 1430 122
rect 1438 114 1440 122
rect 1458 114 1460 122
rect 1468 114 1470 122
rect 1488 114 1490 122
rect 1498 114 1500 122
rect 1358 112 1380 114
rect 1388 112 1410 114
rect 1418 112 1440 114
rect 1448 112 1470 114
rect 1478 112 1500 114
rect 1358 104 1360 112
rect 1368 104 1370 112
rect 1388 104 1390 112
rect 1398 104 1400 112
rect 1418 104 1420 112
rect 1428 104 1430 112
rect 1448 104 1450 112
rect 1458 104 1460 112
rect 1478 104 1480 112
rect 1488 104 1490 112
rect 1358 102 1380 104
rect 1388 102 1410 104
rect 1418 102 1440 104
rect 1448 102 1470 104
rect 1478 102 1500 104
rect 1368 94 1370 102
rect 1378 94 1380 102
rect 1398 94 1400 102
rect 1408 94 1410 102
rect 1428 94 1430 102
rect 1438 94 1440 102
rect 1458 94 1460 102
rect 1468 94 1470 102
rect 1488 94 1490 102
rect 1498 94 1500 102
rect 1358 92 1380 94
rect 1388 92 1410 94
rect 1418 92 1440 94
rect 1448 92 1470 94
rect 1478 92 1500 94
rect 1358 84 1360 92
rect 1368 84 1370 92
rect 1388 84 1390 92
rect 1398 84 1400 92
rect 1418 84 1420 92
rect 1428 84 1430 92
rect 1448 84 1450 92
rect 1458 84 1460 92
rect 1478 84 1480 92
rect 1488 84 1490 92
rect 1358 82 1380 84
rect 1388 82 1410 84
rect 1418 82 1440 84
rect 1448 82 1470 84
rect 1478 82 1500 84
rect 1368 74 1370 82
rect 1378 74 1380 82
rect 1398 74 1400 82
rect 1408 74 1410 82
rect 1428 74 1430 82
rect 1438 74 1440 82
rect 1458 74 1460 82
rect 1468 74 1470 82
rect 1488 74 1490 82
rect 1498 74 1500 82
rect 1358 72 1380 74
rect 1388 72 1410 74
rect 1418 72 1440 74
rect 1448 72 1470 74
rect 1478 72 1500 74
rect 1358 64 1360 72
rect 1368 64 1370 72
rect 1388 64 1390 72
rect 1398 64 1400 72
rect 1418 64 1420 72
rect 1428 64 1430 72
rect 1448 64 1450 72
rect 1458 64 1460 72
rect 1478 64 1480 72
rect 1488 64 1490 72
rect 1358 62 1380 64
rect 1388 62 1410 64
rect 1418 62 1440 64
rect 1448 62 1470 64
rect 1478 62 1500 64
rect 1368 54 1370 62
rect 1378 54 1380 62
rect 1398 54 1400 62
rect 1408 54 1410 62
rect 1428 54 1430 62
rect 1438 54 1440 62
rect 1458 54 1460 62
rect 1468 54 1470 62
rect 1488 54 1490 62
rect 1498 54 1500 62
rect 1358 52 1380 54
rect 1388 52 1410 54
rect 1418 52 1440 54
rect 1448 52 1470 54
rect 1478 52 1500 54
rect 1358 44 1360 52
rect 1368 44 1370 52
rect 1388 44 1390 52
rect 1398 44 1400 52
rect 1418 44 1420 52
rect 1428 44 1430 52
rect 1448 44 1450 52
rect 1458 44 1460 52
rect 1478 44 1480 52
rect 1488 44 1490 52
rect 1358 42 1380 44
rect 1388 42 1410 44
rect 1418 42 1440 44
rect 1448 42 1470 44
rect 1478 42 1500 44
rect 1368 34 1370 42
rect 1378 34 1380 42
rect 1398 34 1400 42
rect 1408 34 1410 42
rect 1428 34 1430 42
rect 1438 34 1440 42
rect 1458 34 1460 42
rect 1468 34 1470 42
rect 1488 34 1490 42
rect 1498 34 1500 42
rect 1358 32 1380 34
rect 1388 32 1410 34
rect 1418 32 1440 34
rect 1448 32 1470 34
rect 1478 32 1500 34
rect 1358 24 1360 32
rect 1368 24 1370 32
rect 1388 24 1390 32
rect 1398 24 1400 32
rect 1418 24 1420 32
rect 1428 24 1430 32
rect 1448 24 1450 32
rect 1458 24 1460 32
rect 1478 24 1480 32
rect 1488 24 1490 32
rect 1358 22 1380 24
rect 1388 22 1410 24
rect 1418 22 1440 24
rect 1448 22 1470 24
rect 1478 22 1500 24
rect 1368 14 1370 22
rect 1378 14 1380 22
rect 1398 14 1400 22
rect 1408 14 1410 22
rect 1428 14 1430 22
rect 1438 14 1440 22
rect 1458 14 1460 22
rect 1468 14 1470 22
rect 1488 14 1490 22
rect 1498 14 1500 22
rect 1358 12 1380 14
rect 1388 12 1410 14
rect 1418 12 1440 14
rect 1448 12 1470 14
rect 1478 12 1500 14
rect 1358 4 1360 12
rect 1368 4 1370 12
rect 1388 4 1390 12
rect 1398 4 1400 12
rect 1418 4 1420 12
rect 1428 4 1430 12
rect 1448 4 1450 12
rect 1458 4 1460 12
rect 1478 4 1480 12
rect 1488 4 1490 12
rect 1998 4 2000 502
rect 1348 0 2000 4
<< m2contact >>
rect 1724 834 1732 842
rect 1754 834 1762 842
rect 1784 834 1792 842
rect 1814 834 1822 842
rect 1844 834 1852 842
rect 1874 834 1882 842
rect 1904 834 1912 842
rect 1934 834 1942 842
rect 1964 834 1972 842
rect 1734 824 1742 832
rect 1764 824 1772 832
rect 1794 824 1802 832
rect 1824 824 1832 832
rect 1854 824 1862 832
rect 1884 824 1892 832
rect 1914 824 1922 832
rect 1944 824 1952 832
rect 1974 824 1982 832
rect 1724 814 1732 822
rect 1754 814 1762 822
rect 1784 814 1792 822
rect 1814 814 1822 822
rect 1844 814 1852 822
rect 1874 814 1882 822
rect 1904 814 1912 822
rect 1934 814 1942 822
rect 1964 814 1972 822
rect 1694 804 1702 812
rect 1734 804 1742 812
rect 1764 804 1772 812
rect 1794 804 1802 812
rect 1824 804 1832 812
rect 1854 804 1862 812
rect 1884 804 1892 812
rect 1914 804 1922 812
rect 1944 804 1952 812
rect 1974 804 1982 812
rect 1684 794 1692 802
rect 1724 794 1732 802
rect 1754 794 1762 802
rect 1784 794 1792 802
rect 1814 794 1822 802
rect 1844 794 1852 802
rect 1874 794 1882 802
rect 1904 794 1912 802
rect 1934 794 1942 802
rect 1964 794 1972 802
rect 1674 784 1682 792
rect 1694 784 1702 792
rect 1734 784 1742 792
rect 1764 784 1772 792
rect 1794 784 1802 792
rect 1824 784 1832 792
rect 1854 784 1862 792
rect 1884 784 1892 792
rect 1914 784 1922 792
rect 1944 784 1952 792
rect 1974 784 1982 792
rect 1664 774 1672 782
rect 1684 774 1692 782
rect 1724 774 1732 782
rect 1754 774 1762 782
rect 1784 774 1792 782
rect 1814 774 1822 782
rect 1844 774 1852 782
rect 1874 774 1882 782
rect 1904 774 1912 782
rect 1934 774 1942 782
rect 1964 774 1972 782
rect 1654 764 1662 772
rect 1674 764 1682 772
rect 1734 764 1742 772
rect 1764 764 1772 772
rect 1794 764 1802 772
rect 1824 764 1832 772
rect 1854 764 1862 772
rect 1884 764 1892 772
rect 1914 764 1922 772
rect 1944 764 1952 772
rect 1974 764 1982 772
rect 1644 754 1652 762
rect 1664 754 1672 762
rect 1694 754 1702 762
rect 1724 754 1732 762
rect 1754 754 1762 762
rect 1784 754 1792 762
rect 1814 754 1822 762
rect 1844 754 1852 762
rect 1874 754 1882 762
rect 1904 754 1912 762
rect 1934 754 1942 762
rect 1964 754 1972 762
rect 1634 744 1642 752
rect 1654 744 1662 752
rect 1684 744 1692 752
rect 1734 744 1742 752
rect 1764 744 1772 752
rect 1794 744 1802 752
rect 1824 744 1832 752
rect 1854 744 1862 752
rect 1884 744 1892 752
rect 1914 744 1922 752
rect 1944 744 1952 752
rect 1974 744 1982 752
rect 1624 734 1632 742
rect 1644 734 1652 742
rect 1674 734 1682 742
rect 1724 734 1732 742
rect 1754 734 1762 742
rect 1784 734 1792 742
rect 1814 734 1822 742
rect 1844 734 1852 742
rect 1874 734 1882 742
rect 1904 734 1912 742
rect 1934 734 1942 742
rect 1964 734 1972 742
rect 1614 724 1622 732
rect 1634 724 1642 732
rect 1664 724 1672 732
rect 1734 724 1742 732
rect 1764 724 1772 732
rect 1794 724 1802 732
rect 1824 724 1832 732
rect 1854 724 1862 732
rect 1884 724 1892 732
rect 1914 724 1922 732
rect 1944 724 1952 732
rect 1974 724 1982 732
rect 1604 714 1612 722
rect 1624 714 1632 722
rect 1654 714 1662 722
rect 1724 714 1732 722
rect 1754 714 1762 722
rect 1784 714 1792 722
rect 1814 714 1822 722
rect 1844 714 1852 722
rect 1874 714 1882 722
rect 1904 714 1912 722
rect 1934 714 1942 722
rect 1964 714 1972 722
rect 1594 704 1602 712
rect 1614 704 1622 712
rect 1644 704 1652 712
rect 1734 704 1742 712
rect 1764 704 1772 712
rect 1794 704 1802 712
rect 1824 704 1832 712
rect 1854 704 1862 712
rect 1884 704 1892 712
rect 1914 704 1922 712
rect 1944 704 1952 712
rect 1974 704 1982 712
rect 1584 694 1592 702
rect 1604 694 1612 702
rect 1574 684 1582 692
rect 1594 684 1602 692
rect 1614 684 1622 692
rect 1634 684 1642 702
rect 1694 694 1702 702
rect 1684 684 1692 692
rect 1704 684 1712 692
rect 1724 684 1732 702
rect 1754 694 1762 702
rect 1784 694 1792 702
rect 1814 694 1822 702
rect 1844 694 1852 702
rect 1874 694 1882 702
rect 1904 694 1912 702
rect 1934 694 1942 702
rect 1964 694 1972 702
rect 1744 684 1752 692
rect 1764 684 1772 692
rect 1564 674 1572 682
rect 1584 674 1592 682
rect 1604 674 1612 682
rect 1624 674 1632 682
rect 1674 674 1682 682
rect 1694 674 1702 682
rect 1714 674 1722 682
rect 1734 674 1742 682
rect 1754 674 1762 682
rect 1554 664 1562 672
rect 1574 664 1582 672
rect 1594 664 1602 672
rect 1614 664 1622 672
rect 1664 664 1672 672
rect 1684 664 1692 672
rect 1704 664 1712 672
rect 1724 664 1732 672
rect 1744 664 1752 672
rect 1544 654 1552 662
rect 1564 654 1572 662
rect 1584 654 1592 662
rect 1604 654 1612 662
rect 1654 654 1662 662
rect 1674 654 1682 662
rect 1694 654 1702 662
rect 1714 654 1722 662
rect 1734 654 1742 662
rect 1534 644 1542 652
rect 1554 644 1562 652
rect 1574 644 1582 652
rect 1594 644 1602 652
rect 1644 644 1652 652
rect 1664 644 1672 652
rect 1684 644 1692 652
rect 1704 644 1712 652
rect 1724 644 1732 652
rect 1524 634 1532 642
rect 1544 634 1552 642
rect 1564 634 1572 642
rect 1584 634 1592 642
rect 1634 634 1642 642
rect 1654 634 1662 642
rect 1674 634 1682 642
rect 1694 634 1702 642
rect 1714 634 1722 642
rect 1830 634 1838 642
rect 1860 634 1868 642
rect 1890 634 1898 642
rect 1920 634 1928 642
rect 1950 634 1958 642
rect 1980 634 1988 642
rect 1514 624 1522 632
rect 1534 624 1542 632
rect 1554 624 1562 632
rect 1574 624 1582 632
rect 1624 624 1632 632
rect 1644 624 1652 632
rect 1664 624 1672 632
rect 1684 624 1692 632
rect 1704 624 1712 632
rect 1840 624 1848 632
rect 1870 624 1878 632
rect 1900 624 1908 632
rect 1930 624 1938 632
rect 1960 624 1968 632
rect 1990 624 1998 632
rect 1504 614 1512 622
rect 1524 614 1532 622
rect 1544 614 1552 622
rect 1564 614 1572 622
rect 1614 614 1622 622
rect 1634 614 1642 622
rect 1654 614 1662 622
rect 1674 614 1682 622
rect 1694 614 1702 622
rect 1830 614 1838 622
rect 1860 614 1868 622
rect 1890 614 1898 622
rect 1920 614 1928 622
rect 1950 614 1958 622
rect 1980 614 1988 622
rect 1494 604 1502 612
rect 1514 604 1522 612
rect 1534 604 1542 612
rect 1554 604 1562 612
rect 1604 604 1612 612
rect 1624 604 1632 612
rect 1644 604 1652 612
rect 1664 604 1672 612
rect 1684 604 1692 612
rect 1810 604 1818 612
rect 1840 604 1848 612
rect 1870 604 1878 612
rect 1900 604 1908 612
rect 1930 604 1938 612
rect 1960 604 1968 612
rect 1990 604 1998 612
rect 1484 594 1492 602
rect 1504 594 1512 602
rect 1524 594 1532 602
rect 1544 594 1552 602
rect 1594 594 1602 602
rect 1614 594 1622 602
rect 1634 594 1642 602
rect 1654 594 1662 602
rect 1674 594 1682 602
rect 1800 594 1808 602
rect 1830 594 1838 602
rect 1860 594 1868 602
rect 1890 594 1898 602
rect 1920 594 1928 602
rect 1950 594 1958 602
rect 1980 594 1988 602
rect 1474 584 1482 592
rect 1494 584 1502 592
rect 1514 584 1522 592
rect 1534 584 1542 592
rect 1584 584 1592 592
rect 1604 584 1612 592
rect 1624 584 1632 592
rect 1644 584 1652 592
rect 1664 584 1672 592
rect 1790 584 1798 592
rect 1840 584 1848 592
rect 1464 574 1472 582
rect 1484 574 1492 582
rect 1504 574 1512 582
rect 1524 574 1532 582
rect 1574 574 1582 582
rect 1594 574 1602 582
rect 1614 574 1622 582
rect 1634 574 1642 582
rect 1654 574 1662 582
rect 1780 574 1788 582
rect 1810 574 1818 582
rect 1870 584 1878 592
rect 1900 584 1908 592
rect 1930 584 1938 592
rect 1960 584 1968 592
rect 1990 584 1998 592
rect 1830 574 1838 582
rect 1890 574 1898 582
rect 1920 574 1928 582
rect 1950 574 1958 582
rect 1980 574 1988 582
rect 1454 564 1462 572
rect 1474 564 1482 572
rect 1494 564 1502 572
rect 1514 564 1522 572
rect 1564 564 1572 572
rect 1584 564 1592 572
rect 1604 564 1612 572
rect 1624 564 1632 572
rect 1644 564 1652 572
rect 1770 564 1778 572
rect 1800 564 1808 572
rect 1870 564 1878 572
rect 1900 564 1908 572
rect 1930 564 1938 572
rect 1960 564 1968 572
rect 1990 564 1998 572
rect 1444 554 1452 562
rect 1464 554 1472 562
rect 1484 554 1492 562
rect 1504 554 1512 562
rect 1554 554 1562 562
rect 1574 554 1582 562
rect 1594 554 1602 562
rect 1614 554 1622 562
rect 1634 554 1642 562
rect 1760 554 1768 562
rect 1790 554 1798 562
rect 1860 554 1868 562
rect 1890 554 1898 562
rect 1920 554 1928 562
rect 1950 554 1958 562
rect 1980 554 1988 562
rect 1434 544 1442 552
rect 1454 544 1462 552
rect 1474 544 1482 552
rect 1494 544 1502 552
rect 1544 544 1552 552
rect 1564 544 1572 552
rect 1584 544 1592 552
rect 1604 544 1612 552
rect 1624 544 1632 552
rect 1750 544 1758 552
rect 1780 544 1788 552
rect 1840 544 1848 552
rect 1870 544 1878 552
rect 1900 544 1908 552
rect 1930 544 1938 552
rect 1960 544 1968 552
rect 1990 544 1998 552
rect 1424 534 1432 542
rect 1444 534 1452 542
rect 1464 534 1472 542
rect 1484 534 1492 542
rect 1534 534 1542 542
rect 1554 534 1562 542
rect 1574 534 1582 542
rect 1594 534 1602 542
rect 1614 534 1622 542
rect 1740 534 1748 542
rect 1770 534 1778 542
rect 1830 534 1838 542
rect 1860 534 1868 542
rect 1890 534 1898 542
rect 1920 534 1928 542
rect 1950 534 1958 542
rect 1980 534 1988 542
rect 1414 524 1422 532
rect 1434 524 1442 532
rect 1454 524 1462 532
rect 1474 524 1482 532
rect 1524 524 1532 532
rect 1544 524 1552 532
rect 1564 524 1572 532
rect 1584 524 1592 532
rect 1604 524 1612 532
rect 1730 524 1738 532
rect 1760 524 1768 532
rect 1840 524 1848 532
rect 1870 524 1878 532
rect 1900 524 1908 532
rect 1930 524 1938 532
rect 1960 524 1968 532
rect 1990 524 1998 532
rect 1404 514 1412 522
rect 1424 514 1432 522
rect 1444 514 1452 522
rect 1464 514 1472 522
rect 1514 514 1522 522
rect 1534 514 1542 522
rect 1554 514 1562 522
rect 1574 514 1582 522
rect 1594 514 1602 522
rect 1720 514 1728 522
rect 1750 514 1758 522
rect 1810 514 1818 522
rect 1830 514 1838 522
rect 1860 514 1868 522
rect 1890 514 1898 522
rect 1920 514 1928 522
rect 1950 514 1958 522
rect 1980 514 1988 522
rect 1394 504 1402 512
rect 1414 504 1422 512
rect 1434 504 1442 512
rect 1454 504 1462 512
rect 1504 504 1512 512
rect 1524 504 1532 512
rect 1544 504 1552 512
rect 1564 504 1572 512
rect 1584 504 1592 512
rect 1710 504 1718 512
rect 1740 504 1748 512
rect 1800 504 1808 512
rect 1840 504 1848 512
rect 1870 504 1878 512
rect 1900 504 1908 512
rect 1930 504 1938 512
rect 1960 504 1968 512
rect 1990 504 1998 512
rect 1384 494 1392 502
rect 1404 494 1412 502
rect 1424 494 1432 502
rect 1444 494 1452 502
rect 1494 494 1502 502
rect 1514 494 1522 502
rect 1534 494 1542 502
rect 1554 494 1562 502
rect 1574 494 1582 502
rect 1374 484 1382 492
rect 1394 484 1402 492
rect 1414 484 1422 492
rect 1434 484 1442 492
rect 1484 484 1492 492
rect 1504 484 1512 492
rect 1524 484 1532 492
rect 1544 484 1552 492
rect 1564 484 1572 492
rect 1680 484 1688 492
rect 1700 484 1708 492
rect 1720 484 1728 492
rect 1740 484 1748 492
rect 1790 484 1798 492
rect 1810 484 1818 492
rect 1830 484 1838 492
rect 1850 484 1858 492
rect 1870 484 1878 492
rect 1364 474 1372 482
rect 1384 474 1392 482
rect 1404 474 1412 482
rect 1424 474 1432 482
rect 1474 474 1482 482
rect 1494 474 1502 482
rect 1514 474 1522 482
rect 1534 474 1542 482
rect 1554 474 1562 482
rect 1670 474 1678 482
rect 1690 474 1698 482
rect 1710 474 1718 482
rect 1730 474 1738 482
rect 1780 474 1788 482
rect 1800 474 1808 482
rect 1820 474 1828 482
rect 1840 474 1848 482
rect 1860 474 1868 482
rect 1354 464 1362 472
rect 1374 464 1382 472
rect 1394 464 1402 472
rect 1414 464 1422 472
rect 1464 464 1472 472
rect 1484 464 1492 472
rect 1504 464 1512 472
rect 1524 464 1532 472
rect 1544 464 1552 472
rect 1660 464 1668 472
rect 1680 464 1688 472
rect 1700 464 1708 472
rect 1720 464 1728 472
rect 1770 464 1778 472
rect 1790 464 1798 472
rect 1810 464 1818 472
rect 1830 464 1838 472
rect 1850 464 1858 472
rect 1344 454 1352 462
rect 1364 454 1372 462
rect 1384 454 1392 462
rect 1404 454 1412 462
rect 1454 454 1462 462
rect 1474 454 1482 462
rect 1494 454 1502 462
rect 1514 454 1522 462
rect 1534 454 1542 462
rect 1650 454 1658 462
rect 1670 454 1678 462
rect 1690 454 1698 462
rect 1710 454 1718 462
rect 1760 454 1768 462
rect 1780 454 1788 462
rect 1800 454 1808 462
rect 1820 454 1828 462
rect 1840 454 1848 462
rect 1334 444 1342 452
rect 1354 444 1362 452
rect 1374 444 1382 452
rect 1394 444 1402 452
rect 1444 444 1452 452
rect 1464 444 1472 452
rect 1484 444 1492 452
rect 1504 444 1512 452
rect 1524 444 1532 452
rect 1640 444 1648 452
rect 1660 444 1668 452
rect 1680 444 1688 452
rect 1700 444 1708 452
rect 1750 444 1758 452
rect 1770 444 1778 452
rect 1790 444 1798 452
rect 1810 444 1818 452
rect 1830 444 1838 452
rect 1324 434 1332 442
rect 1344 434 1352 442
rect 1364 434 1372 442
rect 1384 434 1392 442
rect 1434 434 1442 442
rect 1454 434 1462 442
rect 1474 434 1482 442
rect 1494 434 1502 442
rect 1514 434 1522 442
rect 1630 434 1638 442
rect 1650 434 1658 442
rect 1670 434 1678 442
rect 1690 434 1698 442
rect 1740 434 1748 442
rect 1760 434 1768 442
rect 1780 434 1788 442
rect 1800 434 1808 442
rect 1820 434 1828 442
rect 1314 424 1322 432
rect 1334 424 1342 432
rect 1354 424 1362 432
rect 1374 424 1382 432
rect 1424 424 1432 432
rect 1444 424 1452 432
rect 1464 424 1472 432
rect 1484 424 1492 432
rect 1504 424 1512 432
rect 1620 424 1628 432
rect 1640 424 1648 432
rect 1660 424 1668 432
rect 1680 424 1688 432
rect 1730 424 1738 432
rect 1750 424 1758 432
rect 1770 424 1778 432
rect 1790 424 1798 432
rect 1810 424 1818 432
rect 1304 414 1312 422
rect 1324 414 1332 422
rect 1344 414 1352 422
rect 1364 414 1372 422
rect 1414 414 1422 422
rect 1434 414 1442 422
rect 1454 414 1462 422
rect 1474 414 1482 422
rect 1494 414 1502 422
rect 1610 414 1618 422
rect 1630 414 1638 422
rect 1650 414 1658 422
rect 1670 414 1678 422
rect 1720 414 1728 422
rect 1740 414 1748 422
rect 1760 414 1768 422
rect 1780 414 1788 422
rect 1800 414 1808 422
rect 1294 404 1302 412
rect 1314 404 1322 412
rect 1334 404 1342 412
rect 1354 404 1362 412
rect 1404 404 1412 412
rect 1424 404 1432 412
rect 1444 404 1452 412
rect 1464 404 1472 412
rect 1484 404 1492 412
rect 1600 404 1608 412
rect 1620 404 1628 412
rect 1640 404 1648 412
rect 1660 404 1668 412
rect 1710 404 1718 412
rect 1730 404 1738 412
rect 1750 404 1758 412
rect 1770 404 1778 412
rect 1790 404 1798 412
rect 1284 394 1292 402
rect 1304 394 1312 402
rect 1324 394 1332 402
rect 1344 394 1352 402
rect 1394 394 1402 402
rect 1414 394 1422 402
rect 1434 394 1442 402
rect 1454 394 1462 402
rect 1474 394 1482 402
rect 1590 394 1598 402
rect 1610 394 1618 402
rect 1630 394 1638 402
rect 1650 394 1658 402
rect 1700 394 1708 402
rect 1720 394 1728 402
rect 1740 394 1748 402
rect 1760 394 1768 402
rect 1780 394 1788 402
rect 1274 384 1282 392
rect 1294 384 1302 392
rect 1314 384 1322 392
rect 1334 384 1342 392
rect 1384 384 1392 392
rect 1404 384 1412 392
rect 1424 384 1432 392
rect 1444 384 1452 392
rect 1464 384 1472 392
rect 1580 384 1588 392
rect 1600 384 1608 392
rect 1620 384 1628 392
rect 1640 384 1648 392
rect 1690 384 1698 392
rect 1710 384 1718 392
rect 1730 384 1738 392
rect 1750 384 1758 392
rect 1770 384 1778 392
rect 1264 374 1272 382
rect 1284 374 1292 382
rect 1304 374 1312 382
rect 1324 374 1332 382
rect 1374 374 1382 382
rect 1394 374 1402 382
rect 1414 374 1422 382
rect 1434 374 1442 382
rect 1454 374 1462 382
rect 1570 374 1578 382
rect 1590 374 1598 382
rect 1610 374 1618 382
rect 1630 374 1638 382
rect 1680 374 1688 382
rect 1700 374 1708 382
rect 1720 374 1728 382
rect 1740 374 1748 382
rect 1760 374 1768 382
rect 1254 364 1262 372
rect 1274 364 1282 372
rect 1294 364 1302 372
rect 1314 364 1322 372
rect 1364 364 1372 372
rect 1384 364 1392 372
rect 1404 364 1412 372
rect 1424 364 1432 372
rect 1444 364 1452 372
rect 1560 364 1568 372
rect 1580 364 1588 372
rect 1600 364 1608 372
rect 1620 364 1628 372
rect 1670 364 1678 372
rect 1690 364 1698 372
rect 1710 364 1718 372
rect 1730 364 1738 372
rect 1750 364 1758 372
rect 1244 354 1252 362
rect 1264 354 1272 362
rect 1284 354 1292 362
rect 1304 354 1312 362
rect 1354 354 1362 362
rect 1374 354 1382 362
rect 1394 354 1402 362
rect 1414 354 1422 362
rect 1434 354 1442 362
rect 1550 354 1558 362
rect 1570 354 1578 362
rect 1590 354 1598 362
rect 1610 354 1618 362
rect 1660 354 1668 362
rect 1680 354 1688 362
rect 1700 354 1708 362
rect 1720 354 1728 362
rect 1740 354 1748 362
rect 1234 344 1242 352
rect 1254 344 1262 352
rect 1274 344 1282 352
rect 1294 344 1302 352
rect 1344 344 1352 352
rect 1364 344 1372 352
rect 1384 344 1392 352
rect 1404 344 1412 352
rect 1424 344 1432 352
rect 1540 344 1548 352
rect 1560 344 1568 352
rect 1580 344 1588 352
rect 1600 344 1608 352
rect 1650 344 1658 352
rect 1670 344 1678 352
rect 1690 344 1698 352
rect 1710 344 1718 352
rect 1730 344 1738 352
rect 1224 334 1232 342
rect 1244 334 1252 342
rect 1264 334 1272 342
rect 1284 334 1292 342
rect 1334 334 1342 342
rect 1354 334 1362 342
rect 1374 334 1382 342
rect 1394 334 1402 342
rect 1414 334 1422 342
rect 1530 334 1538 342
rect 1550 334 1558 342
rect 1570 334 1578 342
rect 1590 334 1598 342
rect 1640 334 1648 342
rect 1660 334 1668 342
rect 1680 334 1688 342
rect 1700 334 1708 342
rect 1720 334 1728 342
rect 1214 324 1222 332
rect 1234 324 1242 332
rect 1254 324 1262 332
rect 1274 324 1282 332
rect 1324 324 1332 332
rect 1344 324 1352 332
rect 1364 324 1372 332
rect 1384 324 1392 332
rect 1404 324 1412 332
rect 1520 324 1528 332
rect 1540 324 1548 332
rect 1560 324 1568 332
rect 1580 324 1588 332
rect 1630 324 1638 332
rect 1650 324 1658 332
rect 1670 324 1678 332
rect 1690 324 1698 332
rect 1710 324 1718 332
rect 1204 314 1212 322
rect 1224 314 1232 322
rect 1244 314 1252 322
rect 1264 314 1272 322
rect 1314 314 1322 322
rect 1334 314 1342 322
rect 1354 314 1362 322
rect 1374 314 1382 322
rect 1394 314 1402 322
rect 1510 314 1518 322
rect 1530 314 1538 322
rect 1550 314 1558 322
rect 1570 314 1578 322
rect 1620 314 1628 322
rect 1640 314 1648 322
rect 1660 314 1668 322
rect 1680 314 1688 322
rect 1700 314 1708 322
rect 1194 304 1202 312
rect 1214 304 1222 312
rect 1234 304 1242 312
rect 1254 304 1262 312
rect 1304 304 1312 312
rect 1324 304 1332 312
rect 1344 304 1352 312
rect 1364 304 1372 312
rect 1384 304 1392 312
rect 1500 304 1508 312
rect 1520 304 1528 312
rect 1540 304 1548 312
rect 1560 304 1568 312
rect 1610 304 1618 312
rect 1630 304 1638 312
rect 1650 304 1658 312
rect 1670 304 1678 312
rect 1690 304 1698 312
rect 1184 294 1192 302
rect 1204 294 1212 302
rect 1224 294 1232 302
rect 1244 294 1252 302
rect 1294 294 1302 302
rect 1314 294 1322 302
rect 1334 294 1342 302
rect 1354 294 1362 302
rect 1374 294 1382 302
rect 1490 294 1498 302
rect 1510 294 1518 302
rect 1530 294 1538 302
rect 1550 294 1558 302
rect 1600 294 1608 302
rect 1620 294 1628 302
rect 1640 294 1648 302
rect 1660 294 1668 302
rect 1680 294 1688 302
rect 1174 284 1182 292
rect 1194 284 1202 292
rect 1214 284 1222 292
rect 1234 284 1242 292
rect 1284 284 1292 292
rect 1304 284 1312 292
rect 1324 284 1332 292
rect 1344 284 1352 292
rect 1364 284 1372 292
rect 1480 284 1488 292
rect 1500 284 1508 292
rect 1520 284 1528 292
rect 1540 284 1548 292
rect 1590 284 1598 292
rect 1610 284 1618 292
rect 1630 284 1638 292
rect 1650 284 1658 292
rect 1670 284 1678 292
rect 1164 274 1172 282
rect 1184 274 1192 282
rect 1204 274 1212 282
rect 1224 274 1232 282
rect 1274 274 1282 282
rect 1294 274 1302 282
rect 1314 274 1322 282
rect 1334 274 1342 282
rect 1354 274 1362 282
rect 1470 274 1478 282
rect 1490 274 1498 282
rect 1510 274 1518 282
rect 1530 274 1538 282
rect 1580 274 1588 282
rect 1600 274 1608 282
rect 1620 274 1628 282
rect 1640 274 1648 282
rect 1660 274 1668 282
rect 1154 244 1162 272
rect 1174 244 1182 272
rect 1194 264 1202 272
rect 1214 264 1222 272
rect 1204 244 1212 262
rect 1234 244 1242 262
rect 1264 244 1272 272
rect 1284 264 1292 272
rect 1304 264 1312 272
rect 1294 244 1302 262
rect 1324 244 1332 272
rect 1344 264 1352 272
rect 1460 264 1468 272
rect 1480 264 1488 272
rect 1500 264 1508 272
rect 1520 264 1528 272
rect 1570 264 1578 272
rect 1590 264 1598 272
rect 1610 264 1618 272
rect 1630 264 1638 272
rect 1650 264 1658 272
rect 1450 254 1458 262
rect 1470 254 1478 262
rect 1490 254 1498 262
rect 1510 254 1518 262
rect 1560 254 1568 262
rect 1580 254 1588 262
rect 1600 254 1608 262
rect 1620 254 1628 262
rect 1640 254 1648 262
rect 1440 244 1448 252
rect 1460 244 1468 252
rect 1480 244 1488 252
rect 1500 244 1508 252
rect 1550 244 1558 252
rect 1570 244 1578 252
rect 1590 244 1598 252
rect 1610 244 1618 252
rect 1630 244 1638 252
rect 1164 234 1172 242
rect 1194 234 1202 242
rect 1224 234 1232 242
rect 1254 234 1262 242
rect 1284 234 1292 242
rect 1314 234 1322 242
rect 1430 234 1438 242
rect 1450 234 1458 242
rect 1470 234 1478 242
rect 1490 234 1498 242
rect 1540 234 1548 242
rect 1560 234 1568 242
rect 1580 234 1588 242
rect 1600 234 1608 242
rect 1620 234 1628 242
rect 1174 224 1182 232
rect 1204 224 1212 232
rect 1234 224 1242 232
rect 1264 224 1272 232
rect 1294 224 1302 232
rect 1420 224 1428 232
rect 1440 224 1448 232
rect 1460 224 1468 232
rect 1480 224 1488 232
rect 1530 224 1538 232
rect 1550 224 1558 232
rect 1570 224 1578 232
rect 1590 224 1598 232
rect 1610 224 1618 232
rect 1164 214 1172 222
rect 1194 214 1202 222
rect 1224 214 1232 222
rect 1254 214 1262 222
rect 1284 214 1292 222
rect 1410 214 1418 222
rect 1430 214 1438 222
rect 1450 214 1458 222
rect 1470 214 1478 222
rect 1520 214 1528 222
rect 1540 214 1548 222
rect 1560 214 1568 222
rect 1580 214 1588 222
rect 1600 214 1608 222
rect 1174 204 1182 212
rect 1204 204 1212 212
rect 1234 204 1242 212
rect 1264 204 1272 212
rect 1294 204 1302 212
rect 1400 204 1408 212
rect 1420 204 1428 212
rect 1440 204 1448 212
rect 1460 204 1468 212
rect 1510 204 1518 212
rect 1530 204 1538 212
rect 1550 204 1558 212
rect 1570 204 1578 212
rect 1590 204 1598 212
rect 1164 194 1172 202
rect 1194 194 1202 202
rect 1224 194 1232 202
rect 1254 194 1262 202
rect 1284 194 1292 202
rect 1390 194 1398 202
rect 1410 194 1418 202
rect 1430 194 1438 202
rect 1450 194 1458 202
rect 1500 194 1508 202
rect 1520 194 1528 202
rect 1540 194 1548 202
rect 1560 194 1568 202
rect 1580 194 1588 202
rect 1174 184 1182 192
rect 1204 184 1212 192
rect 1234 184 1242 192
rect 1264 184 1272 192
rect 1294 184 1302 192
rect 1380 184 1388 192
rect 1400 184 1408 192
rect 1420 184 1428 192
rect 1440 184 1448 192
rect 1490 184 1498 192
rect 1510 184 1518 192
rect 1530 184 1538 192
rect 1550 184 1558 192
rect 1570 184 1578 192
rect 1164 174 1172 182
rect 1194 174 1202 182
rect 1224 174 1232 182
rect 1254 174 1262 182
rect 1284 174 1292 182
rect 1174 164 1182 172
rect 1204 164 1212 172
rect 1234 164 1242 172
rect 1264 164 1272 172
rect 1294 164 1302 172
rect 1164 154 1172 162
rect 1194 154 1202 162
rect 1224 154 1232 162
rect 1254 154 1262 162
rect 1284 154 1292 162
rect 1174 144 1182 152
rect 1204 144 1212 152
rect 1234 144 1242 152
rect 1264 144 1272 152
rect 1294 144 1302 152
rect 1164 134 1172 142
rect 1194 134 1202 142
rect 1224 134 1232 142
rect 1254 134 1262 142
rect 1284 134 1292 142
rect 1174 124 1182 132
rect 1204 124 1212 132
rect 1234 124 1242 132
rect 1264 124 1272 132
rect 1294 124 1302 132
rect 1164 114 1172 122
rect 1194 114 1202 122
rect 1224 114 1232 122
rect 1254 114 1262 122
rect 1284 114 1292 122
rect 1174 104 1182 112
rect 1204 104 1212 112
rect 1234 104 1242 112
rect 1264 104 1272 112
rect 1294 104 1302 112
rect 1164 94 1172 102
rect 1194 94 1202 102
rect 1224 94 1232 102
rect 1254 94 1262 102
rect 1284 94 1292 102
rect 1174 84 1182 92
rect 1204 84 1212 92
rect 1234 84 1242 92
rect 1264 84 1272 92
rect 1294 84 1302 92
rect 1164 74 1172 82
rect 1194 74 1202 82
rect 1224 74 1232 82
rect 1254 74 1262 82
rect 1284 74 1292 82
rect 1174 64 1182 72
rect 1204 64 1212 72
rect 1234 64 1242 72
rect 1264 64 1272 72
rect 1294 64 1302 72
rect 1164 54 1172 62
rect 1194 54 1202 62
rect 1224 54 1232 62
rect 1254 54 1262 62
rect 1284 54 1292 62
rect 1174 44 1182 52
rect 1204 44 1212 52
rect 1234 44 1242 52
rect 1264 44 1272 52
rect 1294 44 1302 52
rect 1164 34 1172 42
rect 1194 34 1202 42
rect 1224 34 1232 42
rect 1254 34 1262 42
rect 1284 34 1292 42
rect 1174 24 1182 32
rect 1204 24 1212 32
rect 1234 24 1242 32
rect 1264 24 1272 32
rect 1294 24 1302 32
rect 1164 14 1172 22
rect 1194 14 1202 22
rect 1224 14 1232 22
rect 1254 14 1262 22
rect 1284 14 1292 22
rect 1174 4 1182 12
rect 1204 4 1212 12
rect 1234 4 1242 12
rect 1264 4 1272 12
rect 1294 4 1302 12
rect 1360 144 1368 172
rect 1380 144 1388 172
rect 1370 134 1378 142
rect 1400 134 1408 172
rect 1420 144 1428 172
rect 1470 144 1478 172
rect 1430 134 1438 142
rect 1460 134 1468 142
rect 1490 134 1498 172
rect 1510 144 1518 172
rect 1530 144 1538 172
rect 1550 164 1558 172
rect 1360 124 1368 132
rect 1390 124 1398 132
rect 1420 124 1428 132
rect 1450 124 1458 132
rect 1480 124 1488 132
rect 1370 114 1378 122
rect 1400 114 1408 122
rect 1430 114 1438 122
rect 1460 114 1468 122
rect 1490 114 1498 122
rect 1360 104 1368 112
rect 1390 104 1398 112
rect 1420 104 1428 112
rect 1450 104 1458 112
rect 1480 104 1488 112
rect 1370 94 1378 102
rect 1400 94 1408 102
rect 1430 94 1438 102
rect 1460 94 1468 102
rect 1490 94 1498 102
rect 1360 84 1368 92
rect 1390 84 1398 92
rect 1420 84 1428 92
rect 1450 84 1458 92
rect 1480 84 1488 92
rect 1370 74 1378 82
rect 1400 74 1408 82
rect 1430 74 1438 82
rect 1460 74 1468 82
rect 1490 74 1498 82
rect 1360 64 1368 72
rect 1390 64 1398 72
rect 1420 64 1428 72
rect 1450 64 1458 72
rect 1480 64 1488 72
rect 1370 54 1378 62
rect 1400 54 1408 62
rect 1430 54 1438 62
rect 1460 54 1468 62
rect 1490 54 1498 62
rect 1360 44 1368 52
rect 1390 44 1398 52
rect 1420 44 1428 52
rect 1450 44 1458 52
rect 1480 44 1488 52
rect 1370 34 1378 42
rect 1400 34 1408 42
rect 1430 34 1438 42
rect 1460 34 1468 42
rect 1490 34 1498 42
rect 1360 24 1368 32
rect 1390 24 1398 32
rect 1420 24 1428 32
rect 1450 24 1458 32
rect 1480 24 1488 32
rect 1370 14 1378 22
rect 1400 14 1408 22
rect 1430 14 1438 22
rect 1460 14 1468 22
rect 1490 14 1498 22
rect 1360 4 1368 12
rect 1390 4 1398 12
rect 1420 4 1428 12
rect 1450 4 1458 12
rect 1480 4 1488 12
<< metal2 >>
tri 1496 1252 1584 1340 se
rect 1584 1252 2000 1340
tri 1332 1088 1496 1252 se
rect 1496 1190 2000 1252
rect 1496 1180 1740 1190
rect 1958 1180 2000 1190
rect 1496 1088 2000 1180
tri 1158 914 1332 1088 se
rect 1332 1078 2000 1088
rect 1332 1070 1488 1078
tri 1488 1070 1496 1078 nw
tri 1496 1070 1504 1078 ne
rect 1332 1054 1472 1070
tri 1472 1054 1488 1070 nw
tri 1488 1054 1504 1070 se
rect 1504 1054 2000 1078
rect 1332 1038 1456 1054
tri 1456 1038 1472 1054 nw
tri 1472 1038 1488 1054 se
rect 1488 1040 2000 1054
rect 1488 1038 1740 1040
rect 1332 1022 1440 1038
tri 1440 1022 1456 1038 nw
tri 1456 1022 1472 1038 se
rect 1472 1030 1740 1038
rect 1958 1030 2000 1040
rect 1472 1022 2000 1030
rect 1332 1006 1424 1022
tri 1424 1006 1440 1022 nw
tri 1440 1006 1456 1022 se
rect 1456 1006 2000 1022
rect 1332 990 1408 1006
tri 1408 990 1424 1006 nw
tri 1424 990 1440 1006 se
rect 1440 990 2000 1006
rect 1332 978 1396 990
tri 1396 978 1408 990 nw
tri 1412 978 1424 990 se
rect 1424 978 2000 990
rect 1332 962 1380 978
tri 1380 962 1396 978 nw
tri 1396 962 1412 978 se
rect 1412 962 2000 978
rect 1332 946 1364 962
tri 1364 946 1380 962 nw
tri 1380 946 1396 962 se
rect 1396 961 2000 962
rect 1396 953 1583 961
tri 1583 953 1591 961 nw
tri 1591 953 1599 961 ne
rect 1396 946 1567 953
rect 1332 930 1348 946
tri 1348 930 1364 946 nw
tri 1364 930 1380 946 se
rect 1380 937 1567 946
tri 1567 937 1583 953 nw
tri 1583 937 1599 953 se
rect 1599 937 2000 961
rect 1380 930 1551 937
tri 1332 914 1348 930 nw
tri 1348 914 1364 930 se
rect 1364 921 1551 930
tri 1551 921 1567 937 nw
tri 1567 921 1583 937 se
rect 1583 921 2000 937
rect 1364 914 1544 921
tri 1544 914 1551 921 nw
tri 1560 914 1567 921 se
rect 1567 914 2000 921
tri 1092 848 1158 914 se
rect 1158 898 1316 914
tri 1316 898 1332 914 nw
tri 1332 898 1348 914 se
rect 1348 898 1528 914
tri 1528 898 1544 914 nw
tri 1544 898 1560 914 se
rect 1560 898 2000 914
rect 1158 882 1300 898
tri 1300 882 1316 898 nw
tri 1316 882 1332 898 se
rect 1332 882 1512 898
tri 1512 882 1528 898 nw
tri 1528 882 1544 898 se
rect 1544 882 2000 898
rect 1158 866 1284 882
tri 1284 866 1300 882 nw
tri 1300 866 1316 882 se
rect 1316 874 1504 882
tri 1504 874 1512 882 nw
tri 1520 874 1528 882 se
rect 1528 880 2000 882
rect 1528 874 1671 880
rect 1316 866 1488 874
rect 1158 864 1282 866
tri 1282 864 1284 866 nw
tri 1298 864 1300 866 se
rect 1300 864 1488 866
rect 1158 848 1266 864
tri 1266 848 1282 864 nw
tri 1282 848 1298 864 se
rect 1298 858 1488 864
tri 1488 858 1504 874 nw
tri 1504 858 1520 874 se
rect 1520 858 1671 874
tri 1671 858 1693 880 nw
rect 1298 853 1483 858
tri 1483 853 1488 858 nw
tri 1499 853 1504 858 se
rect 1504 853 1666 858
tri 1666 853 1671 858 nw
rect 1298 848 1478 853
tri 1478 848 1483 853 nw
tri 1494 848 1499 853 se
rect 1499 848 1661 853
tri 1661 848 1666 853 nw
tri 1086 842 1092 848 se
rect 1092 842 1260 848
tri 1260 842 1266 848 nw
tri 1276 842 1282 848 se
rect 1282 842 1472 848
tri 1472 842 1478 848 nw
tri 1488 842 1494 848 se
rect 1494 842 1655 848
tri 1655 842 1661 848 nw
tri 1716 842 1722 848 se
rect 1722 842 2000 848
tri 1078 834 1086 842 se
rect 1086 834 1252 842
tri 1252 834 1260 842 nw
tri 1268 834 1276 842 se
rect 1276 834 1464 842
tri 1464 834 1472 842 nw
tri 1480 834 1488 842 se
rect 1488 834 1647 842
tri 1647 834 1655 842 nw
tri 1708 834 1716 842 se
rect 1716 834 1724 842
rect 1732 834 1754 842
rect 1762 834 1784 842
rect 1792 834 1814 842
rect 1822 834 1844 842
rect 1852 834 1874 842
rect 1882 834 1904 842
rect 1912 834 1934 842
rect 1942 834 1964 842
rect 1972 834 2000 842
tri 1076 832 1078 834 se
rect 1078 832 1250 834
tri 1250 832 1252 834 nw
tri 1266 832 1268 834 se
rect 1268 832 1462 834
tri 1462 832 1464 834 nw
tri 1478 832 1480 834 se
rect 1480 832 1645 834
tri 1645 832 1647 834 nw
tri 1706 832 1708 834 se
rect 1708 832 2000 834
tri 1068 824 1076 832 se
rect 1076 824 1242 832
tri 1242 824 1250 832 nw
tri 1258 824 1266 832 se
rect 1266 824 1454 832
tri 1454 824 1462 832 nw
tri 1470 824 1478 832 se
rect 1478 824 1637 832
tri 1637 824 1645 832 nw
tri 1698 824 1706 832 se
rect 1706 824 1734 832
rect 1742 824 1764 832
rect 1772 824 1794 832
rect 1802 824 1824 832
rect 1832 824 1854 832
rect 1862 824 1884 832
rect 1892 824 1914 832
rect 1922 824 1944 832
rect 1952 824 1974 832
rect 1982 824 2000 832
tri 1066 822 1068 824 se
rect 1068 822 1240 824
tri 1240 822 1242 824 nw
tri 1256 822 1258 824 se
rect 1258 822 1452 824
tri 1452 822 1454 824 nw
tri 1468 822 1470 824 se
rect 1470 822 1635 824
tri 1635 822 1637 824 nw
tri 1696 822 1698 824 se
rect 1698 822 2000 824
tri 1058 814 1066 822 se
rect 1066 814 1232 822
tri 1232 814 1240 822 nw
tri 1248 814 1256 822 se
rect 1256 814 1444 822
tri 1444 814 1452 822 nw
tri 1460 814 1468 822 se
rect 1468 819 1632 822
tri 1632 819 1635 822 nw
tri 1693 819 1696 822 se
rect 1696 819 1724 822
rect 1468 814 1627 819
tri 1627 814 1632 819 nw
tri 1688 814 1693 819 se
rect 1693 814 1724 819
rect 1732 814 1754 822
rect 1762 814 1784 822
rect 1792 814 1814 822
rect 1822 814 1844 822
rect 1852 814 1874 822
rect 1882 814 1904 822
rect 1912 814 1934 822
rect 1942 814 1964 822
rect 1972 814 2000 822
tri 1056 812 1058 814 se
rect 1058 812 1230 814
tri 1230 812 1232 814 nw
tri 1246 812 1248 814 se
rect 1248 812 1442 814
tri 1442 812 1444 814 nw
tri 1458 812 1460 814 se
rect 1460 812 1625 814
tri 1625 812 1627 814 nw
tri 1686 812 1688 814 se
rect 1688 812 2000 814
tri 1048 804 1056 812 se
rect 1056 804 1222 812
tri 1222 804 1230 812 nw
tri 1238 804 1246 812 se
rect 1246 804 1434 812
tri 1434 804 1442 812 nw
tri 1450 804 1458 812 se
rect 1458 804 1617 812
tri 1617 804 1625 812 nw
tri 1678 804 1686 812 se
rect 1686 804 1694 812
rect 1702 804 1734 812
rect 1742 804 1764 812
rect 1772 804 1794 812
rect 1802 804 1824 812
rect 1832 804 1854 812
rect 1862 804 1884 812
rect 1892 804 1914 812
rect 1922 804 1944 812
rect 1952 804 1974 812
rect 1982 804 2000 812
tri 1046 802 1048 804 se
rect 1048 802 1220 804
tri 1220 802 1222 804 nw
tri 1236 802 1238 804 se
rect 1238 802 1432 804
tri 1432 802 1434 804 nw
tri 1448 802 1450 804 se
rect 1450 802 1615 804
tri 1615 802 1617 804 nw
tri 1676 802 1678 804 se
rect 1678 802 2000 804
tri 1038 794 1046 802 se
rect 1046 794 1212 802
tri 1212 794 1220 802 nw
tri 1228 794 1236 802 se
rect 1236 794 1424 802
tri 1424 794 1432 802 nw
tri 1440 794 1448 802 se
rect 1448 794 1607 802
tri 1607 794 1615 802 nw
tri 1668 794 1676 802 se
rect 1676 794 1684 802
rect 1692 794 1724 802
rect 1732 794 1754 802
rect 1762 794 1784 802
rect 1792 794 1814 802
rect 1822 794 1844 802
rect 1852 794 1874 802
rect 1882 794 1904 802
rect 1912 794 1934 802
rect 1942 794 1964 802
rect 1972 794 2000 802
tri 1036 792 1038 794 se
rect 1038 792 1210 794
tri 1210 792 1212 794 nw
tri 1226 792 1228 794 se
rect 1228 792 1422 794
tri 1422 792 1424 794 nw
tri 1438 792 1440 794 se
rect 1440 792 1605 794
tri 1605 792 1607 794 nw
tri 1666 792 1668 794 se
rect 1668 792 2000 794
tri 1028 784 1036 792 se
rect 1036 784 1202 792
tri 1202 784 1210 792 nw
tri 1218 784 1226 792 se
rect 1226 784 1414 792
tri 1414 784 1422 792 nw
tri 1430 784 1438 792 se
rect 1438 786 1599 792
tri 1599 786 1605 792 nw
tri 1660 786 1666 792 se
rect 1666 786 1674 792
rect 1438 784 1597 786
tri 1597 784 1599 786 nw
tri 1658 784 1660 786 se
rect 1660 784 1674 786
rect 1682 784 1694 792
rect 1702 784 1734 792
rect 1742 784 1764 792
rect 1772 784 1794 792
rect 1802 784 1824 792
rect 1832 784 1854 792
rect 1862 784 1884 792
rect 1892 784 1914 792
rect 1922 784 1944 792
rect 1952 784 1974 792
rect 1982 784 2000 792
tri 1026 782 1028 784 se
rect 1028 782 1200 784
tri 1200 782 1202 784 nw
tri 1216 782 1218 784 se
rect 1218 782 1412 784
tri 1412 782 1414 784 nw
tri 1428 782 1430 784 se
rect 1430 782 1595 784
tri 1595 782 1597 784 nw
tri 1656 782 1658 784 se
rect 1658 782 2000 784
tri 1018 774 1026 782 se
rect 1026 774 1192 782
tri 1192 774 1200 782 nw
tri 1208 774 1216 782 se
rect 1216 774 1404 782
tri 1404 774 1412 782 nw
tri 1420 774 1428 782 se
rect 1428 774 1587 782
tri 1587 774 1595 782 nw
tri 1648 774 1656 782 se
rect 1656 774 1664 782
rect 1672 774 1684 782
rect 1692 774 1724 782
rect 1732 774 1754 782
rect 1762 774 1784 782
rect 1792 774 1814 782
rect 1822 774 1844 782
rect 1852 774 1874 782
rect 1882 774 1904 782
rect 1912 774 1934 782
rect 1942 774 1964 782
rect 1972 774 2000 782
tri 1016 772 1018 774 se
rect 1018 772 1190 774
tri 1190 772 1192 774 nw
tri 1206 772 1208 774 se
rect 1208 772 1402 774
tri 1402 772 1404 774 nw
tri 1418 772 1420 774 se
rect 1420 772 1585 774
tri 1585 772 1587 774 nw
tri 1646 772 1648 774 se
rect 1648 772 2000 774
tri 1008 764 1016 772 se
rect 1016 764 1182 772
tri 1182 764 1190 772 nw
tri 1198 764 1206 772 se
rect 1206 764 1394 772
tri 1394 764 1402 772 nw
tri 1410 764 1418 772 se
rect 1418 764 1577 772
tri 1577 764 1585 772 nw
tri 1638 764 1646 772 se
rect 1646 764 1654 772
rect 1662 764 1674 772
rect 1682 764 1734 772
rect 1742 764 1764 772
rect 1772 764 1794 772
rect 1802 764 1824 772
rect 1832 764 1854 772
rect 1862 764 1884 772
rect 1892 764 1914 772
rect 1922 764 1944 772
rect 1952 764 1974 772
rect 1982 764 2000 772
tri 1006 762 1008 764 se
rect 1008 762 1180 764
tri 1180 762 1182 764 nw
tri 1196 762 1198 764 se
rect 1198 762 1392 764
tri 1392 762 1394 764 nw
tri 1408 762 1410 764 se
rect 1410 762 1575 764
tri 1575 762 1577 764 nw
tri 1636 762 1638 764 se
rect 1638 762 2000 764
tri 998 754 1006 762 se
rect 1006 754 1172 762
tri 1172 754 1180 762 nw
tri 1188 754 1196 762 se
rect 1196 754 1384 762
tri 1384 754 1392 762 nw
tri 1400 754 1408 762 se
rect 1408 754 1567 762
tri 1567 754 1575 762 nw
tri 1628 754 1636 762 se
rect 1636 754 1644 762
rect 1652 754 1664 762
rect 1672 754 1694 762
rect 1702 754 1724 762
rect 1732 754 1754 762
rect 1762 754 1784 762
rect 1792 754 1814 762
rect 1822 754 1844 762
rect 1852 754 1874 762
rect 1882 754 1904 762
rect 1912 754 1934 762
rect 1942 754 1964 762
rect 1972 754 2000 762
tri 996 752 998 754 se
rect 998 752 1170 754
tri 1170 752 1172 754 nw
tri 1186 752 1188 754 se
rect 1188 752 1382 754
tri 1382 752 1384 754 nw
tri 1398 752 1400 754 se
rect 1400 752 1565 754
tri 1565 752 1567 754 nw
tri 1626 752 1628 754 se
rect 1628 752 2000 754
tri 988 744 996 752 se
rect 996 744 1162 752
tri 1162 744 1170 752 nw
tri 1178 744 1186 752 se
rect 1186 744 1374 752
tri 1374 744 1382 752 nw
tri 1390 744 1398 752 se
rect 1398 744 1557 752
tri 1557 744 1565 752 nw
tri 1618 744 1626 752 se
rect 1626 744 1634 752
rect 1642 744 1654 752
rect 1662 744 1684 752
rect 1692 744 1734 752
rect 1742 744 1764 752
rect 1772 744 1794 752
rect 1802 744 1824 752
rect 1832 744 1854 752
rect 1862 744 1884 752
rect 1892 744 1914 752
rect 1922 744 1944 752
rect 1952 744 1974 752
rect 1982 744 2000 752
tri 986 742 988 744 se
rect 988 742 1160 744
tri 1160 742 1162 744 nw
tri 1176 742 1178 744 se
rect 1178 742 1372 744
tri 1372 742 1374 744 nw
tri 1388 742 1390 744 se
rect 1390 742 1555 744
tri 1555 742 1557 744 nw
tri 1616 742 1618 744 se
rect 1618 742 2000 744
tri 984 740 986 742 se
rect 986 740 1158 742
tri 1158 740 1160 742 nw
tri 1174 740 1176 742 se
rect 1176 740 1364 742
tri 978 734 984 740 se
rect 984 734 1152 740
tri 1152 734 1158 740 nw
tri 1168 734 1174 740 se
rect 1174 734 1364 740
tri 1364 734 1372 742 nw
tri 1380 734 1388 742 se
rect 1388 734 1547 742
tri 1547 734 1555 742 nw
tri 1608 734 1616 742 se
rect 1616 734 1624 742
rect 1632 734 1644 742
rect 1652 734 1674 742
rect 1682 738 1724 742
rect 1682 734 1704 738
tri 1704 734 1708 738 nw
tri 1708 734 1712 738 ne
rect 1712 734 1724 738
rect 1732 734 1754 742
rect 1762 734 1784 742
rect 1792 734 1814 742
rect 1822 734 1844 742
rect 1852 734 1874 742
rect 1882 734 1904 742
rect 1912 734 1934 742
rect 1942 734 1964 742
rect 1972 734 2000 742
tri 976 732 978 734 se
rect 978 732 1150 734
tri 1150 732 1152 734 nw
tri 1166 732 1168 734 se
rect 1168 732 1362 734
tri 1362 732 1364 734 nw
tri 1378 732 1380 734 se
rect 1380 732 1545 734
tri 1545 732 1547 734 nw
tri 1606 732 1608 734 se
rect 1608 732 1702 734
tri 1702 732 1704 734 nw
tri 1712 732 1714 734 ne
rect 1714 732 2000 734
tri 968 724 976 732 se
rect 976 724 1142 732
tri 1142 724 1150 732 nw
tri 1158 724 1166 732 se
rect 1166 724 1354 732
tri 1354 724 1362 732 nw
tri 1370 724 1378 732 se
rect 1378 725 1538 732
tri 1538 725 1545 732 nw
tri 1599 725 1606 732 se
rect 1606 725 1614 732
rect 1378 724 1537 725
tri 1537 724 1538 725 nw
tri 1598 724 1599 725 se
rect 1599 724 1614 725
rect 1622 724 1634 732
rect 1642 724 1664 732
rect 1672 728 1698 732
tri 1698 728 1702 732 nw
tri 1714 728 1718 732 ne
rect 1672 724 1694 728
tri 1694 724 1698 728 nw
tri 1714 724 1718 728 se
rect 1718 724 1734 732
rect 1742 724 1764 732
rect 1772 724 1794 732
rect 1802 724 1824 732
rect 1832 724 1854 732
rect 1862 724 1884 732
rect 1892 724 1914 732
rect 1922 724 1944 732
rect 1952 724 1974 732
rect 1982 724 2000 732
tri 966 722 968 724 se
rect 968 722 1140 724
tri 1140 722 1142 724 nw
tri 1156 722 1158 724 se
rect 1158 722 1352 724
tri 1352 722 1354 724 nw
tri 1368 722 1370 724 se
rect 1370 722 1535 724
tri 1535 722 1537 724 nw
tri 1596 722 1598 724 se
rect 1598 722 1692 724
tri 1692 722 1694 724 nw
tri 1712 722 1714 724 se
rect 1714 722 2000 724
tri 958 714 966 722 se
rect 966 714 1132 722
tri 1132 714 1140 722 nw
tri 1148 714 1156 722 se
rect 1156 714 1344 722
tri 1344 714 1352 722 nw
tri 1360 714 1368 722 se
rect 1368 714 1527 722
tri 1527 714 1535 722 nw
tri 1588 714 1596 722 se
rect 1596 714 1604 722
rect 1612 714 1624 722
rect 1632 714 1654 722
rect 1662 714 1684 722
tri 1684 714 1692 722 nw
tri 1704 714 1712 722 se
rect 1712 714 1724 722
rect 1732 714 1754 722
rect 1762 714 1784 722
rect 1792 714 1814 722
rect 1822 714 1844 722
rect 1852 714 1874 722
rect 1882 714 1904 722
rect 1912 714 1934 722
rect 1942 714 1964 722
rect 1972 714 2000 722
tri 956 712 958 714 se
rect 958 712 1130 714
tri 1130 712 1132 714 nw
tri 1146 712 1148 714 se
rect 1148 712 1342 714
tri 1342 712 1344 714 nw
tri 1358 712 1360 714 se
rect 1360 712 1525 714
tri 1525 712 1527 714 nw
tri 1586 712 1588 714 se
rect 1588 712 1682 714
tri 1682 712 1684 714 nw
tri 1702 712 1704 714 se
rect 1704 712 2000 714
tri 948 704 956 712 se
rect 956 704 1122 712
tri 1122 704 1130 712 nw
tri 1138 704 1146 712 se
rect 1146 704 1334 712
tri 1334 704 1342 712 nw
tri 1350 704 1358 712 se
rect 1358 704 1517 712
tri 1517 704 1525 712 nw
tri 1578 704 1586 712 se
rect 1586 704 1594 712
rect 1602 704 1614 712
rect 1622 704 1644 712
rect 1652 704 1674 712
tri 1674 704 1682 712 nw
tri 1694 704 1702 712 se
rect 1702 704 1734 712
rect 1742 704 1764 712
rect 1772 704 1794 712
rect 1802 704 1824 712
rect 1832 704 1854 712
rect 1862 704 1884 712
rect 1892 704 1914 712
rect 1922 704 1944 712
rect 1952 704 1974 712
rect 1982 704 2000 712
tri 946 702 948 704 se
rect 948 702 1120 704
tri 1120 702 1122 704 nw
tri 1136 702 1138 704 se
rect 1138 702 1332 704
tri 1332 702 1334 704 nw
tri 1348 702 1350 704 se
rect 1350 702 1515 704
tri 1515 702 1517 704 nw
tri 1576 702 1578 704 se
rect 1578 702 1672 704
tri 1672 702 1674 704 nw
tri 1692 702 1694 704 se
rect 1694 702 2000 704
tri 938 694 946 702 se
rect 946 694 1112 702
tri 1112 694 1120 702 nw
tri 1128 694 1136 702 se
rect 1136 694 1324 702
tri 1324 694 1332 702 nw
tri 1340 694 1348 702 se
rect 1348 694 1507 702
tri 1507 694 1515 702 nw
tri 1568 694 1576 702 se
rect 1576 694 1584 702
rect 1592 694 1604 702
rect 1612 694 1634 702
tri 936 692 938 694 se
rect 938 692 1110 694
tri 1110 692 1112 694 nw
tri 1126 692 1128 694 se
rect 1128 692 1322 694
tri 1322 692 1324 694 nw
tri 1338 692 1340 694 se
rect 1340 692 1505 694
tri 1505 692 1507 694 nw
tri 1566 692 1568 694 se
rect 1568 692 1634 694
tri 928 684 936 692 se
rect 936 684 1102 692
tri 1102 684 1110 692 nw
tri 1118 684 1126 692 se
rect 1126 684 1314 692
tri 1314 684 1322 692 nw
tri 1332 686 1338 692 se
rect 1338 686 1499 692
tri 1499 686 1505 692 nw
tri 1560 686 1566 692 se
rect 1566 686 1574 692
tri 1330 684 1332 686 se
rect 1332 684 1497 686
tri 1497 684 1499 686 nw
tri 1558 684 1560 686 se
rect 1560 684 1574 686
rect 1582 684 1594 692
rect 1602 684 1614 692
rect 1622 684 1634 692
rect 1642 694 1664 702
tri 1664 694 1672 702 nw
tri 1684 694 1692 702 se
rect 1692 694 1694 702
rect 1702 694 1724 702
rect 1642 692 1662 694
tri 1662 692 1664 694 nw
tri 1682 692 1684 694 se
rect 1684 692 1724 694
rect 1642 684 1654 692
tri 1654 684 1662 692 nw
tri 1674 684 1682 692 se
rect 1682 684 1684 692
rect 1692 684 1704 692
rect 1712 684 1724 692
rect 1732 694 1754 702
rect 1762 694 1784 702
rect 1792 694 1814 702
rect 1822 694 1844 702
rect 1852 694 1874 702
rect 1882 694 1904 702
rect 1912 694 1934 702
rect 1942 694 1964 702
rect 1972 694 2000 702
rect 1732 692 2000 694
rect 1732 684 1744 692
rect 1752 684 1764 692
rect 1772 688 2000 692
rect 1772 684 1784 688
tri 1784 684 1788 688 nw
tri 926 682 928 684 se
rect 928 682 1100 684
tri 1100 682 1102 684 nw
tri 1116 682 1118 684 se
rect 1118 682 1312 684
tri 1312 682 1314 684 nw
tri 1328 682 1330 684 se
rect 1330 682 1495 684
tri 1495 682 1497 684 nw
tri 1556 682 1558 684 se
rect 1558 682 1652 684
tri 1652 682 1654 684 nw
tri 1672 682 1674 684 se
rect 1674 682 1782 684
tri 1782 682 1784 684 nw
tri 922 678 926 682 se
rect 926 678 1096 682
tri 1096 678 1100 682 nw
tri 1112 678 1116 682 se
rect 1116 679 1309 682
tri 1309 679 1312 682 nw
tri 1325 679 1328 682 se
rect 1328 679 1492 682
tri 1492 679 1495 682 nw
tri 1553 679 1556 682 se
rect 1556 679 1564 682
rect 1116 678 1308 679
tri 1308 678 1309 679 nw
tri 1324 678 1325 679 se
rect 1325 678 1491 679
tri 1491 678 1492 679 nw
tri 1552 678 1553 679 se
rect 1553 678 1564 679
tri 918 674 922 678 se
rect 922 674 1092 678
tri 1092 674 1096 678 nw
tri 1108 674 1112 678 se
rect 1112 674 1304 678
tri 1304 674 1308 678 nw
tri 1320 674 1324 678 se
rect 1324 674 1487 678
tri 1487 674 1491 678 nw
tri 1548 674 1552 678 se
rect 1552 674 1564 678
rect 1572 674 1584 682
rect 1592 674 1604 682
rect 1612 674 1624 682
rect 1632 678 1648 682
tri 1648 678 1652 682 nw
tri 1668 678 1672 682 se
rect 1672 678 1674 682
rect 1632 674 1644 678
tri 1644 674 1648 678 nw
tri 1664 674 1668 678 se
rect 1668 674 1674 678
rect 1682 674 1694 682
rect 1702 674 1714 682
rect 1722 674 1734 682
rect 1742 674 1754 682
rect 1762 674 1774 682
tri 1774 674 1782 682 nw
tri 916 672 918 674 se
rect 918 672 1090 674
tri 1090 672 1092 674 nw
tri 1106 672 1108 674 se
rect 1108 672 1302 674
tri 1302 672 1304 674 nw
tri 1318 672 1320 674 se
rect 1320 672 1485 674
tri 1485 672 1487 674 nw
tri 1546 672 1548 674 se
rect 1548 672 1642 674
tri 1642 672 1644 674 nw
tri 1662 672 1664 674 se
rect 1664 672 1772 674
tri 1772 672 1774 674 nw
tri 908 664 916 672 se
rect 916 664 1082 672
tri 1082 664 1090 672 nw
tri 1098 664 1106 672 se
rect 1106 664 1294 672
tri 1294 664 1302 672 nw
tri 1310 664 1318 672 se
rect 1318 664 1477 672
tri 1477 664 1485 672 nw
tri 1538 664 1546 672 se
rect 1546 664 1554 672
rect 1562 664 1574 672
rect 1582 664 1594 672
rect 1602 664 1614 672
rect 1622 664 1634 672
tri 1634 664 1642 672 nw
tri 1654 664 1662 672 se
rect 1662 664 1664 672
rect 1672 664 1684 672
rect 1692 664 1704 672
rect 1712 664 1724 672
rect 1732 664 1744 672
rect 1752 664 1764 672
tri 1764 664 1772 672 nw
tri 906 662 908 664 se
rect 908 662 1080 664
tri 1080 662 1082 664 nw
tri 1096 662 1098 664 se
rect 1098 662 1292 664
tri 1292 662 1294 664 nw
tri 1308 662 1310 664 se
rect 1310 662 1475 664
tri 1475 662 1477 664 nw
tri 1536 662 1538 664 se
rect 1538 662 1632 664
tri 1632 662 1634 664 nw
tri 1652 662 1654 664 se
rect 1654 662 1762 664
tri 1762 662 1764 664 nw
tri 898 654 906 662 se
rect 906 654 1072 662
tri 1072 654 1080 662 nw
tri 1088 654 1096 662 se
rect 1096 654 1284 662
tri 1284 654 1292 662 nw
tri 1300 654 1308 662 se
rect 1308 654 1467 662
tri 1467 654 1475 662 nw
tri 1528 654 1536 662 se
rect 1536 654 1544 662
rect 1552 654 1564 662
rect 1572 654 1584 662
rect 1592 654 1604 662
rect 1612 658 1628 662
tri 1628 658 1632 662 nw
tri 1648 658 1652 662 se
rect 1652 658 1654 662
rect 1612 654 1624 658
tri 1624 654 1628 658 nw
tri 1644 654 1648 658 se
rect 1648 654 1654 658
rect 1662 654 1674 662
rect 1682 654 1694 662
rect 1702 654 1714 662
rect 1722 654 1734 662
rect 1742 654 1754 662
tri 1754 654 1762 662 nw
tri 896 652 898 654 se
rect 898 652 1070 654
tri 1070 652 1072 654 nw
tri 1086 652 1088 654 se
rect 1088 652 1282 654
tri 1282 652 1284 654 nw
tri 1298 652 1300 654 se
rect 1300 652 1465 654
tri 1465 652 1467 654 nw
tri 1526 652 1528 654 se
rect 1528 652 1622 654
tri 1622 652 1624 654 nw
tri 1642 652 1644 654 se
rect 1644 652 1752 654
tri 1752 652 1754 654 nw
tri 888 644 896 652 se
rect 896 644 1062 652
tri 1062 644 1070 652 nw
tri 1078 644 1086 652 se
rect 1086 644 1274 652
tri 1274 644 1282 652 nw
tri 1290 644 1298 652 se
rect 1298 644 1457 652
tri 1457 644 1465 652 nw
tri 1518 644 1526 652 se
rect 1526 644 1534 652
rect 1542 644 1554 652
rect 1562 644 1574 652
rect 1582 644 1594 652
rect 1602 644 1614 652
tri 1614 644 1622 652 nw
tri 1634 644 1642 652 se
rect 1642 644 1644 652
rect 1652 644 1664 652
rect 1672 644 1684 652
rect 1692 644 1704 652
rect 1712 644 1724 652
rect 1732 644 1744 652
tri 1744 644 1752 652 nw
tri 1814 644 1822 652 se
rect 1822 644 2000 652
tri 886 642 888 644 se
rect 888 642 1060 644
tri 1060 642 1062 644 nw
tri 1076 642 1078 644 se
rect 1078 642 1272 644
tri 1272 642 1274 644 nw
tri 1288 642 1290 644 se
rect 1290 642 1455 644
tri 1455 642 1457 644 nw
tri 1516 642 1518 644 se
rect 1518 642 1612 644
tri 1612 642 1614 644 nw
tri 1632 642 1634 644 se
rect 1634 642 1742 644
tri 1742 642 1744 644 nw
tri 1812 642 1814 644 se
rect 1814 642 2000 644
tri 878 634 886 642 se
rect 886 634 1052 642
tri 1052 634 1060 642 nw
tri 1068 634 1076 642 se
rect 1076 634 1264 642
tri 1264 634 1272 642 nw
tri 1280 634 1288 642 se
rect 1288 634 1447 642
tri 1447 634 1455 642 nw
tri 1508 634 1516 642 se
rect 1516 634 1524 642
rect 1532 634 1544 642
rect 1552 634 1564 642
rect 1572 634 1584 642
rect 1592 634 1604 642
tri 1604 634 1612 642 nw
tri 1624 634 1632 642 se
rect 1632 634 1634 642
rect 1642 634 1654 642
rect 1662 634 1674 642
rect 1682 634 1694 642
rect 1702 634 1714 642
rect 1722 634 1734 642
tri 1734 634 1742 642 nw
tri 1804 634 1812 642 se
rect 1812 634 1830 642
rect 1838 634 1860 642
rect 1868 634 1890 642
rect 1898 634 1920 642
rect 1928 634 1950 642
rect 1958 634 1980 642
rect 1988 634 2000 642
tri 876 632 878 634 se
rect 878 632 1050 634
tri 1050 632 1052 634 nw
tri 1066 632 1068 634 se
rect 1068 632 1262 634
tri 1262 632 1264 634 nw
tri 1278 632 1280 634 se
rect 1280 632 1445 634
tri 1445 632 1447 634 nw
tri 1506 632 1508 634 se
rect 1508 632 1602 634
tri 1602 632 1604 634 nw
tri 1622 632 1624 634 se
rect 1624 632 1732 634
tri 1732 632 1734 634 nw
tri 1802 632 1804 634 se
rect 1804 632 2000 634
tri 868 624 876 632 se
rect 876 624 1042 632
tri 1042 624 1050 632 nw
tri 1058 624 1066 632 se
rect 1066 624 1254 632
tri 1254 624 1262 632 nw
tri 1270 624 1278 632 se
rect 1278 625 1438 632
tri 1438 625 1445 632 nw
tri 1499 625 1506 632 se
rect 1506 625 1514 632
rect 1278 624 1437 625
tri 1437 624 1438 625 nw
tri 1498 624 1499 625 se
rect 1499 624 1514 625
rect 1522 624 1534 632
rect 1542 624 1554 632
rect 1562 624 1574 632
rect 1582 624 1594 632
tri 1594 624 1602 632 nw
tri 1614 624 1622 632 se
rect 1622 624 1624 632
rect 1632 624 1644 632
rect 1652 624 1664 632
rect 1672 624 1684 632
rect 1692 624 1704 632
rect 1712 624 1724 632
tri 1724 624 1732 632 nw
tri 1794 624 1802 632 se
rect 1802 624 1840 632
rect 1848 624 1870 632
rect 1878 624 1900 632
rect 1908 624 1930 632
rect 1938 624 1960 632
rect 1968 624 1990 632
rect 1998 624 2000 632
tri 866 622 868 624 se
rect 868 622 1040 624
tri 1040 622 1042 624 nw
tri 1056 622 1058 624 se
rect 1058 622 1252 624
tri 1252 622 1254 624 nw
tri 1268 622 1270 624 se
rect 1270 622 1435 624
tri 1435 622 1437 624 nw
tri 1496 622 1498 624 se
rect 1498 622 1592 624
tri 1592 622 1594 624 nw
tri 1612 622 1614 624 se
rect 1614 622 1722 624
tri 1722 622 1724 624 nw
tri 1792 622 1794 624 se
rect 1794 622 2000 624
tri 858 614 866 622 se
rect 866 614 1032 622
tri 1032 614 1040 622 nw
tri 1048 614 1056 622 se
rect 1056 614 1244 622
tri 1244 614 1252 622 nw
tri 1260 614 1268 622 se
rect 1268 614 1427 622
tri 1427 614 1435 622 nw
tri 1488 614 1496 622 se
rect 1496 614 1504 622
rect 1512 614 1524 622
rect 1532 614 1544 622
rect 1552 614 1564 622
rect 1572 614 1584 622
tri 1584 614 1592 622 nw
tri 1604 614 1612 622 se
rect 1612 614 1614 622
rect 1622 614 1634 622
rect 1642 614 1654 622
rect 1662 614 1674 622
rect 1682 614 1694 622
rect 1702 618 1718 622
tri 1718 618 1722 622 nw
tri 1788 618 1792 622 se
rect 1792 618 1830 622
rect 1702 614 1714 618
tri 1714 614 1718 618 nw
tri 1784 614 1788 618 se
rect 1788 614 1830 618
rect 1838 614 1860 622
rect 1868 614 1890 622
rect 1898 614 1920 622
rect 1928 614 1950 622
rect 1958 614 1980 622
rect 1988 614 2000 622
tri 856 612 858 614 se
rect 858 612 1030 614
tri 1030 612 1032 614 nw
tri 1046 612 1048 614 se
rect 1048 612 1242 614
tri 1242 612 1244 614 nw
tri 1258 612 1260 614 se
rect 1260 612 1425 614
tri 1425 612 1427 614 nw
tri 1486 612 1488 614 se
rect 1488 612 1582 614
tri 1582 612 1584 614 nw
tri 1602 612 1604 614 se
rect 1604 612 1712 614
tri 1712 612 1714 614 nw
tri 1782 612 1784 614 se
rect 1784 612 2000 614
tri 848 604 856 612 se
rect 856 604 1022 612
tri 1022 604 1030 612 nw
tri 1038 604 1046 612 se
rect 1046 604 1234 612
tri 1234 604 1242 612 nw
tri 1250 604 1258 612 se
rect 1258 604 1417 612
tri 1417 604 1425 612 nw
tri 1478 604 1486 612 se
rect 1486 604 1494 612
rect 1502 604 1514 612
rect 1522 604 1534 612
rect 1542 604 1554 612
rect 1562 604 1574 612
tri 1574 604 1582 612 nw
tri 1594 604 1602 612 se
rect 1602 604 1604 612
rect 1612 604 1624 612
rect 1632 604 1644 612
rect 1652 604 1664 612
rect 1672 604 1684 612
rect 1692 604 1704 612
tri 1704 604 1712 612 nw
tri 1774 604 1782 612 se
rect 1782 604 1810 612
rect 1818 604 1840 612
rect 1848 604 1870 612
rect 1878 604 1900 612
rect 1908 604 1930 612
rect 1938 604 1960 612
rect 1968 604 1990 612
rect 1998 604 2000 612
tri 846 602 848 604 se
rect 848 602 1020 604
tri 1020 602 1022 604 nw
tri 1036 602 1038 604 se
rect 1038 602 1232 604
tri 1232 602 1234 604 nw
tri 1248 602 1250 604 se
rect 1250 602 1415 604
tri 1415 602 1417 604 nw
tri 1476 602 1478 604 se
rect 1478 602 1572 604
tri 1572 602 1574 604 nw
tri 1592 602 1594 604 se
rect 1594 602 1702 604
tri 1702 602 1704 604 nw
tri 1772 602 1774 604 se
rect 1774 602 2000 604
tri 838 594 846 602 se
rect 846 594 1012 602
tri 1012 594 1020 602 nw
tri 1028 594 1036 602 se
rect 1036 594 1224 602
tri 1224 594 1232 602 nw
tri 1240 594 1248 602 se
rect 1248 594 1407 602
tri 1407 594 1415 602 nw
tri 1468 594 1476 602 se
rect 1476 594 1484 602
rect 1492 594 1504 602
rect 1512 594 1524 602
rect 1532 594 1544 602
rect 1552 594 1564 602
tri 1564 594 1572 602 nw
tri 1584 594 1592 602 se
rect 1592 594 1594 602
rect 1602 594 1614 602
rect 1622 594 1634 602
rect 1642 594 1654 602
rect 1662 594 1674 602
rect 1682 600 1700 602
tri 1700 600 1702 602 nw
tri 1770 600 1772 602 se
rect 1772 600 1800 602
rect 1682 594 1694 600
tri 1694 594 1700 600 nw
tri 1764 594 1770 600 se
rect 1770 594 1800 600
rect 1808 594 1830 602
rect 1838 594 1860 602
rect 1868 594 1890 602
rect 1898 594 1920 602
rect 1928 594 1950 602
rect 1958 594 1980 602
rect 1988 594 2000 602
tri 836 592 838 594 se
rect 838 592 1010 594
tri 1010 592 1012 594 nw
tri 1026 592 1028 594 se
rect 1028 592 1222 594
tri 1222 592 1224 594 nw
tri 1238 592 1240 594 se
rect 1240 592 1405 594
tri 1405 592 1407 594 nw
tri 1466 592 1468 594 se
rect 1468 592 1562 594
tri 1562 592 1564 594 nw
tri 1582 592 1584 594 se
rect 1584 592 1692 594
tri 1692 592 1694 594 nw
tri 1762 592 1764 594 se
rect 1764 592 2000 594
tri 828 584 836 592 se
rect 836 584 1002 592
tri 1002 584 1010 592 nw
tri 1018 584 1026 592 se
rect 1026 584 1214 592
tri 1214 584 1222 592 nw
tri 1230 584 1238 592 se
rect 1238 584 1397 592
tri 1397 584 1405 592 nw
tri 1458 584 1466 592 se
rect 1466 584 1474 592
rect 1482 584 1494 592
rect 1502 584 1514 592
rect 1522 584 1534 592
rect 1542 584 1554 592
tri 1554 584 1562 592 nw
tri 1574 584 1582 592 se
rect 1582 584 1584 592
rect 1592 584 1604 592
rect 1612 584 1624 592
rect 1632 584 1644 592
rect 1652 584 1664 592
rect 1672 584 1684 592
tri 1684 584 1692 592 nw
tri 1754 584 1762 592 se
rect 1762 584 1790 592
rect 1798 584 1840 592
rect 1848 584 1870 592
rect 1878 584 1900 592
rect 1908 584 1930 592
rect 1938 584 1960 592
rect 1968 584 1990 592
rect 1998 584 2000 592
tri 826 582 828 584 se
rect 828 582 1000 584
tri 1000 582 1002 584 nw
tri 1016 582 1018 584 se
rect 1018 582 1212 584
tri 1212 582 1214 584 nw
tri 1228 582 1230 584 se
rect 1230 582 1395 584
tri 1395 582 1397 584 nw
tri 1456 582 1458 584 se
rect 1458 582 1552 584
tri 1552 582 1554 584 nw
tri 1572 582 1574 584 se
rect 1574 582 1682 584
tri 1682 582 1684 584 nw
tri 1752 582 1754 584 se
rect 1754 582 1850 584
tri 1850 582 1852 584 nw
tri 1852 582 1854 584 ne
rect 1854 582 2000 584
tri 818 574 826 582 se
rect 826 574 992 582
tri 992 574 1000 582 nw
tri 1008 574 1016 582 se
rect 1016 574 1204 582
tri 1204 574 1212 582 nw
tri 1220 574 1228 582 se
rect 1228 574 1387 582
tri 1387 574 1395 582 nw
tri 1448 574 1456 582 se
rect 1456 574 1464 582
rect 1472 574 1484 582
rect 1492 574 1504 582
rect 1512 574 1524 582
rect 1532 574 1544 582
tri 1544 574 1552 582 nw
tri 1564 574 1572 582 se
rect 1572 574 1574 582
rect 1582 574 1594 582
rect 1602 574 1614 582
rect 1622 574 1634 582
rect 1642 574 1654 582
rect 1662 574 1674 582
tri 1674 574 1682 582 nw
tri 1744 574 1752 582 se
rect 1752 574 1780 582
rect 1788 574 1810 582
rect 1818 574 1830 582
rect 1838 576 1844 582
tri 1844 576 1850 582 nw
tri 1854 576 1860 582 ne
rect 1838 574 1842 576
tri 1842 574 1844 576 nw
tri 1858 574 1860 576 se
rect 1860 574 1890 582
rect 1898 574 1920 582
rect 1928 574 1950 582
rect 1958 574 1980 582
rect 1988 574 2000 582
tri 816 572 818 574 se
rect 818 572 990 574
tri 990 572 992 574 nw
tri 1006 572 1008 574 se
rect 1008 572 1202 574
tri 1202 572 1204 574 nw
tri 1218 572 1220 574 se
rect 1220 572 1385 574
tri 1385 572 1387 574 nw
tri 1446 572 1448 574 se
rect 1448 572 1542 574
tri 1542 572 1544 574 nw
tri 1562 572 1564 574 se
rect 1564 572 1672 574
tri 1672 572 1674 574 nw
tri 1742 572 1744 574 se
rect 1744 572 1840 574
tri 1840 572 1842 574 nw
tri 1856 572 1858 574 se
rect 1858 572 2000 574
tri 810 566 816 572 se
rect 816 566 984 572
tri 984 566 990 572 nw
tri 1000 566 1006 572 se
rect 1006 566 1194 572
tri 808 564 810 566 se
rect 810 564 982 566
tri 982 564 984 566 nw
tri 998 564 1000 566 se
rect 1000 564 1194 566
tri 1194 564 1202 572 nw
tri 1210 564 1218 572 se
rect 1218 564 1377 572
tri 1377 564 1385 572 nw
tri 1438 564 1446 572 se
rect 1446 564 1454 572
rect 1462 564 1474 572
rect 1482 564 1494 572
rect 1502 564 1514 572
rect 1522 564 1534 572
tri 1534 564 1542 572 nw
tri 1554 564 1562 572 se
rect 1562 564 1564 572
rect 1572 564 1584 572
rect 1592 564 1604 572
rect 1612 564 1624 572
rect 1632 564 1644 572
rect 1652 564 1664 572
tri 1664 564 1672 572 nw
tri 1734 564 1742 572 se
rect 1742 564 1770 572
rect 1778 564 1800 572
rect 1808 564 1832 572
tri 1832 564 1840 572 nw
tri 1848 564 1856 572 se
rect 1856 564 1870 572
rect 1878 564 1900 572
rect 1908 564 1930 572
rect 1938 564 1960 572
rect 1968 564 1990 572
rect 1998 564 2000 572
tri 806 562 808 564 se
rect 808 562 980 564
tri 980 562 982 564 nw
tri 996 562 998 564 se
rect 998 562 1192 564
tri 1192 562 1194 564 nw
tri 1208 562 1210 564 se
rect 1210 562 1375 564
tri 1375 562 1377 564 nw
tri 1436 562 1438 564 se
rect 1438 562 1532 564
tri 1532 562 1534 564 nw
tri 1552 562 1554 564 se
rect 1554 562 1662 564
tri 1662 562 1664 564 nw
tri 1732 562 1734 564 se
rect 1734 562 1830 564
tri 1830 562 1832 564 nw
tri 1846 562 1848 564 se
rect 1848 562 2000 564
tri 798 554 806 562 se
rect 806 554 972 562
tri 972 554 980 562 nw
tri 988 554 996 562 se
rect 996 554 1184 562
tri 1184 554 1192 562 nw
tri 1200 554 1208 562 se
rect 1208 554 1367 562
tri 1367 554 1375 562 nw
tri 1428 554 1436 562 se
rect 1436 554 1444 562
rect 1452 554 1464 562
rect 1472 554 1484 562
rect 1492 554 1504 562
rect 1512 554 1524 562
tri 1524 554 1532 562 nw
tri 1544 554 1552 562 se
rect 1552 554 1554 562
rect 1562 554 1574 562
rect 1582 554 1594 562
rect 1602 554 1614 562
rect 1622 554 1634 562
rect 1642 554 1654 562
tri 1654 554 1662 562 nw
tri 1724 554 1732 562 se
rect 1732 554 1760 562
rect 1768 554 1790 562
rect 1798 554 1822 562
tri 1822 554 1830 562 nw
tri 1838 554 1846 562 se
rect 1846 554 1860 562
rect 1868 554 1890 562
rect 1898 554 1920 562
rect 1928 554 1950 562
rect 1958 554 1980 562
rect 1988 554 2000 562
tri 796 552 798 554 se
rect 798 552 970 554
tri 970 552 972 554 nw
tri 986 552 988 554 se
rect 988 552 1182 554
tri 1182 552 1184 554 nw
tri 1198 552 1200 554 se
rect 1200 552 1365 554
tri 1365 552 1367 554 nw
tri 1426 552 1428 554 se
rect 1428 552 1522 554
tri 1522 552 1524 554 nw
tri 1542 552 1544 554 se
rect 1544 552 1652 554
tri 1652 552 1654 554 nw
tri 1722 552 1724 554 se
rect 1724 552 1820 554
tri 1820 552 1822 554 nw
tri 1836 552 1838 554 se
rect 1838 552 2000 554
tri 788 544 796 552 se
rect 796 550 968 552
tri 968 550 970 552 nw
tri 984 550 986 552 se
rect 986 550 1180 552
tri 1180 550 1182 552 nw
tri 1196 550 1198 552 se
rect 1198 550 1357 552
rect 796 544 962 550
tri 962 544 968 550 nw
tri 978 544 984 550 se
rect 984 544 1174 550
tri 1174 544 1180 550 nw
tri 1190 544 1196 550 se
rect 1196 544 1357 550
tri 1357 544 1365 552 nw
tri 1418 544 1426 552 se
rect 1426 544 1434 552
rect 1442 544 1454 552
rect 1462 544 1474 552
rect 1482 544 1494 552
rect 1502 544 1514 552
tri 1514 544 1522 552 nw
tri 1534 544 1542 552 se
rect 1542 544 1544 552
rect 1552 544 1564 552
rect 1572 544 1584 552
rect 1592 544 1604 552
rect 1612 544 1624 552
rect 1632 548 1648 552
tri 1648 548 1652 552 nw
tri 1718 548 1722 552 se
rect 1722 548 1750 552
rect 1632 544 1644 548
tri 1644 544 1648 548 nw
tri 1714 544 1718 548 se
rect 1718 544 1750 548
rect 1758 544 1780 552
rect 1788 544 1812 552
tri 1812 544 1820 552 nw
tri 1828 544 1836 552 se
rect 1836 544 1840 552
rect 1848 544 1870 552
rect 1878 544 1900 552
rect 1908 544 1930 552
rect 1938 544 1960 552
rect 1968 544 1990 552
rect 1998 544 2000 552
tri 786 542 788 544 se
rect 788 542 960 544
tri 960 542 962 544 nw
tri 976 542 978 544 se
rect 978 542 1172 544
tri 1172 542 1174 544 nw
tri 1188 542 1190 544 se
rect 1190 542 1355 544
tri 1355 542 1357 544 nw
tri 1416 542 1418 544 se
rect 1418 542 1512 544
tri 1512 542 1514 544 nw
tri 1532 542 1534 544 se
rect 1534 542 1642 544
tri 1642 542 1644 544 nw
tri 1712 542 1714 544 se
rect 1714 542 1810 544
tri 1810 542 1812 544 nw
tri 1826 542 1828 544 se
rect 1828 542 2000 544
tri 778 534 786 542 se
rect 786 534 952 542
tri 952 534 960 542 nw
tri 968 534 976 542 se
rect 976 534 1164 542
tri 1164 534 1172 542 nw
tri 1180 534 1188 542 se
rect 1188 534 1347 542
tri 1347 534 1355 542 nw
tri 1408 534 1416 542 se
rect 1416 534 1424 542
rect 1432 534 1444 542
rect 1452 534 1464 542
rect 1472 534 1484 542
rect 1492 534 1504 542
tri 1504 534 1512 542 nw
tri 1524 534 1532 542 se
rect 1532 534 1534 542
rect 1542 534 1554 542
rect 1562 534 1574 542
rect 1582 534 1594 542
rect 1602 534 1614 542
rect 1622 534 1634 542
tri 1634 534 1642 542 nw
tri 1704 534 1712 542 se
rect 1712 534 1740 542
rect 1748 534 1770 542
rect 1778 534 1802 542
tri 1802 534 1810 542 nw
tri 1818 534 1826 542 se
rect 1826 534 1830 542
rect 1838 534 1860 542
rect 1868 534 1890 542
rect 1898 534 1920 542
rect 1928 534 1950 542
rect 1958 534 1980 542
rect 1988 534 2000 542
tri 776 532 778 534 se
rect 778 532 950 534
tri 950 532 952 534 nw
tri 966 532 968 534 se
rect 968 532 1162 534
tri 1162 532 1164 534 nw
tri 1178 532 1180 534 se
rect 1180 532 1345 534
tri 1345 532 1347 534 nw
tri 1406 532 1408 534 se
rect 1408 532 1502 534
tri 1502 532 1504 534 nw
tri 1522 532 1524 534 se
rect 1524 532 1632 534
tri 1632 532 1634 534 nw
tri 1702 532 1704 534 se
rect 1704 532 1800 534
tri 1800 532 1802 534 nw
tri 1816 532 1818 534 se
rect 1818 532 2000 534
tri 768 524 776 532 se
rect 776 526 944 532
tri 944 526 950 532 nw
tri 960 526 966 532 se
rect 966 528 1158 532
tri 1158 528 1162 532 nw
tri 1174 528 1178 532 se
rect 1178 528 1337 532
rect 966 526 1156 528
tri 1156 526 1158 528 nw
tri 1172 526 1174 528 se
rect 1174 526 1337 528
rect 776 524 942 526
tri 942 524 944 526 nw
tri 958 524 960 526 se
rect 960 524 1154 526
tri 1154 524 1156 526 nw
tri 1170 524 1172 526 se
rect 1172 524 1337 526
tri 1337 524 1345 532 nw
tri 1398 524 1406 532 se
rect 1406 524 1414 532
rect 1422 524 1434 532
rect 1442 524 1454 532
rect 1462 524 1474 532
rect 1482 529 1499 532
tri 1499 529 1502 532 nw
tri 1519 529 1522 532 se
rect 1522 529 1524 532
rect 1482 524 1494 529
tri 1494 524 1499 529 nw
tri 1514 524 1519 529 se
rect 1519 524 1524 529
rect 1532 524 1544 532
rect 1552 524 1564 532
rect 1572 524 1584 532
rect 1592 524 1604 532
rect 1612 524 1624 532
tri 1624 524 1632 532 nw
tri 1694 524 1702 532 se
rect 1702 524 1730 532
rect 1738 524 1760 532
rect 1768 524 1792 532
tri 1792 524 1800 532 nw
tri 1808 524 1816 532 se
rect 1816 524 1840 532
rect 1848 524 1870 532
rect 1878 524 1900 532
rect 1908 524 1930 532
rect 1938 524 1960 532
rect 1968 524 1990 532
rect 1998 524 2000 532
tri 766 522 768 524 se
rect 768 522 940 524
tri 940 522 942 524 nw
tri 956 522 958 524 se
rect 958 522 1152 524
tri 1152 522 1154 524 nw
tri 1168 522 1170 524 se
rect 1170 522 1335 524
tri 1335 522 1337 524 nw
tri 1396 522 1398 524 se
rect 1398 522 1492 524
tri 1492 522 1494 524 nw
tri 1512 522 1514 524 se
rect 1514 522 1622 524
tri 1622 522 1624 524 nw
tri 1692 522 1694 524 se
rect 1694 522 1790 524
tri 1790 522 1792 524 nw
tri 1806 522 1808 524 se
rect 1808 522 2000 524
tri 758 514 766 522 se
rect 766 514 932 522
tri 932 514 940 522 nw
tri 948 514 956 522 se
rect 956 514 1144 522
tri 1144 514 1152 522 nw
tri 1160 514 1168 522 se
rect 1168 519 1332 522
tri 1332 519 1335 522 nw
tri 1393 519 1396 522 se
rect 1396 519 1404 522
rect 1168 514 1327 519
tri 1327 514 1332 519 nw
tri 1388 514 1393 519 se
rect 1393 514 1404 519
rect 1412 514 1424 522
rect 1432 514 1444 522
rect 1452 514 1464 522
rect 1472 519 1489 522
tri 1489 519 1492 522 nw
tri 1509 519 1512 522 se
rect 1512 519 1514 522
rect 1472 514 1484 519
tri 1484 514 1489 519 nw
tri 1504 514 1509 519 se
rect 1509 514 1514 519
rect 1522 514 1534 522
rect 1542 514 1554 522
rect 1562 514 1574 522
rect 1582 514 1594 522
rect 1602 514 1614 522
tri 1614 514 1622 522 nw
tri 1684 514 1692 522 se
rect 1692 514 1720 522
rect 1728 514 1750 522
rect 1758 514 1782 522
tri 1782 514 1790 522 nw
tri 1798 514 1806 522 se
rect 1806 514 1810 522
rect 1818 514 1830 522
rect 1838 514 1860 522
rect 1868 514 1890 522
rect 1898 514 1920 522
rect 1928 514 1950 522
rect 1958 514 1980 522
rect 1988 514 2000 522
tri 756 512 758 514 se
rect 758 513 931 514
tri 931 513 932 514 nw
tri 947 513 948 514 se
rect 948 513 1142 514
rect 758 512 930 513
tri 930 512 931 513 nw
tri 946 512 947 513 se
rect 947 512 1142 513
tri 1142 512 1144 514 nw
tri 1158 512 1160 514 se
rect 1160 512 1325 514
tri 1325 512 1327 514 nw
tri 1386 512 1388 514 se
rect 1388 512 1482 514
tri 1482 512 1484 514 nw
tri 1502 512 1504 514 se
rect 1504 512 1612 514
tri 1612 512 1614 514 nw
tri 1682 512 1684 514 se
rect 1684 512 1780 514
tri 1780 512 1782 514 nw
tri 1796 512 1798 514 se
rect 1798 512 2000 514
tri 748 504 756 512 se
rect 756 504 923 512
tri 923 505 930 512 nw
tri 939 505 946 512 se
rect 946 505 1134 512
tri 923 504 924 505 sw
tri 938 504 939 505 se
rect 939 504 1134 505
tri 1134 504 1142 512 nw
tri 1150 504 1158 512 se
rect 1158 504 1317 512
tri 1317 504 1325 512 nw
tri 1378 504 1386 512 se
rect 1386 504 1394 512
rect 1402 504 1414 512
rect 1422 504 1434 512
rect 1442 504 1454 512
rect 1462 504 1474 512
tri 1474 504 1482 512 nw
tri 1494 504 1502 512 se
rect 1502 504 1504 512
rect 1512 504 1524 512
rect 1532 504 1544 512
rect 1552 504 1564 512
rect 1572 504 1584 512
rect 1592 504 1604 512
tri 1604 504 1612 512 nw
tri 1674 504 1682 512 se
rect 1682 504 1710 512
rect 1718 504 1740 512
rect 1748 504 1772 512
tri 1772 504 1780 512 nw
tri 1788 504 1796 512 se
rect 1796 504 1800 512
rect 1808 504 1840 512
rect 1848 504 1870 512
rect 1878 504 1900 512
rect 1908 504 1930 512
rect 1938 504 1960 512
rect 1968 504 1990 512
rect 1998 504 2000 512
tri 746 502 748 504 se
rect 748 502 924 504
tri 924 502 926 504 sw
tri 936 502 938 504 se
rect 938 502 1132 504
tri 1132 502 1134 504 nw
tri 1148 502 1150 504 se
rect 1150 502 1315 504
tri 1315 502 1317 504 nw
tri 1376 502 1378 504 se
rect 1378 502 1472 504
tri 1472 502 1474 504 nw
tri 1492 502 1494 504 se
rect 1494 502 1602 504
tri 1602 502 1604 504 nw
tri 1672 502 1674 504 se
rect 1674 502 1770 504
tri 1770 502 1772 504 nw
tri 1786 502 1788 504 se
rect 1788 502 2000 504
tri 738 494 746 502 se
rect 746 497 926 502
tri 926 497 931 502 sw
tri 931 497 936 502 se
rect 936 497 1127 502
tri 1127 497 1132 502 nw
tri 1143 497 1148 502 se
rect 1148 497 1307 502
rect 746 494 1124 497
tri 1124 494 1127 497 nw
tri 1140 494 1143 497 se
rect 1143 494 1307 497
tri 1307 494 1315 502 nw
tri 1368 494 1376 502 se
rect 1376 494 1384 502
rect 1392 494 1404 502
rect 1412 494 1424 502
rect 1432 494 1444 502
rect 1452 494 1464 502
tri 1464 494 1472 502 nw
tri 1484 494 1492 502 se
rect 1492 494 1494 502
rect 1502 494 1514 502
rect 1522 494 1534 502
rect 1542 494 1554 502
rect 1562 494 1574 502
rect 1582 494 1594 502
tri 1594 494 1602 502 nw
tri 1664 494 1672 502 se
rect 1672 494 1760 502
tri 736 492 738 494 se
rect 738 492 1122 494
tri 1122 492 1124 494 nw
tri 1138 492 1140 494 se
rect 1140 492 1305 494
tri 1305 492 1307 494 nw
tri 1366 492 1368 494 se
rect 1368 492 1462 494
tri 1462 492 1464 494 nw
tri 1482 492 1484 494 se
rect 1484 492 1592 494
tri 1592 492 1594 494 nw
tri 1662 492 1664 494 se
rect 1664 492 1760 494
tri 1760 492 1770 502 nw
tri 1776 492 1786 502 se
rect 1786 492 2000 502
tri 730 486 736 492 se
rect 736 486 1116 492
tri 1116 486 1122 492 nw
tri 1132 486 1138 492 se
rect 1138 486 1299 492
tri 1299 486 1305 492 nw
tri 1360 486 1366 492 se
rect 1366 486 1374 492
tri 728 484 730 486 se
rect 730 484 1114 486
tri 1114 484 1116 486 nw
tri 1130 484 1132 486 se
rect 1132 484 1297 486
tri 1297 484 1299 486 nw
tri 1358 484 1360 486 se
rect 1360 484 1374 486
rect 1382 484 1394 492
rect 1402 484 1414 492
rect 1422 484 1434 492
rect 1442 486 1456 492
tri 1456 486 1462 492 nw
tri 1476 486 1482 492 se
rect 1482 486 1484 492
rect 1442 484 1454 486
tri 1454 484 1456 486 nw
tri 1474 484 1476 486 se
rect 1476 484 1484 486
rect 1492 484 1504 492
rect 1512 484 1524 492
rect 1532 484 1544 492
rect 1552 484 1564 492
rect 1572 484 1584 492
tri 1584 484 1592 492 nw
tri 1654 484 1662 492 se
rect 1662 484 1680 492
rect 1688 484 1700 492
rect 1708 484 1720 492
rect 1728 484 1740 492
rect 1748 486 1754 492
tri 1754 486 1760 492 nw
tri 1770 486 1776 492 se
rect 1776 486 1790 492
rect 1748 484 1752 486
tri 1752 484 1754 486 nw
tri 1768 484 1770 486 se
rect 1770 484 1790 486
rect 1798 484 1810 492
rect 1818 484 1830 492
rect 1838 484 1850 492
rect 1858 484 1870 492
rect 1878 484 1880 492
tri 1880 484 1888 492 nw
tri 726 482 728 484 se
rect 728 482 1112 484
tri 1112 482 1114 484 nw
tri 1128 482 1130 484 se
rect 1130 482 1295 484
tri 1295 482 1297 484 nw
tri 1356 482 1358 484 se
rect 1358 482 1452 484
tri 1452 482 1454 484 nw
tri 1472 482 1474 484 se
rect 1474 482 1582 484
tri 1582 482 1584 484 nw
tri 1652 482 1654 484 se
rect 1654 482 1750 484
tri 1750 482 1752 484 nw
tri 1766 482 1768 484 se
rect 1768 482 1878 484
tri 1878 482 1880 484 nw
tri 718 474 726 482 se
rect 726 474 1104 482
tri 1104 474 1112 482 nw
tri 1120 474 1128 482 se
rect 1128 474 1287 482
tri 1287 474 1295 482 nw
tri 1348 474 1356 482 se
rect 1356 474 1364 482
rect 1372 474 1384 482
rect 1392 474 1404 482
rect 1412 474 1424 482
rect 1432 474 1444 482
tri 1444 474 1452 482 nw
tri 1464 474 1472 482 se
rect 1472 474 1474 482
rect 1482 474 1494 482
rect 1502 474 1514 482
rect 1522 474 1534 482
rect 1542 474 1554 482
rect 1562 474 1574 482
tri 1574 474 1582 482 nw
tri 1644 474 1652 482 se
rect 1652 474 1670 482
rect 1678 474 1690 482
rect 1698 474 1710 482
rect 1718 474 1730 482
rect 1738 474 1742 482
tri 1742 474 1750 482 nw
tri 1758 474 1766 482 se
rect 1766 474 1780 482
rect 1788 474 1800 482
rect 1808 474 1820 482
rect 1828 474 1840 482
rect 1848 474 1860 482
rect 1868 474 1870 482
tri 1870 474 1878 482 nw
tri 716 472 718 474 se
rect 718 472 1102 474
tri 1102 472 1104 474 nw
tri 1118 472 1120 474 se
rect 1120 472 1285 474
tri 1285 472 1287 474 nw
tri 1346 472 1348 474 se
rect 1348 472 1442 474
tri 1442 472 1444 474 nw
tri 1462 472 1464 474 se
rect 1464 472 1572 474
tri 1572 472 1574 474 nw
tri 1642 472 1644 474 se
rect 1644 472 1740 474
tri 1740 472 1742 474 nw
tri 1756 472 1758 474 se
rect 1758 472 1868 474
tri 1868 472 1870 474 nw
tri 708 464 716 472 se
rect 716 464 1094 472
tri 1094 464 1102 472 nw
tri 1110 464 1118 472 se
rect 1118 464 1277 472
tri 1277 464 1285 472 nw
tri 1338 464 1346 472 se
rect 1346 464 1354 472
rect 1362 464 1374 472
rect 1382 464 1394 472
rect 1402 464 1414 472
rect 1422 466 1436 472
tri 1436 466 1442 472 nw
tri 1456 466 1462 472 se
rect 1462 466 1464 472
rect 1422 464 1434 466
tri 1434 464 1436 466 nw
tri 1454 464 1456 466 se
rect 1456 464 1464 466
rect 1472 464 1484 472
rect 1492 464 1504 472
rect 1512 464 1524 472
rect 1532 464 1544 472
rect 1552 464 1564 472
tri 1564 464 1572 472 nw
tri 1634 464 1642 472 se
rect 1642 464 1660 472
rect 1668 464 1680 472
rect 1688 464 1700 472
rect 1708 464 1720 472
rect 1728 464 1732 472
tri 1732 464 1740 472 nw
tri 1748 464 1756 472 se
rect 1756 464 1770 472
rect 1778 464 1790 472
rect 1798 464 1810 472
rect 1818 464 1830 472
rect 1838 464 1850 472
rect 1858 464 1860 472
tri 1860 464 1868 472 nw
tri 706 462 708 464 se
rect 708 462 1092 464
tri 1092 462 1094 464 nw
tri 1108 462 1110 464 se
rect 1110 462 1275 464
tri 1275 462 1277 464 nw
tri 1336 462 1338 464 se
rect 1338 462 1432 464
tri 1432 462 1434 464 nw
tri 1452 462 1454 464 se
rect 1454 462 1562 464
tri 1562 462 1564 464 nw
tri 1632 462 1634 464 se
rect 1634 462 1730 464
tri 1730 462 1732 464 nw
tri 1746 462 1748 464 se
rect 1748 462 1858 464
tri 1858 462 1860 464 nw
tri 698 454 706 462 se
rect 706 454 1084 462
tri 1084 454 1092 462 nw
tri 1100 454 1108 462 se
rect 1108 454 1267 462
tri 1267 454 1275 462 nw
tri 1328 454 1336 462 se
rect 1336 454 1344 462
rect 1352 454 1364 462
rect 1372 454 1384 462
rect 1392 454 1404 462
rect 1412 454 1424 462
tri 1424 454 1432 462 nw
tri 1444 454 1452 462 se
rect 1452 454 1454 462
rect 1462 454 1474 462
rect 1482 454 1494 462
rect 1502 454 1514 462
rect 1522 454 1534 462
rect 1542 454 1554 462
tri 1554 454 1562 462 nw
tri 1624 454 1632 462 se
rect 1632 454 1650 462
rect 1658 454 1670 462
rect 1678 454 1690 462
rect 1698 454 1710 462
rect 1718 454 1722 462
tri 1722 454 1730 462 nw
tri 1738 454 1746 462 se
rect 1746 454 1760 462
rect 1768 454 1780 462
rect 1788 454 1800 462
rect 1808 454 1820 462
rect 1828 454 1840 462
rect 1848 460 1856 462
tri 1856 460 1858 462 nw
rect 1848 454 1850 460
tri 1850 454 1856 460 nw
tri 1914 454 1920 460 se
rect 1920 454 2000 460
tri 696 452 698 454 se
rect 698 452 1082 454
tri 1082 452 1084 454 nw
tri 1098 452 1100 454 se
rect 1100 452 1265 454
tri 1265 452 1267 454 nw
tri 1326 452 1328 454 se
rect 1328 452 1422 454
tri 1422 452 1424 454 nw
tri 1442 452 1444 454 se
rect 1444 452 1552 454
tri 1552 452 1554 454 nw
tri 1622 452 1624 454 se
rect 1624 452 1720 454
tri 1720 452 1722 454 nw
tri 1736 452 1738 454 se
rect 1738 452 1848 454
tri 1848 452 1850 454 nw
tri 1912 452 1914 454 se
rect 1914 452 2000 454
tri 688 444 696 452 se
rect 696 444 1074 452
tri 1074 444 1082 452 nw
tri 1090 444 1098 452 se
rect 1098 451 1264 452
tri 1264 451 1265 452 nw
tri 1325 451 1326 452 se
rect 1326 451 1334 452
rect 1098 444 1257 451
tri 1257 444 1264 451 nw
tri 1318 444 1325 451 se
rect 1325 444 1334 451
rect 1342 444 1354 452
rect 1362 444 1374 452
rect 1382 444 1394 452
rect 1402 444 1414 452
tri 1414 444 1422 452 nw
tri 1434 444 1442 452 se
rect 1442 444 1444 452
rect 1452 444 1464 452
rect 1472 444 1484 452
rect 1492 444 1504 452
rect 1512 444 1524 452
rect 1532 444 1544 452
tri 1544 444 1552 452 nw
tri 1614 444 1622 452 se
rect 1622 444 1640 452
rect 1648 444 1660 452
rect 1668 444 1680 452
rect 1688 444 1700 452
rect 1708 444 1712 452
tri 1712 444 1720 452 nw
tri 1728 444 1736 452 se
rect 1736 444 1750 452
rect 1758 444 1770 452
rect 1778 444 1790 452
rect 1798 444 1810 452
rect 1818 444 1830 452
rect 1838 444 1840 452
tri 1840 444 1848 452 nw
tri 1904 444 1912 452 se
rect 1912 444 2000 452
tri 686 442 688 444 se
rect 688 442 1072 444
tri 1072 442 1074 444 nw
tri 1088 442 1090 444 se
rect 1090 442 1255 444
tri 1255 442 1257 444 nw
tri 1316 442 1318 444 se
rect 1318 442 1412 444
tri 1412 442 1414 444 nw
tri 1432 442 1434 444 se
rect 1434 442 1542 444
tri 1542 442 1544 444 nw
tri 1612 442 1614 444 se
rect 1614 442 1710 444
tri 1710 442 1712 444 nw
tri 1726 442 1728 444 se
rect 1728 442 1838 444
tri 1838 442 1840 444 nw
tri 1902 442 1904 444 se
rect 1904 442 2000 444
tri 678 434 686 442 se
rect 686 434 1064 442
tri 1064 434 1072 442 nw
tri 1080 434 1088 442 se
rect 1088 434 1247 442
tri 1247 434 1255 442 nw
tri 1308 434 1316 442 se
rect 1316 434 1324 442
rect 1332 434 1344 442
rect 1352 434 1364 442
rect 1372 434 1384 442
rect 1392 434 1404 442
tri 1404 434 1412 442 nw
tri 1424 434 1432 442 se
rect 1432 434 1434 442
rect 1442 434 1454 442
rect 1462 434 1474 442
rect 1482 434 1494 442
rect 1502 434 1514 442
rect 1522 434 1534 442
tri 1534 434 1542 442 nw
tri 1604 434 1612 442 se
rect 1612 434 1630 442
rect 1638 434 1650 442
rect 1658 434 1670 442
rect 1678 434 1690 442
rect 1698 434 1702 442
tri 1702 434 1710 442 nw
tri 1718 434 1726 442 se
rect 1726 434 1740 442
rect 1748 434 1760 442
rect 1768 434 1780 442
rect 1788 434 1800 442
rect 1808 434 1820 442
rect 1828 434 1830 442
tri 1830 434 1838 442 nw
tri 1894 434 1902 442 se
rect 1902 434 2000 442
tri 676 432 678 434 se
rect 678 432 1062 434
tri 1062 432 1064 434 nw
tri 1078 432 1080 434 se
rect 1080 432 1245 434
tri 1245 432 1247 434 nw
tri 1306 432 1308 434 se
rect 1308 432 1402 434
tri 1402 432 1404 434 nw
tri 1422 432 1424 434 se
rect 1424 432 1532 434
tri 1532 432 1534 434 nw
tri 1602 432 1604 434 se
rect 1604 432 1700 434
tri 1700 432 1702 434 nw
tri 1716 432 1718 434 se
rect 1718 432 1828 434
tri 1828 432 1830 434 nw
tri 1892 432 1894 434 se
rect 1894 432 2000 434
tri 668 424 676 432 se
rect 676 424 1054 432
tri 1054 424 1062 432 nw
tri 1070 424 1078 432 se
rect 1078 424 1237 432
tri 1237 424 1245 432 nw
tri 1298 424 1306 432 se
rect 1306 424 1314 432
rect 1322 424 1334 432
rect 1342 424 1354 432
rect 1362 424 1374 432
rect 1382 424 1394 432
tri 1394 424 1402 432 nw
tri 1414 424 1422 432 se
rect 1422 424 1424 432
rect 1432 424 1444 432
rect 1452 424 1464 432
rect 1472 424 1484 432
rect 1492 424 1504 432
rect 1512 424 1524 432
tri 1524 424 1532 432 nw
tri 1594 424 1602 432 se
rect 1602 424 1620 432
rect 1628 424 1640 432
rect 1648 424 1660 432
rect 1668 424 1680 432
rect 1688 424 1692 432
tri 1692 424 1700 432 nw
tri 1708 424 1716 432 se
rect 1716 424 1730 432
rect 1738 424 1750 432
rect 1758 424 1770 432
rect 1778 424 1790 432
rect 1798 424 1810 432
rect 1818 424 1820 432
tri 1820 424 1828 432 nw
tri 1884 424 1892 432 se
rect 1892 424 2000 432
tri 666 422 668 424 se
rect 668 422 1052 424
tri 1052 422 1054 424 nw
tri 1068 422 1070 424 se
rect 1070 422 1235 424
tri 1235 422 1237 424 nw
tri 1296 422 1298 424 se
rect 1298 422 1392 424
tri 1392 422 1394 424 nw
tri 1412 422 1414 424 se
rect 1414 422 1522 424
tri 1522 422 1524 424 nw
tri 1592 422 1594 424 se
rect 1594 422 1690 424
tri 1690 422 1692 424 nw
tri 1706 422 1708 424 se
rect 1708 422 1818 424
tri 1818 422 1820 424 nw
tri 1882 422 1884 424 se
rect 1884 422 2000 424
tri 660 416 666 422 se
rect 666 416 1046 422
tri 1046 416 1052 422 nw
tri 1062 416 1068 422 se
rect 1068 416 1227 422
rect 660 414 1044 416
tri 1044 414 1046 416 nw
tri 1060 414 1062 416 se
rect 1062 414 1227 416
tri 1227 414 1235 422 nw
tri 1288 414 1296 422 se
rect 1296 414 1304 422
rect 1312 414 1324 422
rect 1332 414 1344 422
rect 1352 414 1364 422
rect 1372 414 1384 422
tri 1384 414 1392 422 nw
tri 1404 414 1412 422 se
rect 1412 414 1414 422
rect 1422 414 1434 422
rect 1442 414 1454 422
rect 1462 414 1474 422
rect 1482 414 1494 422
rect 1502 414 1514 422
tri 1514 414 1522 422 nw
tri 1584 414 1592 422 se
rect 1592 414 1610 422
rect 1618 414 1630 422
rect 1638 414 1650 422
rect 1658 414 1670 422
rect 1678 414 1682 422
tri 1682 414 1690 422 nw
tri 1698 414 1706 422 se
rect 1706 414 1720 422
rect 1728 414 1740 422
rect 1748 414 1760 422
rect 1768 414 1780 422
rect 1788 414 1800 422
rect 1808 414 1810 422
tri 1810 414 1818 422 nw
tri 1874 414 1882 422 se
rect 1882 414 2000 422
rect 660 412 1042 414
tri 1042 412 1044 414 nw
tri 1058 412 1060 414 se
rect 1060 412 1225 414
tri 1225 412 1227 414 nw
tri 1286 412 1288 414 se
rect 1288 412 1382 414
tri 1382 412 1384 414 nw
tri 1402 412 1404 414 se
rect 1404 412 1512 414
tri 1512 412 1514 414 nw
tri 1582 412 1584 414 se
rect 1584 412 1680 414
tri 1680 412 1682 414 nw
tri 1696 412 1698 414 se
rect 1698 412 1808 414
tri 1808 412 1810 414 nw
tri 1872 412 1874 414 se
rect 1874 412 2000 414
rect 660 406 1036 412
tri 1036 406 1042 412 nw
tri 1052 406 1058 412 se
rect 1058 406 1217 412
rect 660 404 1034 406
tri 1034 404 1036 406 nw
tri 1050 404 1052 406 se
rect 1052 404 1217 406
tri 1217 404 1225 412 nw
tri 1278 404 1286 412 se
rect 1286 404 1294 412
rect 1302 404 1314 412
rect 1322 404 1334 412
rect 1342 404 1354 412
rect 1362 404 1374 412
tri 1374 404 1382 412 nw
tri 1394 404 1402 412 se
rect 1402 404 1404 412
rect 1412 404 1424 412
rect 1432 404 1444 412
rect 1452 404 1464 412
rect 1472 404 1484 412
rect 1492 404 1504 412
tri 1504 404 1512 412 nw
tri 1574 404 1582 412 se
rect 1582 404 1600 412
rect 1608 404 1620 412
rect 1628 404 1640 412
rect 1648 404 1660 412
rect 1668 404 1672 412
tri 1672 404 1680 412 nw
tri 1688 404 1696 412 se
rect 1696 404 1710 412
rect 1718 404 1730 412
rect 1738 404 1750 412
rect 1758 404 1770 412
rect 1778 404 1790 412
rect 1798 404 1800 412
tri 1800 404 1808 412 nw
tri 1864 404 1872 412 se
rect 1872 404 2000 412
rect 660 402 1032 404
tri 1032 402 1034 404 nw
tri 1048 402 1050 404 se
rect 1050 402 1215 404
tri 1215 402 1217 404 nw
tri 1276 402 1278 404 se
rect 1278 402 1372 404
tri 1372 402 1374 404 nw
tri 1392 402 1394 404 se
rect 1394 402 1502 404
tri 1502 402 1504 404 nw
tri 1572 402 1574 404 se
rect 1574 402 1670 404
tri 1670 402 1672 404 nw
tri 1686 402 1688 404 se
rect 1688 402 1798 404
tri 1798 402 1800 404 nw
tri 1862 402 1864 404 se
rect 1864 402 2000 404
rect 660 394 1028 402
tri 1028 398 1032 402 nw
tri 1028 394 1032 398 sw
tri 1040 394 1048 402 se
rect 1048 394 1207 402
tri 1207 394 1215 402 nw
tri 1268 394 1276 402 se
rect 1276 394 1284 402
rect 1292 394 1304 402
rect 1312 394 1324 402
rect 1332 394 1344 402
rect 1352 394 1364 402
tri 1364 394 1372 402 nw
tri 1384 394 1392 402 se
rect 1392 394 1394 402
rect 1402 394 1414 402
rect 1422 394 1434 402
rect 1442 394 1454 402
rect 1462 394 1474 402
rect 1482 394 1494 402
tri 1494 394 1502 402 nw
tri 1564 394 1572 402 se
rect 1572 394 1590 402
rect 1598 394 1610 402
rect 1618 394 1630 402
rect 1638 394 1650 402
rect 1658 394 1662 402
tri 1662 394 1670 402 nw
tri 1678 394 1686 402 se
rect 1686 394 1700 402
rect 1708 394 1720 402
rect 1728 394 1740 402
rect 1748 394 1760 402
rect 1768 394 1780 402
rect 1788 394 1790 402
tri 1790 394 1798 402 nw
tri 1854 394 1862 402 se
rect 1862 394 2000 402
rect 660 392 1032 394
tri 1032 392 1034 394 sw
tri 1038 392 1040 394 se
rect 1040 392 1205 394
tri 1205 392 1207 394 nw
tri 1266 392 1268 394 se
rect 1268 392 1362 394
tri 1362 392 1364 394 nw
tri 1382 392 1384 394 se
rect 1384 392 1492 394
tri 1492 392 1494 394 nw
tri 1562 392 1564 394 se
rect 1564 392 1660 394
tri 1660 392 1662 394 nw
tri 1676 392 1678 394 se
rect 1678 392 1788 394
tri 1788 392 1790 394 nw
tri 1852 392 1854 394 se
rect 1854 392 2000 394
rect 660 390 1034 392
tri 1034 390 1036 392 sw
tri 1036 390 1038 392 se
rect 1038 390 1203 392
tri 1203 390 1205 392 nw
tri 1264 390 1266 392 se
rect 1266 390 1274 392
rect 660 384 1197 390
tri 1197 384 1203 390 nw
tri 1258 384 1264 390 se
rect 1264 384 1274 390
rect 1282 384 1294 392
rect 1302 384 1314 392
rect 1322 384 1334 392
rect 1342 390 1360 392
tri 1360 390 1362 392 nw
tri 1380 390 1382 392 se
rect 1382 390 1384 392
rect 1342 384 1354 390
tri 1354 384 1360 390 nw
tri 1374 384 1380 390 se
rect 1380 384 1384 390
rect 1392 384 1404 392
rect 1412 384 1424 392
rect 1432 384 1444 392
rect 1452 384 1464 392
rect 1472 384 1484 392
tri 1484 384 1492 392 nw
tri 1554 384 1562 392 se
rect 1562 384 1580 392
rect 1588 384 1600 392
rect 1608 384 1620 392
rect 1628 384 1640 392
rect 1648 388 1656 392
tri 1656 388 1660 392 nw
tri 1672 388 1676 392 se
rect 1676 388 1690 392
rect 1648 384 1652 388
tri 1652 384 1656 388 nw
tri 1668 384 1672 388 se
rect 1672 384 1690 388
rect 1698 384 1710 392
rect 1718 384 1730 392
rect 1738 384 1750 392
rect 1758 384 1770 392
rect 1778 384 1780 392
tri 1780 384 1788 392 nw
tri 1844 384 1852 392 se
rect 1852 384 2000 392
rect 660 382 1195 384
tri 1195 382 1197 384 nw
tri 1256 382 1258 384 se
rect 1258 382 1352 384
tri 1352 382 1354 384 nw
tri 1372 382 1374 384 se
rect 1374 382 1482 384
tri 1482 382 1484 384 nw
tri 1552 382 1554 384 se
rect 1554 382 1650 384
tri 1650 382 1652 384 nw
tri 1666 382 1668 384 se
rect 1668 382 1778 384
tri 1778 382 1780 384 nw
tri 1842 382 1844 384 se
rect 1844 382 2000 384
rect 660 374 1187 382
tri 1187 374 1195 382 nw
tri 1248 374 1256 382 se
rect 1256 374 1264 382
rect 1272 374 1284 382
rect 1292 374 1304 382
rect 1312 374 1324 382
rect 1332 378 1348 382
tri 1348 378 1352 382 nw
tri 1368 378 1372 382 se
rect 1372 378 1374 382
rect 1332 374 1344 378
tri 1344 374 1348 378 nw
tri 1364 374 1368 378 se
rect 1368 374 1374 378
rect 1382 374 1394 382
rect 1402 374 1414 382
rect 1422 374 1434 382
rect 1442 374 1454 382
rect 1462 374 1474 382
tri 1474 374 1482 382 nw
tri 1544 374 1552 382 se
rect 1552 374 1570 382
rect 1578 374 1590 382
rect 1598 374 1610 382
rect 1618 374 1630 382
rect 1638 374 1642 382
tri 1642 374 1650 382 nw
tri 1658 374 1666 382 se
rect 1666 374 1680 382
rect 1688 374 1700 382
rect 1708 374 1720 382
rect 1728 374 1740 382
rect 1748 374 1760 382
rect 1768 374 1770 382
tri 1770 374 1778 382 nw
tri 1834 374 1842 382 se
rect 1842 374 2000 382
rect 660 372 1185 374
tri 1185 372 1187 374 nw
tri 1246 372 1248 374 se
rect 1248 372 1342 374
tri 1342 372 1344 374 nw
tri 1362 372 1364 374 se
rect 1364 372 1472 374
tri 1472 372 1474 374 nw
tri 1542 372 1544 374 se
rect 1544 372 1640 374
tri 1640 372 1642 374 nw
tri 1656 372 1658 374 se
rect 1658 372 1768 374
tri 1768 372 1770 374 nw
tri 1832 372 1834 374 se
rect 1834 372 2000 374
rect 660 364 1177 372
tri 1177 364 1185 372 nw
tri 1238 364 1246 372 se
rect 1246 364 1254 372
rect 1262 364 1274 372
rect 1282 364 1294 372
rect 1302 364 1314 372
rect 1322 370 1340 372
tri 1340 370 1342 372 nw
tri 1360 370 1362 372 se
rect 1362 370 1364 372
rect 1322 364 1334 370
tri 1334 364 1340 370 nw
tri 1354 364 1360 370 se
rect 1360 364 1364 370
rect 1372 364 1384 372
rect 1392 364 1404 372
rect 1412 364 1424 372
rect 1432 364 1444 372
rect 1452 370 1470 372
tri 1470 370 1472 372 nw
tri 1540 370 1542 372 se
rect 1542 370 1560 372
rect 1452 364 1464 370
tri 1464 364 1470 370 nw
tri 1534 364 1540 370 se
rect 1540 364 1560 370
rect 1568 364 1580 372
rect 1588 364 1600 372
rect 1608 364 1620 372
rect 1628 364 1632 372
tri 1632 364 1640 372 nw
tri 1648 364 1656 372 se
rect 1656 364 1670 372
rect 1678 364 1690 372
rect 1698 364 1710 372
rect 1718 364 1730 372
rect 1738 364 1750 372
rect 1758 364 1760 372
tri 1760 364 1768 372 nw
tri 1824 364 1832 372 se
rect 1832 364 2000 372
rect 660 362 1175 364
tri 1175 362 1177 364 nw
tri 1236 362 1238 364 se
rect 1238 362 1332 364
tri 1332 362 1334 364 nw
tri 1352 362 1354 364 se
rect 1354 362 1462 364
tri 1462 362 1464 364 nw
tri 1532 362 1534 364 se
rect 1534 362 1630 364
tri 1630 362 1632 364 nw
tri 1646 362 1648 364 se
rect 1648 362 1758 364
tri 1758 362 1760 364 nw
tri 1822 362 1824 364 se
rect 1824 362 2000 364
rect 660 354 1167 362
tri 1167 354 1175 362 nw
tri 1228 354 1236 362 se
rect 1236 354 1244 362
rect 1252 354 1264 362
rect 1272 354 1284 362
rect 1292 354 1304 362
rect 1312 355 1325 362
tri 1325 355 1332 362 nw
tri 1348 358 1352 362 se
rect 1352 358 1354 362
tri 1345 355 1348 358 se
rect 1348 355 1354 358
rect 1312 354 1324 355
tri 1324 354 1325 355 nw
tri 1344 354 1345 355 se
rect 1345 354 1354 355
rect 1362 354 1374 362
rect 1382 354 1394 362
rect 1402 354 1414 362
rect 1422 354 1434 362
rect 1442 356 1456 362
tri 1456 356 1462 362 nw
tri 1526 356 1532 362 se
rect 1532 356 1550 362
rect 1442 354 1454 356
tri 1454 354 1456 356 nw
tri 1524 354 1526 356 se
rect 1526 354 1550 356
rect 1558 354 1570 362
rect 1578 354 1590 362
rect 1598 354 1610 362
rect 1618 354 1622 362
tri 1622 354 1630 362 nw
tri 1638 354 1646 362 se
rect 1646 354 1660 362
rect 1668 354 1680 362
rect 1688 354 1700 362
rect 1708 354 1720 362
rect 1728 354 1740 362
rect 1748 354 1750 362
tri 1750 354 1758 362 nw
tri 1814 354 1822 362 se
rect 1822 354 2000 362
rect 660 352 1165 354
tri 1165 352 1167 354 nw
tri 1226 352 1228 354 se
rect 1228 352 1322 354
tri 1322 352 1324 354 nw
tri 1342 352 1344 354 se
rect 1344 352 1452 354
tri 1452 352 1454 354 nw
tri 1522 352 1524 354 se
rect 1524 352 1620 354
tri 1620 352 1622 354 nw
tri 1636 352 1638 354 se
rect 1638 352 1748 354
tri 1748 352 1750 354 nw
tri 1812 352 1814 354 se
rect 1814 352 2000 354
rect 660 345 1158 352
tri 1158 345 1165 352 nw
tri 1219 345 1226 352 se
rect 1226 345 1234 352
rect 660 344 1157 345
tri 1157 344 1158 345 nw
tri 1218 344 1219 345 se
rect 1219 344 1234 345
rect 1242 344 1254 352
rect 1262 344 1274 352
rect 1282 344 1294 352
rect 1302 345 1315 352
tri 1315 345 1322 352 nw
tri 1335 345 1342 352 se
rect 1342 345 1344 352
rect 1302 344 1314 345
tri 1314 344 1315 345 nw
tri 1334 344 1335 345 se
rect 1335 344 1344 345
rect 1352 344 1364 352
rect 1372 344 1384 352
rect 1392 344 1404 352
rect 1412 344 1424 352
rect 1432 344 1444 352
tri 1444 344 1452 352 nw
tri 1514 344 1522 352 se
rect 1522 344 1540 352
rect 1548 344 1560 352
rect 1568 344 1580 352
rect 1588 344 1600 352
rect 1608 344 1612 352
tri 1612 344 1620 352 nw
tri 1628 344 1636 352 se
rect 1636 344 1650 352
rect 1658 344 1670 352
rect 1678 344 1690 352
rect 1698 344 1710 352
rect 1718 344 1730 352
rect 1738 344 1740 352
tri 1740 344 1748 352 nw
tri 1804 344 1812 352 se
rect 1812 344 2000 352
rect 660 342 1155 344
tri 1155 342 1157 344 nw
tri 1216 342 1218 344 se
rect 1218 342 1312 344
tri 1312 342 1314 344 nw
tri 1332 342 1334 344 se
rect 1334 342 1442 344
tri 1442 342 1444 344 nw
tri 1512 342 1514 344 se
rect 1514 342 1610 344
tri 1610 342 1612 344 nw
tri 1626 342 1628 344 se
rect 1628 342 1738 344
tri 1738 342 1740 344 nw
tri 1802 342 1804 344 se
rect 1804 342 2000 344
rect 660 334 1147 342
tri 1147 334 1155 342 nw
tri 1208 334 1216 342 se
rect 1216 334 1224 342
rect 1232 334 1244 342
rect 1252 334 1264 342
rect 1272 334 1284 342
rect 1292 334 1304 342
tri 1304 334 1312 342 nw
tri 1324 334 1332 342 se
rect 1332 334 1334 342
rect 1342 334 1354 342
rect 1362 334 1374 342
rect 1382 334 1394 342
rect 1402 334 1414 342
rect 1422 334 1434 342
tri 1434 334 1442 342 nw
tri 1504 334 1512 342 se
rect 1512 334 1530 342
rect 1538 334 1550 342
rect 1558 334 1570 342
rect 1578 334 1590 342
rect 1598 334 1602 342
tri 1602 334 1610 342 nw
tri 1618 334 1626 342 se
rect 1626 334 1640 342
rect 1648 334 1660 342
rect 1668 334 1680 342
rect 1688 334 1700 342
rect 1708 334 1720 342
rect 1728 334 1730 342
tri 1730 334 1738 342 nw
tri 1794 334 1802 342 se
rect 1802 334 2000 342
rect 660 332 1145 334
tri 1145 332 1147 334 nw
tri 1206 332 1208 334 se
rect 1208 332 1302 334
tri 1302 332 1304 334 nw
tri 1322 332 1324 334 se
rect 1324 332 1432 334
tri 1432 332 1434 334 nw
tri 1502 332 1504 334 se
rect 1504 332 1600 334
tri 1600 332 1602 334 nw
tri 1616 332 1618 334 se
rect 1618 332 1728 334
tri 1728 332 1730 334 nw
tri 1792 332 1794 334 se
rect 1794 332 2000 334
rect 660 324 1137 332
tri 1137 324 1145 332 nw
tri 1198 324 1206 332 se
rect 1206 324 1214 332
rect 1222 324 1234 332
rect 1242 324 1254 332
rect 1262 324 1274 332
rect 1282 324 1294 332
tri 1294 324 1302 332 nw
tri 1314 324 1322 332 se
rect 1322 324 1324 332
rect 1332 324 1344 332
rect 1352 324 1364 332
rect 1372 324 1384 332
rect 1392 324 1404 332
rect 1412 324 1424 332
tri 1424 324 1432 332 nw
tri 1494 324 1502 332 se
rect 1502 324 1520 332
rect 1528 324 1540 332
rect 1548 324 1560 332
rect 1568 324 1580 332
rect 1588 324 1592 332
tri 1592 324 1600 332 nw
tri 1608 324 1616 332 se
rect 1616 324 1630 332
rect 1638 324 1650 332
rect 1658 324 1670 332
rect 1678 324 1690 332
rect 1698 324 1710 332
rect 1718 324 1720 332
tri 1720 324 1728 332 nw
tri 1784 324 1792 332 se
rect 1792 324 2000 332
rect 660 322 1135 324
tri 1135 322 1137 324 nw
tri 1196 322 1198 324 se
rect 1198 322 1292 324
tri 1292 322 1294 324 nw
tri 1312 322 1314 324 se
rect 1314 322 1422 324
tri 1422 322 1424 324 nw
tri 1492 322 1494 324 se
rect 1494 322 1590 324
tri 1590 322 1592 324 nw
tri 1606 322 1608 324 se
rect 1608 322 1718 324
tri 1718 322 1720 324 nw
tri 1782 322 1784 324 se
rect 1784 322 2000 324
rect 660 314 1127 322
tri 1127 314 1135 322 nw
tri 1188 314 1196 322 se
rect 1196 314 1204 322
rect 1212 314 1224 322
rect 1232 314 1244 322
rect 1252 314 1264 322
rect 1272 314 1284 322
tri 1284 314 1292 322 nw
tri 1304 314 1312 322 se
rect 1312 314 1314 322
rect 1322 314 1334 322
rect 1342 314 1354 322
rect 1362 314 1374 322
rect 1382 314 1394 322
rect 1402 314 1414 322
tri 1414 314 1422 322 nw
tri 1484 314 1492 322 se
rect 1492 314 1510 322
rect 1518 314 1530 322
rect 1538 314 1550 322
rect 1558 314 1570 322
rect 1578 314 1582 322
tri 1582 314 1590 322 nw
tri 1598 314 1606 322 se
rect 1606 314 1620 322
rect 1628 314 1640 322
rect 1648 314 1660 322
rect 1668 314 1680 322
rect 1688 314 1700 322
rect 1708 314 1710 322
tri 1710 314 1718 322 nw
tri 1774 314 1782 322 se
rect 1782 314 2000 322
rect 660 312 1125 314
tri 1125 312 1127 314 nw
tri 1186 312 1188 314 se
rect 1188 312 1282 314
tri 1282 312 1284 314 nw
tri 1302 312 1304 314 se
rect 1304 312 1412 314
tri 1412 312 1414 314 nw
tri 1482 312 1484 314 se
rect 1484 312 1580 314
tri 1580 312 1582 314 nw
tri 1596 312 1598 314 se
rect 1598 312 1708 314
tri 1708 312 1710 314 nw
tri 1772 312 1774 314 se
rect 1774 312 2000 314
rect 660 260 1120 312
tri 1120 307 1125 312 nw
tri 1181 307 1186 312 se
rect 1186 307 1194 312
tri 1178 304 1181 307 se
rect 1181 304 1194 307
rect 1202 304 1214 312
rect 1222 304 1234 312
rect 1242 304 1254 312
rect 1262 304 1274 312
tri 1274 304 1282 312 nw
tri 1294 304 1302 312 se
rect 1302 304 1304 312
rect 1312 304 1324 312
rect 1332 304 1344 312
rect 1352 304 1364 312
rect 1372 304 1384 312
rect 1392 304 1404 312
tri 1404 304 1412 312 nw
tri 1476 306 1482 312 se
rect 1482 306 1500 312
rect 1456 304 1500 306
rect 1508 304 1520 312
rect 1528 304 1540 312
rect 1548 304 1560 312
rect 1568 304 1574 312
tri 1574 306 1580 312 nw
tri 1590 306 1596 312 se
rect 1596 306 1610 312
tri 1588 304 1590 306 se
rect 1590 304 1610 306
rect 1618 304 1630 312
rect 1638 304 1650 312
rect 1658 304 1670 312
rect 1678 304 1690 312
rect 1698 304 1700 312
tri 1700 304 1708 312 nw
tri 1764 304 1772 312 se
rect 1772 304 2000 312
tri 1176 302 1178 304 se
rect 1178 302 1272 304
tri 1272 302 1274 304 nw
tri 1292 302 1294 304 se
rect 1294 302 1402 304
tri 1402 302 1404 304 nw
rect 1456 302 1574 304
tri 1586 302 1588 304 se
rect 1588 302 1698 304
tri 1698 302 1700 304 nw
tri 1762 302 1764 304 se
rect 1764 302 2000 304
tri 1168 294 1176 302 se
rect 1176 294 1184 302
rect 1192 294 1204 302
rect 1212 294 1224 302
rect 1232 294 1244 302
rect 1252 296 1266 302
tri 1266 296 1272 302 nw
tri 1286 296 1292 302 se
rect 1292 296 1294 302
rect 1252 294 1264 296
tri 1264 294 1266 296 nw
tri 1284 294 1286 296 se
rect 1286 294 1294 296
rect 1302 294 1314 302
rect 1322 294 1334 302
rect 1342 294 1354 302
rect 1362 294 1374 302
rect 1382 294 1394 302
tri 1394 294 1402 302 nw
rect 1456 294 1490 302
rect 1498 294 1510 302
rect 1518 294 1530 302
rect 1538 294 1550 302
rect 1558 294 1574 302
tri 1578 294 1586 302 se
rect 1586 294 1600 302
rect 1608 294 1620 302
rect 1628 294 1640 302
rect 1648 294 1660 302
rect 1668 294 1680 302
rect 1688 294 1690 302
tri 1690 294 1698 302 nw
tri 1754 294 1762 302 se
rect 1762 294 2000 302
tri 1166 292 1168 294 se
rect 1168 292 1264 294
tri 1282 292 1284 294 se
rect 1284 292 1392 294
tri 1392 292 1394 294 nw
rect 1456 292 1574 294
tri 1576 292 1578 294 se
rect 1578 292 1688 294
tri 1688 292 1690 294 nw
tri 1752 292 1754 294 se
rect 1754 292 2000 294
tri 1158 284 1166 292 se
rect 1166 284 1174 292
rect 1182 284 1194 292
rect 1202 284 1214 292
rect 1222 284 1234 292
rect 1242 284 1264 292
tri 1274 284 1282 292 se
rect 1282 284 1284 292
rect 1292 284 1304 292
rect 1312 284 1324 292
rect 1332 284 1344 292
rect 1352 284 1364 292
rect 1372 284 1384 292
tri 1384 284 1392 292 nw
tri 1454 284 1456 286 se
rect 1456 284 1480 292
rect 1488 284 1500 292
rect 1508 284 1520 292
rect 1528 284 1540 292
rect 1548 290 1574 292
tri 1574 290 1576 292 se
rect 1576 290 1590 292
rect 1548 284 1590 290
rect 1598 284 1610 292
rect 1618 284 1630 292
rect 1638 284 1650 292
rect 1658 284 1670 292
rect 1678 290 1686 292
tri 1686 290 1688 292 nw
tri 1750 290 1752 292 se
rect 1752 290 2000 292
rect 1678 284 1680 290
tri 1680 284 1686 290 nw
tri 1744 284 1750 290 se
rect 1750 284 2000 290
tri 1156 282 1158 284 se
rect 1158 282 1264 284
tri 1272 282 1274 284 se
rect 1274 282 1382 284
tri 1382 282 1384 284 nw
tri 1452 282 1454 284 se
rect 1454 282 1678 284
tri 1678 282 1680 284 nw
tri 1742 282 1744 284 se
rect 1744 282 2000 284
rect 660 42 810 260
rect 820 42 960 260
rect 970 42 1120 260
rect 660 0 1120 42
tri 1152 278 1156 282 se
rect 1156 278 1164 282
rect 1152 274 1164 278
rect 1172 274 1184 282
rect 1192 274 1204 282
rect 1212 274 1224 282
rect 1232 276 1264 282
tri 1268 278 1272 282 se
rect 1272 278 1274 282
tri 1264 276 1266 278 sw
tri 1266 276 1268 278 se
rect 1268 276 1274 278
rect 1232 274 1274 276
rect 1282 274 1294 282
rect 1302 274 1314 282
rect 1322 274 1334 282
rect 1342 274 1354 282
rect 1362 274 1374 282
tri 1374 274 1382 282 nw
tri 1444 274 1452 282 se
rect 1452 274 1470 282
rect 1478 274 1490 282
rect 1498 274 1510 282
rect 1518 274 1530 282
rect 1538 274 1580 282
rect 1588 274 1600 282
rect 1608 274 1620 282
rect 1628 274 1640 282
rect 1648 274 1660 282
rect 1668 276 1672 282
tri 1672 276 1678 282 nw
tri 1736 276 1742 282 se
rect 1742 276 2000 282
rect 1668 274 1670 276
tri 1670 274 1672 276 nw
tri 1734 274 1736 276 se
rect 1736 274 2000 276
rect 1152 272 1372 274
tri 1372 272 1374 274 nw
tri 1442 272 1444 274 se
rect 1444 272 1668 274
tri 1668 272 1670 274 nw
tri 1732 272 1734 274 se
rect 1734 272 2000 274
rect 1152 244 1154 272
rect 1162 244 1174 272
rect 1182 264 1194 272
rect 1202 264 1214 272
rect 1222 264 1264 272
rect 1182 262 1264 264
rect 1182 244 1204 262
rect 1212 244 1234 262
rect 1242 244 1264 262
rect 1272 264 1284 272
rect 1292 264 1304 272
rect 1312 264 1324 272
rect 1272 262 1324 264
rect 1272 244 1294 262
rect 1302 244 1324 262
rect 1332 264 1344 272
rect 1352 264 1364 272
tri 1364 264 1372 272 nw
tri 1434 264 1442 272 se
rect 1442 264 1460 272
rect 1468 264 1480 272
rect 1488 264 1500 272
rect 1508 264 1520 272
rect 1528 264 1570 272
rect 1578 264 1590 272
rect 1598 264 1610 272
rect 1618 264 1630 272
rect 1638 264 1650 272
rect 1658 264 1660 272
tri 1660 264 1668 272 nw
tri 1724 264 1732 272 se
rect 1732 264 2000 272
rect 1332 262 1362 264
tri 1362 262 1364 264 nw
tri 1432 262 1434 264 se
rect 1434 262 1658 264
tri 1658 262 1660 264 nw
tri 1722 262 1724 264 se
rect 1724 262 2000 264
rect 1332 260 1360 262
tri 1360 260 1362 262 nw
tri 1430 260 1432 262 se
rect 1432 260 1450 262
rect 1332 254 1354 260
tri 1354 254 1360 260 nw
tri 1424 254 1430 260 se
rect 1430 254 1450 260
rect 1458 254 1470 262
rect 1478 254 1490 262
rect 1498 254 1510 262
rect 1518 254 1560 262
rect 1568 254 1580 262
rect 1588 254 1600 262
rect 1608 254 1620 262
rect 1628 254 1640 262
rect 1648 254 1650 262
tri 1650 254 1658 262 nw
tri 1714 254 1722 262 se
rect 1722 254 2000 262
rect 1332 252 1352 254
tri 1352 252 1354 254 nw
tri 1422 252 1424 254 se
rect 1424 252 1648 254
tri 1648 252 1650 254 nw
tri 1712 252 1714 254 se
rect 1714 252 2000 254
rect 1332 248 1348 252
tri 1348 248 1352 252 nw
tri 1418 248 1422 252 se
rect 1422 248 1440 252
rect 1332 244 1344 248
tri 1344 244 1348 248 nw
tri 1414 244 1418 248 se
rect 1418 244 1440 248
rect 1448 244 1460 252
rect 1468 244 1480 252
rect 1488 244 1500 252
rect 1508 244 1550 252
rect 1558 244 1570 252
rect 1578 244 1590 252
rect 1598 244 1610 252
rect 1618 244 1630 252
rect 1638 244 1640 252
tri 1640 244 1648 252 nw
tri 1704 244 1712 252 se
rect 1712 246 1916 252
tri 1916 246 1922 252 nw
tri 1922 246 1928 252 ne
rect 1712 244 1908 246
rect 1152 242 1342 244
tri 1342 242 1344 244 nw
tri 1412 242 1414 244 se
rect 1414 242 1638 244
tri 1638 242 1640 244 nw
tri 1702 242 1704 244 se
rect 1704 242 1908 244
rect 1152 234 1164 242
rect 1172 234 1194 242
rect 1202 234 1224 242
rect 1232 234 1254 242
rect 1262 234 1284 242
rect 1292 234 1314 242
rect 1322 234 1334 242
tri 1334 234 1342 242 nw
tri 1404 234 1412 242 se
rect 1412 234 1430 242
rect 1438 234 1450 242
rect 1458 234 1470 242
rect 1478 234 1490 242
rect 1498 234 1540 242
rect 1548 234 1560 242
rect 1568 234 1580 242
rect 1588 234 1600 242
rect 1608 234 1620 242
rect 1628 234 1630 242
tri 1630 234 1638 242 nw
tri 1694 234 1702 242 se
rect 1702 238 1908 242
tri 1908 238 1916 246 nw
tri 1920 238 1928 246 se
rect 1928 238 2000 252
rect 1702 234 1896 238
rect 1152 232 1332 234
tri 1332 232 1334 234 nw
tri 1402 232 1404 234 se
rect 1404 232 1628 234
tri 1628 232 1630 234 nw
tri 1692 232 1694 234 se
rect 1694 232 1896 234
rect 1152 224 1174 232
rect 1182 224 1204 232
rect 1212 224 1234 232
rect 1242 224 1264 232
rect 1272 224 1294 232
rect 1302 224 1324 232
tri 1324 224 1332 232 nw
tri 1394 224 1402 232 se
rect 1402 224 1420 232
rect 1428 224 1440 232
rect 1448 224 1460 232
rect 1468 224 1480 232
rect 1488 224 1530 232
rect 1538 224 1550 232
rect 1558 224 1570 232
rect 1578 224 1590 232
rect 1598 224 1610 232
rect 1618 224 1620 232
tri 1620 224 1628 232 nw
tri 1684 224 1692 232 se
rect 1692 226 1896 232
tri 1896 226 1908 238 nw
tri 1908 226 1920 238 se
rect 1920 226 2000 238
rect 1692 224 1884 226
rect 1152 222 1322 224
tri 1322 222 1324 224 nw
tri 1392 222 1394 224 se
rect 1394 222 1618 224
tri 1618 222 1620 224 nw
tri 1682 222 1684 224 se
rect 1684 222 1884 224
rect 1152 214 1164 222
rect 1172 214 1194 222
rect 1202 214 1224 222
rect 1232 214 1254 222
rect 1262 214 1284 222
rect 1292 214 1314 222
tri 1314 214 1322 222 nw
tri 1384 214 1392 222 se
rect 1392 214 1410 222
rect 1418 214 1430 222
rect 1438 214 1450 222
rect 1458 214 1470 222
rect 1478 214 1520 222
rect 1528 214 1540 222
rect 1548 214 1560 222
rect 1568 214 1580 222
rect 1588 214 1600 222
rect 1608 214 1610 222
tri 1610 214 1618 222 nw
tri 1674 214 1682 222 se
rect 1682 214 1884 222
tri 1884 214 1896 226 nw
tri 1896 214 1908 226 se
rect 1908 214 2000 226
rect 1152 212 1312 214
tri 1312 212 1314 214 nw
tri 1382 212 1384 214 se
rect 1384 212 1608 214
tri 1608 212 1610 214 nw
tri 1672 212 1674 214 se
rect 1674 212 1872 214
rect 1152 204 1174 212
rect 1182 204 1204 212
rect 1212 204 1234 212
rect 1242 204 1264 212
rect 1272 204 1294 212
rect 1302 204 1312 212
tri 1374 204 1382 212 se
rect 1382 204 1400 212
rect 1408 204 1420 212
rect 1428 204 1440 212
rect 1448 204 1460 212
rect 1468 204 1510 212
rect 1518 204 1530 212
rect 1538 204 1550 212
rect 1558 204 1570 212
rect 1578 204 1590 212
rect 1598 204 1600 212
tri 1600 204 1608 212 nw
tri 1664 204 1672 212 se
rect 1672 204 1872 212
rect 1152 202 1312 204
tri 1372 202 1374 204 se
rect 1374 202 1598 204
tri 1598 202 1600 204 nw
tri 1662 202 1664 204 se
rect 1664 202 1872 204
tri 1872 202 1884 214 nw
tri 1884 202 1896 214 se
rect 1896 202 2000 214
rect 1152 194 1164 202
rect 1172 194 1194 202
rect 1202 194 1224 202
rect 1232 194 1254 202
rect 1262 194 1284 202
rect 1292 194 1312 202
tri 1364 194 1372 202 se
rect 1372 194 1390 202
rect 1398 194 1410 202
rect 1418 194 1430 202
rect 1438 194 1450 202
rect 1458 194 1500 202
rect 1508 194 1520 202
rect 1528 194 1540 202
rect 1548 194 1560 202
rect 1568 194 1580 202
rect 1588 194 1590 202
tri 1590 194 1598 202 nw
tri 1654 194 1662 202 se
rect 1662 194 1860 202
rect 1152 192 1312 194
tri 1362 192 1364 194 se
rect 1364 192 1588 194
tri 1588 192 1590 194 nw
tri 1652 192 1654 194 se
rect 1654 192 1860 194
rect 1152 184 1174 192
rect 1182 184 1204 192
rect 1212 184 1234 192
rect 1242 184 1264 192
rect 1272 184 1294 192
rect 1302 184 1312 192
tri 1354 184 1362 192 se
rect 1362 184 1380 192
rect 1388 184 1400 192
rect 1408 184 1420 192
rect 1428 184 1440 192
rect 1448 184 1490 192
rect 1498 184 1510 192
rect 1518 184 1530 192
rect 1538 184 1550 192
rect 1558 184 1570 192
rect 1578 184 1580 192
tri 1580 184 1588 192 nw
tri 1644 184 1652 192 se
rect 1652 190 1860 192
tri 1860 190 1872 202 nw
tri 1872 190 1884 202 se
rect 1884 190 2000 202
rect 1652 184 1848 190
rect 1152 182 1312 184
rect 1152 174 1164 182
rect 1172 174 1194 182
rect 1202 174 1224 182
rect 1232 174 1254 182
rect 1262 174 1284 182
rect 1292 174 1312 182
rect 1152 172 1312 174
rect 1152 164 1174 172
rect 1182 164 1204 172
rect 1212 164 1234 172
rect 1242 164 1264 172
rect 1272 164 1294 172
rect 1302 164 1312 172
rect 1152 162 1312 164
rect 1152 154 1164 162
rect 1172 154 1194 162
rect 1202 154 1224 162
rect 1232 154 1254 162
rect 1262 154 1284 162
rect 1292 154 1312 162
rect 1152 152 1312 154
rect 1152 144 1174 152
rect 1182 144 1204 152
rect 1212 144 1234 152
rect 1242 144 1264 152
rect 1272 144 1294 152
rect 1302 144 1312 152
rect 1152 142 1312 144
rect 1152 134 1164 142
rect 1172 134 1194 142
rect 1202 134 1224 142
rect 1232 134 1254 142
rect 1262 134 1284 142
rect 1292 134 1312 142
rect 1152 132 1312 134
rect 1152 124 1174 132
rect 1182 124 1204 132
rect 1212 124 1234 132
rect 1242 124 1264 132
rect 1272 124 1294 132
rect 1302 124 1312 132
rect 1152 122 1312 124
rect 1152 114 1164 122
rect 1172 114 1194 122
rect 1202 114 1224 122
rect 1232 114 1254 122
rect 1262 114 1284 122
rect 1292 114 1312 122
rect 1152 112 1312 114
rect 1152 104 1174 112
rect 1182 104 1204 112
rect 1212 104 1234 112
rect 1242 104 1264 112
rect 1272 104 1294 112
rect 1302 104 1312 112
rect 1152 102 1312 104
rect 1152 94 1164 102
rect 1172 94 1194 102
rect 1202 94 1224 102
rect 1232 94 1254 102
rect 1262 94 1284 102
rect 1292 94 1312 102
rect 1152 92 1312 94
rect 1152 84 1174 92
rect 1182 84 1204 92
rect 1212 84 1234 92
rect 1242 84 1264 92
rect 1272 84 1294 92
rect 1302 84 1312 92
rect 1152 82 1312 84
rect 1152 74 1164 82
rect 1172 74 1194 82
rect 1202 74 1224 82
rect 1232 74 1254 82
rect 1262 74 1284 82
rect 1292 74 1312 82
rect 1152 72 1312 74
rect 1152 64 1174 72
rect 1182 64 1204 72
rect 1212 64 1234 72
rect 1242 64 1264 72
rect 1272 64 1294 72
rect 1302 64 1312 72
rect 1152 62 1312 64
rect 1152 54 1164 62
rect 1172 54 1194 62
rect 1202 54 1224 62
rect 1232 54 1254 62
rect 1262 54 1284 62
rect 1292 54 1312 62
rect 1152 52 1312 54
rect 1152 44 1174 52
rect 1182 44 1204 52
rect 1212 44 1234 52
rect 1242 44 1264 52
rect 1272 44 1294 52
rect 1302 44 1312 52
rect 1152 42 1312 44
rect 1152 34 1164 42
rect 1172 34 1194 42
rect 1202 34 1224 42
rect 1232 34 1254 42
rect 1262 34 1284 42
rect 1292 34 1312 42
rect 1152 32 1312 34
rect 1152 24 1174 32
rect 1182 24 1204 32
rect 1212 24 1234 32
rect 1242 24 1264 32
rect 1272 24 1294 32
rect 1302 24 1312 32
rect 1152 22 1312 24
rect 1152 14 1164 22
rect 1172 14 1194 22
rect 1202 14 1224 22
rect 1232 14 1254 22
rect 1262 14 1284 22
rect 1292 14 1312 22
rect 1152 12 1312 14
rect 1152 4 1174 12
rect 1182 4 1204 12
rect 1212 4 1234 12
rect 1242 4 1264 12
rect 1272 4 1294 12
rect 1302 4 1312 12
rect 1152 0 1312 4
tri 1348 178 1354 184 se
rect 1354 178 1574 184
tri 1574 178 1580 184 nw
tri 1638 178 1644 184 se
rect 1644 178 1848 184
tri 1848 178 1860 190 nw
tri 1860 178 1872 190 se
rect 1872 178 2000 190
rect 1348 172 1568 178
tri 1568 172 1574 178 nw
tri 1632 172 1638 178 se
rect 1638 172 1836 178
rect 1348 144 1360 172
rect 1368 144 1380 172
rect 1388 144 1400 172
rect 1348 142 1400 144
rect 1348 134 1370 142
rect 1378 134 1400 142
rect 1408 144 1420 172
rect 1428 144 1470 172
rect 1478 144 1490 172
rect 1408 142 1490 144
rect 1408 134 1430 142
rect 1438 134 1460 142
rect 1468 134 1490 142
rect 1498 144 1510 172
rect 1518 144 1530 172
rect 1538 164 1550 172
rect 1558 164 1560 172
tri 1560 164 1568 172 nw
tri 1624 164 1632 172 se
rect 1632 166 1836 172
tri 1836 166 1848 178 nw
tri 1848 166 1860 178 se
rect 1860 166 2000 178
rect 1632 164 1826 166
rect 1538 162 1558 164
tri 1558 162 1560 164 nw
tri 1622 162 1624 164 se
rect 1624 162 1826 164
rect 1538 154 1550 162
tri 1550 154 1558 162 nw
tri 1614 154 1622 162 se
rect 1622 156 1826 162
tri 1826 156 1836 166 nw
tri 1838 156 1848 166 se
rect 1848 156 2000 166
rect 1622 154 1814 156
rect 1538 152 1548 154
tri 1548 152 1550 154 nw
tri 1612 152 1614 154 se
rect 1614 152 1814 154
rect 1538 144 1540 152
tri 1540 144 1548 152 nw
tri 1604 144 1612 152 se
rect 1612 144 1814 152
tri 1814 144 1826 156 nw
tri 1826 144 1838 156 se
rect 1838 144 2000 156
rect 1498 142 1538 144
tri 1538 142 1540 144 nw
tri 1602 142 1604 144 se
rect 1604 142 1802 144
rect 1498 134 1530 142
tri 1530 134 1538 142 nw
tri 1594 134 1602 142 se
rect 1602 134 1802 142
rect 1348 132 1528 134
tri 1528 132 1530 134 nw
tri 1592 132 1594 134 se
rect 1594 132 1802 134
tri 1802 132 1814 144 nw
tri 1814 132 1826 144 se
rect 1826 132 2000 144
rect 1348 124 1360 132
rect 1368 124 1390 132
rect 1398 124 1420 132
rect 1428 124 1450 132
rect 1458 124 1480 132
rect 1488 124 1520 132
tri 1520 124 1528 132 nw
tri 1584 124 1592 132 se
rect 1592 124 1790 132
rect 1348 122 1518 124
tri 1518 122 1520 124 nw
tri 1582 122 1584 124 se
rect 1584 122 1790 124
rect 1348 114 1370 122
rect 1378 114 1400 122
rect 1408 114 1430 122
rect 1438 114 1460 122
rect 1468 114 1490 122
rect 1498 114 1510 122
tri 1510 114 1518 122 nw
tri 1574 114 1582 122 se
rect 1582 120 1790 122
tri 1790 120 1802 132 nw
tri 1802 120 1814 132 se
rect 1814 124 2000 132
rect 1814 120 1964 124
rect 1582 114 1778 120
rect 1348 112 1508 114
tri 1508 112 1510 114 nw
tri 1572 112 1574 114 se
rect 1574 112 1778 114
rect 1348 104 1360 112
rect 1368 104 1390 112
rect 1398 104 1420 112
rect 1428 104 1450 112
rect 1458 104 1480 112
rect 1488 104 1508 112
rect 1348 102 1508 104
rect 1348 94 1370 102
rect 1378 94 1400 102
rect 1408 94 1430 102
rect 1438 94 1460 102
rect 1468 94 1490 102
rect 1498 94 1508 102
rect 1348 92 1508 94
rect 1348 84 1360 92
rect 1368 84 1390 92
rect 1398 84 1420 92
rect 1428 84 1450 92
rect 1458 84 1480 92
rect 1488 84 1508 92
rect 1348 82 1508 84
rect 1348 74 1370 82
rect 1378 74 1400 82
rect 1408 74 1430 82
rect 1438 74 1460 82
rect 1468 74 1490 82
rect 1498 74 1508 82
rect 1348 72 1508 74
rect 1348 64 1360 72
rect 1368 64 1390 72
rect 1398 64 1420 72
rect 1428 64 1450 72
rect 1458 64 1480 72
rect 1488 64 1508 72
rect 1348 62 1508 64
rect 1348 54 1370 62
rect 1378 54 1400 62
rect 1408 54 1430 62
rect 1438 54 1460 62
rect 1468 54 1490 62
rect 1498 54 1508 62
rect 1348 52 1508 54
rect 1348 44 1360 52
rect 1368 44 1390 52
rect 1398 44 1420 52
rect 1428 44 1450 52
rect 1458 44 1480 52
rect 1488 44 1508 52
rect 1348 42 1508 44
rect 1348 34 1370 42
rect 1378 34 1400 42
rect 1408 34 1430 42
rect 1438 34 1460 42
rect 1468 34 1490 42
rect 1498 34 1508 42
rect 1348 32 1508 34
rect 1348 24 1360 32
rect 1368 24 1390 32
rect 1398 24 1420 32
rect 1428 24 1450 32
rect 1458 24 1480 32
rect 1488 24 1508 32
rect 1348 22 1508 24
rect 1348 14 1370 22
rect 1378 14 1400 22
rect 1408 14 1430 22
rect 1438 14 1460 22
rect 1468 14 1490 22
rect 1498 14 1508 22
rect 1348 12 1508 14
rect 1348 4 1360 12
rect 1368 4 1390 12
rect 1398 4 1420 12
rect 1428 4 1450 12
rect 1458 4 1480 12
rect 1488 4 1508 12
rect 1348 0 1508 4
tri 1540 80 1572 112 se
rect 1572 108 1778 112
tri 1778 108 1790 120 nw
tri 1790 108 1802 120 se
rect 1802 116 1964 120
tri 1964 116 1972 124 nw
tri 1972 116 1980 124 ne
rect 1802 108 1948 116
rect 1572 96 1766 108
tri 1766 96 1778 108 nw
tri 1778 96 1790 108 se
rect 1790 100 1948 108
tri 1948 100 1964 116 nw
tri 1964 100 1980 116 se
rect 1980 100 2000 124
rect 1790 96 1936 100
rect 1572 84 1754 96
tri 1754 84 1766 96 nw
tri 1766 84 1778 96 se
rect 1778 88 1936 96
tri 1936 88 1948 100 nw
tri 1952 88 1964 100 se
rect 1964 88 2000 100
rect 1778 84 1920 88
rect 1572 80 1750 84
tri 1750 80 1754 84 nw
tri 1762 80 1766 84 se
rect 1766 80 1920 84
rect 1540 72 1748 80
tri 1748 78 1750 80 nw
tri 1760 78 1762 80 se
rect 1762 78 1920 80
tri 1748 72 1754 78 sw
tri 1754 72 1760 78 se
rect 1760 72 1920 78
tri 1920 72 1936 88 nw
tri 1936 72 1952 88 se
rect 1952 72 2000 88
rect 1540 56 1904 72
tri 1904 56 1920 72 nw
tri 1920 56 1936 72 se
rect 1936 56 2000 72
rect 1540 40 1888 56
tri 1888 40 1904 56 nw
tri 1904 40 1920 56 se
rect 1920 40 2000 56
rect 1540 37 1885 40
tri 1885 37 1888 40 nw
tri 1901 37 1904 40 se
rect 1904 37 2000 40
rect 1540 21 1877 37
tri 1877 29 1885 37 nw
tri 1893 29 1901 37 se
rect 1901 29 2000 37
tri 1877 21 1885 29 sw
tri 1885 21 1893 29 se
rect 1893 21 2000 29
rect 1540 0 2000 21
<< labels >>
flabel nwell 2000 -6 2000 -6 6 FreeSans 16 0 0 0 VddNW
flabel nwell 1340 0 1340 0 8 FreeSans 16 270 0 0 VddNW
flabel nsubstratendiff 1346 0 1346 0 8 FreeSans 16 270 0 0 VddAct
flabel metal2 2000 0 2000 0 6 FreeSans 16 0 0 0 VddAct
flabel psubstratepdiff 660 0 660 0 8 FreeSans 16 270 0 0 GndAct
flabel psubstratepdiff 2000 686 2000 686 6 FreeSans 16 0 0 0 GndAct
flabel metal2 1540 0 1540 0 8 FreeSans 16 270 0 0 GndM2A
flabel metal2 2000 0 2000 0 6 FreeSans 16 0 0 0 GndM2A
flabel metal2 2000 688 2000 688 6 FreeSans 16 0 0 0 GndM2B
flabel metal2 1152 0 1152 0 8 FreeSans 16 270 0 0 GndM2B
flabel metal2 660 0 660 0 8 FreeSans 16 270 0 0 VddM2A
flabel metal2 2000 880 2000 880 6 FreeSans 16 0 0 0 VddM2A
flabel metal2 1348 0 1348 0 8 FreeSans 16 270 0 0 VddM2B
flabel metal2 2000 492 2000 492 6 FreeSans 16 0 0 0 VddM2B
<< properties >>
string path 1485.000 936.000 1822.500 1273.500 1822.500 94.500 1845.000 94.500 1845.000 585.000 1822.500 585.000 1822.500 1273.500 3366.000 2817.000 3366.000 2425.500 2076.750 1136.250 2094.750 1118.250 2160.000 1183.500 2160.000 94.500 2182.500 94.500 2182.500 585.000 2160.000 585.000 2160.000 1183.500 3384.000 2407.500 3366.000 2425.500 3366.000 2817.000 3564.000 3015.000 3579.750 3015.000 3579.750 2162.250 2313.000 895.500 2331.000 877.500 3597.750 2144.250 3579.750 2162.250 3579.750 3015.000 3915.000 3015.000 3915.000 2317.500 4405.500 2317.500 4405.500 2340.000 3915.000 2340.000 3915.000 2655.000 4405.500 2655.000 4405.500 2677.500 3915.000 2677.500 3915.000 3015.000 4500.000 3015.000 4500.000 1980.000 3809.250 1980.000 2520.000 690.750 2520.000 0.000 1485.000 0.000 1485.000 936.000 
<< end >>
