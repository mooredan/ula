magic
tech amic5n
timestamp 1625244852
<< nwell >>
rect -130 550 1030 1495
rect 105 150 795 550
<< polysilicon >>
rect 105 1240 795 1290
rect 105 1220 225 1240
rect 105 1170 125 1220
rect 175 1170 225 1220
rect 675 1220 795 1240
rect 105 1120 225 1170
rect 675 1170 725 1220
rect 775 1170 795 1220
rect 105 1070 125 1120
rect 175 1070 225 1120
rect 675 1120 795 1170
rect 675 1070 725 1120
rect 775 1070 795 1120
rect 105 1020 225 1070
rect 675 1020 795 1070
rect 105 970 125 1020
rect 175 970 225 1020
rect 105 920 225 970
rect 675 970 725 1020
rect 775 970 795 1020
rect 105 870 125 920
rect 175 870 225 920
rect 675 920 795 970
rect 105 820 225 870
rect 675 870 725 920
rect 775 870 795 920
rect 105 770 125 820
rect 175 770 225 820
rect 675 820 795 870
rect 105 720 225 770
rect 675 770 725 820
rect 775 770 795 820
rect 105 670 125 720
rect 175 670 225 720
rect 675 720 795 770
rect 105 620 225 670
rect 675 670 725 720
rect 775 670 795 720
rect 105 570 125 620
rect 175 570 225 620
rect 675 620 795 670
rect 105 520 225 570
rect 675 570 725 620
rect 775 570 795 620
rect 675 520 795 570
rect 105 470 125 520
rect 175 470 225 520
rect 675 470 725 520
rect 775 470 795 520
rect 105 420 225 470
rect 105 370 125 420
rect 175 370 225 420
rect 675 420 795 470
rect 105 320 225 370
rect 675 370 725 420
rect 775 370 795 420
rect 105 270 125 320
rect 175 270 225 320
rect 675 320 795 370
rect 105 220 225 270
rect 675 270 725 320
rect 775 270 795 320
rect 105 170 125 220
rect 175 200 225 220
rect 675 220 795 270
rect 675 200 725 220
rect 175 170 725 200
rect 775 170 795 220
rect 105 150 795 170
<< polycontact >>
rect 125 1170 175 1220
rect 725 1170 775 1220
rect 125 1070 175 1120
rect 725 1070 775 1120
rect 125 970 175 1020
rect 725 970 775 1020
rect 125 870 175 920
rect 725 870 775 920
rect 125 770 175 820
rect 725 770 775 820
rect 125 670 175 720
rect 725 670 775 720
rect 125 570 175 620
rect 725 570 775 620
rect 125 470 175 520
rect 725 470 775 520
rect 125 370 175 420
rect 725 370 775 420
rect 125 270 175 320
rect 725 270 775 320
rect 125 170 175 220
rect 725 170 775 220
<< poly2cap >>
rect 225 1180 675 1240
rect 225 1130 275 1180
rect 325 1130 430 1180
rect 480 1130 575 1180
rect 625 1130 675 1180
rect 225 1070 675 1130
rect 225 1020 275 1070
rect 325 1020 430 1070
rect 480 1020 575 1070
rect 625 1020 675 1070
rect 225 960 675 1020
rect 225 910 275 960
rect 325 910 430 960
rect 480 910 575 960
rect 625 910 675 960
rect 225 850 675 910
rect 225 800 275 850
rect 325 800 430 850
rect 480 800 575 850
rect 625 800 675 850
rect 225 740 675 800
rect 225 690 275 740
rect 325 690 430 740
rect 480 690 575 740
rect 625 690 675 740
rect 225 630 675 690
rect 225 580 275 630
rect 325 580 430 630
rect 480 580 575 630
rect 625 580 675 630
rect 225 520 675 580
rect 225 470 275 520
rect 325 470 430 520
rect 480 470 575 520
rect 625 470 675 520
rect 225 410 675 470
rect 225 360 275 410
rect 325 360 430 410
rect 480 360 575 410
rect 625 360 675 410
rect 225 300 675 360
rect 225 250 275 300
rect 325 250 430 300
rect 480 250 575 300
rect 625 250 675 300
rect 225 200 675 250
<< poly2capcontact >>
rect 275 1130 325 1180
rect 430 1130 480 1180
rect 575 1130 625 1180
rect 275 1020 325 1070
rect 430 1020 480 1070
rect 575 1020 625 1070
rect 275 910 325 960
rect 430 910 480 960
rect 575 910 625 960
rect 275 800 325 850
rect 430 800 480 850
rect 575 800 625 850
rect 275 690 325 740
rect 430 690 480 740
rect 575 690 625 740
rect 275 580 325 630
rect 430 580 480 630
rect 575 580 625 630
rect 275 470 325 520
rect 430 470 480 520
rect 575 470 625 520
rect 275 360 325 410
rect 430 360 480 410
rect 575 360 625 410
rect 275 250 325 300
rect 430 250 480 300
rect 575 250 625 300
<< metal1 >>
rect 0 1395 900 1485
rect 165 1305 735 1395
rect 105 1220 195 1240
rect 105 1170 125 1220
rect 175 1170 195 1220
rect 105 1120 195 1170
rect 105 1070 125 1120
rect 175 1070 195 1120
rect 105 1020 195 1070
rect 105 970 125 1020
rect 175 970 195 1020
rect 105 920 195 970
rect 105 870 125 920
rect 175 870 195 920
rect 105 820 195 870
rect 105 770 125 820
rect 175 770 195 820
rect 105 720 195 770
rect 105 670 125 720
rect 175 670 195 720
rect 105 620 195 670
rect 105 570 125 620
rect 175 570 195 620
rect 105 520 195 570
rect 105 470 125 520
rect 175 470 195 520
rect 105 420 195 470
rect 105 370 125 420
rect 175 370 195 420
rect 105 320 195 370
rect 105 270 125 320
rect 175 270 195 320
rect 105 220 195 270
rect 255 1180 645 1305
rect 255 1130 275 1180
rect 325 1130 430 1180
rect 480 1130 575 1180
rect 625 1130 645 1180
rect 255 1070 645 1130
rect 255 1020 275 1070
rect 325 1020 430 1070
rect 480 1020 575 1070
rect 625 1020 645 1070
rect 255 960 645 1020
rect 255 910 275 960
rect 325 910 430 960
rect 480 910 575 960
rect 625 910 645 960
rect 255 850 645 910
rect 255 800 275 850
rect 325 800 430 850
rect 480 800 575 850
rect 625 800 645 850
rect 255 740 645 800
rect 255 690 275 740
rect 325 690 430 740
rect 480 690 575 740
rect 625 690 645 740
rect 255 630 645 690
rect 255 580 275 630
rect 325 580 430 630
rect 480 580 575 630
rect 625 580 645 630
rect 255 520 645 580
rect 255 470 275 520
rect 325 470 430 520
rect 480 470 575 520
rect 625 470 645 520
rect 255 410 645 470
rect 255 360 275 410
rect 325 360 430 410
rect 480 360 575 410
rect 625 360 645 410
rect 255 300 645 360
rect 255 250 275 300
rect 325 250 430 300
rect 480 250 575 300
rect 625 250 645 300
rect 255 230 645 250
rect 705 1220 795 1240
rect 705 1170 725 1220
rect 775 1170 795 1220
rect 705 1120 795 1170
rect 705 1070 725 1120
rect 775 1070 795 1120
rect 705 1020 795 1070
rect 705 970 725 1020
rect 775 970 795 1020
rect 705 920 795 970
rect 705 870 725 920
rect 775 870 795 920
rect 705 820 795 870
rect 705 770 725 820
rect 775 770 795 820
rect 705 720 795 770
rect 705 670 725 720
rect 775 670 795 720
rect 705 620 795 670
rect 705 570 725 620
rect 775 570 795 620
rect 705 520 795 570
rect 705 470 725 520
rect 775 470 795 520
rect 705 420 795 470
rect 705 370 725 420
rect 775 370 795 420
rect 705 320 795 370
rect 705 270 725 320
rect 775 270 795 320
rect 105 170 125 220
rect 175 170 195 220
rect 105 150 195 170
rect 705 220 795 270
rect 705 170 725 220
rect 775 170 795 220
rect 705 150 795 170
rect 105 45 795 150
rect 0 -45 900 45
<< labels >>
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 0 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 1 ne
flabel nwell 5 580 5 580 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFsite core
string LEFclass CORE
string FIXED_BBOX 0 0 900 1440
string LEFsymmetry X Y
<< end >>
