magic
tech amic5n
timestamp 1608415876
<< nwell >>
rect 3880 590 4500 2090
<< ntransistor >>
rect 7050 410 7110 980
rect 4150 -270 4210 300
rect 7050 -350 7110 220
<< ptransistor >>
rect 4150 740 4210 1940
<< nselect >>
rect 6900 380 7260 1010
rect 4000 -300 4360 330
rect 6900 -380 7260 250
<< pselect >>
rect 4000 710 4360 2010
<< ndiffusion >>
rect 6930 750 7050 980
rect 6930 700 6960 750
rect 7010 700 7050 750
rect 6930 410 7050 700
rect 7110 750 7230 980
rect 7110 700 7150 750
rect 7200 700 7230 750
rect 7110 410 7230 700
rect 4030 10 4150 300
rect 4030 -40 4060 10
rect 4110 -40 4150 10
rect 4030 -270 4150 -40
rect 4210 10 4330 300
rect 4210 -40 4250 10
rect 4300 -40 4330 10
rect 4210 -270 4330 -40
rect 6930 -70 7050 220
rect 6930 -120 6960 -70
rect 7010 -120 7050 -70
rect 6930 -350 7050 -120
rect 7110 -70 7230 220
rect 7110 -120 7150 -70
rect 7200 -120 7230 -70
rect 7110 -350 7230 -120
<< pdiffusion >>
rect 4030 1310 4150 1940
rect 4030 1260 4060 1310
rect 4110 1260 4150 1310
rect 4030 740 4150 1260
rect 4210 1310 4330 1940
rect 4210 1260 4250 1310
rect 4300 1260 4330 1310
rect 4210 740 4330 1260
<< ndcontact >>
rect 6960 700 7010 750
rect 7150 700 7200 750
rect 4060 -40 4110 10
rect 4250 -40 4300 10
rect 6960 -120 7010 -70
rect 7150 -120 7200 -70
<< pdcontact >>
rect 4060 1260 4110 1310
rect 4250 1260 4300 1310
<< polysilicon >>
rect 4150 1940 4210 2005
rect 7050 980 7110 1050
rect 4150 480 4210 740
rect 4040 460 4210 480
rect 4040 410 4060 460
rect 4110 410 4210 460
rect 4040 390 4210 410
rect 4150 300 4210 390
rect 7050 345 7110 410
rect 7050 220 7110 285
rect 4150 -335 4210 -270
rect 7050 -420 7110 -350
<< polycontact >>
rect 4060 410 4110 460
<< metal1 >>
rect 5030 2540 5120 2560
rect 5030 2490 5050 2540
rect 5100 2490 5120 2540
rect 5030 2220 5120 2490
rect 5030 2170 5050 2220
rect 5100 2170 5120 2220
rect 4040 1990 4320 2080
rect 4040 1310 4130 1990
rect 5030 1900 5120 2170
rect 5030 1850 5050 1900
rect 5100 1850 5120 1900
rect 5030 1580 5120 1850
rect 5030 1530 5050 1580
rect 5100 1530 5120 1580
rect 4040 1260 4060 1310
rect 4110 1260 4130 1310
rect 4040 750 4130 1260
rect 4230 1310 4320 1330
rect 4230 1260 4250 1310
rect 4300 1260 4320 1310
rect 4040 460 4130 480
rect 4040 410 4060 460
rect 4110 410 4130 460
rect 4040 390 4130 410
rect 4040 10 4130 290
rect 4040 -40 4060 10
rect 4110 -40 4130 10
rect 4040 -320 4130 -40
rect 4230 10 4320 1260
rect 4230 -40 4250 10
rect 4300 -40 4320 10
rect 4230 -60 4320 -40
rect 5030 1260 5120 1530
rect 5030 1210 5050 1260
rect 5100 1210 5120 1260
rect 5030 940 5120 1210
rect 5030 890 5050 940
rect 5100 890 5120 940
rect 5030 620 5120 890
rect 5030 570 5050 620
rect 5100 570 5120 620
rect 5030 300 5120 570
rect 5030 250 5050 300
rect 5100 250 5120 300
rect 5030 -20 5120 250
rect 5030 -70 5050 -20
rect 5100 -70 5120 -20
rect 4040 -410 4320 -320
rect 5030 -340 5120 -70
rect 5030 -390 5050 -340
rect 5100 -390 5120 -340
rect 5030 -500 5120 -390
rect 5030 -550 5050 -500
rect 5100 -550 5120 -500
rect 5030 -820 5120 -550
rect 5030 -870 5050 -820
rect 5100 -870 5120 -820
rect 5030 -1140 5120 -870
rect 5030 -1190 5050 -1140
rect 5100 -1190 5120 -1140
rect 5030 -1210 5120 -1190
rect 5180 2380 5270 2560
rect 5180 2330 5200 2380
rect 5250 2330 5270 2380
rect 5180 2060 5270 2330
rect 5180 2010 5200 2060
rect 5250 2010 5270 2060
rect 5180 1740 5270 2010
rect 5180 1690 5200 1740
rect 5250 1690 5270 1740
rect 5180 1420 5270 1690
rect 5180 1370 5200 1420
rect 5250 1370 5270 1420
rect 5180 1100 5270 1370
rect 5180 1050 5200 1100
rect 5250 1050 5270 1100
rect 5180 780 5270 1050
rect 5180 730 5200 780
rect 5250 730 5270 780
rect 5180 460 5270 730
rect 6940 750 7030 770
rect 6940 700 6960 750
rect 7010 700 7030 750
rect 6940 680 7030 700
rect 7130 750 7220 770
rect 7130 700 7150 750
rect 7200 700 7220 750
rect 5180 410 5200 460
rect 5250 410 5270 460
rect 5180 140 5270 410
rect 5180 90 5200 140
rect 5250 90 5270 140
rect 5180 -180 5270 90
rect 6940 -70 7030 -50
rect 6940 -120 6960 -70
rect 7010 -120 7030 -70
rect 6940 -140 7030 -120
rect 7130 -70 7220 700
rect 7130 -120 7150 -70
rect 7200 -120 7220 -70
rect 7130 -140 7220 -120
rect 5180 -230 5200 -180
rect 5250 -230 5270 -180
rect 5180 -660 5270 -230
rect 5180 -710 5200 -660
rect 5250 -710 5270 -660
rect 5180 -980 5270 -710
rect 5180 -1030 5200 -980
rect 5250 -1030 5270 -980
rect 5180 -1210 5270 -1030
<< via1 >>
rect 5050 2490 5100 2540
rect 5050 2170 5100 2220
rect 5050 1850 5100 1900
rect 5050 1530 5100 1580
rect 5050 1210 5100 1260
rect 5050 890 5100 940
rect 5050 570 5100 620
rect 5050 250 5100 300
rect 5050 -70 5100 -20
rect 5050 -390 5100 -340
rect 5050 -550 5100 -500
rect 5050 -870 5100 -820
rect 5050 -1190 5100 -1140
rect 5200 2330 5250 2380
rect 5200 2010 5250 2060
rect 5200 1690 5250 1740
rect 5200 1370 5250 1420
rect 5200 1050 5250 1100
rect 5200 730 5250 780
rect 5200 410 5250 460
rect 5200 90 5250 140
rect 5200 -230 5250 -180
rect 5200 -710 5250 -660
rect 5200 -1030 5250 -980
<< metal2 >>
rect 4710 2540 5730 2560
rect 4710 2490 5050 2540
rect 5100 2490 5730 2540
rect 4710 2470 5730 2490
rect 4710 2380 5730 2400
rect 4710 2330 5200 2380
rect 5250 2330 5730 2380
rect 4710 2310 5730 2330
rect 4710 2220 5730 2240
rect 4710 2170 5050 2220
rect 5100 2170 5730 2220
rect 4710 2150 5730 2170
rect 4710 2060 5730 2080
rect 4710 2010 5200 2060
rect 5250 2010 5730 2060
rect 4710 1990 5730 2010
rect 4710 1900 5730 1920
rect 4710 1850 5050 1900
rect 5100 1850 5730 1900
rect 4710 1830 5730 1850
rect 4710 1740 5730 1760
rect 4710 1690 5200 1740
rect 5250 1690 5730 1740
rect 4710 1670 5730 1690
rect 4710 1580 5730 1600
rect 4710 1530 5050 1580
rect 5100 1530 5730 1580
rect 4710 1510 5730 1530
rect 4710 1420 5730 1440
rect 4710 1370 5200 1420
rect 5250 1370 5730 1420
rect 4710 1350 5730 1370
rect 4710 1260 5730 1280
rect 4710 1210 5050 1260
rect 5100 1210 5730 1260
rect 4710 1190 5730 1210
rect 4710 1100 5730 1120
rect 4710 1050 5200 1100
rect 5250 1050 5730 1100
rect 4710 1030 5730 1050
rect 4710 940 5730 960
rect 4710 890 5050 940
rect 5100 890 5730 940
rect 4710 870 5730 890
rect 4710 780 5730 800
rect 4710 730 5200 780
rect 5250 730 5730 780
rect 4710 710 5730 730
rect 4710 620 5730 640
rect 4710 570 5050 620
rect 5100 570 5730 620
rect 4710 550 5730 570
rect 4710 460 5730 480
rect 4710 410 5200 460
rect 5250 410 5730 460
rect 4710 390 5730 410
rect 4710 300 5730 320
rect 4710 250 5050 300
rect 5100 250 5730 300
rect 6790 270 7050 360
rect 4710 230 5730 250
rect 4710 140 5730 160
rect 4710 90 5200 140
rect 5250 90 5730 140
rect 4710 70 5730 90
rect 4710 -20 5730 0
rect 4710 -70 5050 -20
rect 5100 -70 5730 -20
rect 4710 -90 5730 -70
rect 4710 -180 5730 -160
rect 4710 -230 5200 -180
rect 5250 -230 5730 -180
rect 4710 -250 5730 -230
rect 4710 -340 5730 -320
rect 4710 -390 5050 -340
rect 5100 -390 5730 -340
rect 4710 -410 5730 -390
rect 4710 -500 5730 -480
rect 4710 -550 5050 -500
rect 5100 -550 5730 -500
rect 4710 -570 5730 -550
rect 4710 -660 5730 -640
rect 4710 -710 5200 -660
rect 5250 -710 5730 -660
rect 4710 -730 5730 -710
rect 4710 -820 5730 -800
rect 4710 -870 5050 -820
rect 5100 -870 5730 -820
rect 4710 -890 5730 -870
rect 4710 -980 5730 -960
rect 4710 -1030 5200 -980
rect 5250 -1030 5730 -980
rect 4710 -1050 5730 -1030
rect 4710 -1140 5730 -1120
rect 4710 -1190 5050 -1140
rect 5100 -1190 5730 -1140
rect 4710 -1210 5730 -1190
<< labels >>
flabel metal1 s 4260 360 4260 360 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 4060 -390 4060 -390 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel nwell 4350 640 4350 640 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 4050 2010 4050 2010 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 4060 400 4060 400 2 FreeSans 400 0 0 0 a
port 2 ne
<< end >>
