magic
tech scmos
timestamp 1540770671
<< nwell >>
rect -12 39 108 81
rect 116 30 175 81
<< ntransistor >>
rect -1 4 1 14
rect 7 4 9 14
rect 15 4 17 14
rect 20 4 22 14
rect 29 4 31 14
rect 34 4 36 14
rect 43 4 45 14
rect 59 4 61 14
rect 64 4 66 14
rect 74 4 76 14
rect 79 4 81 14
rect 87 4 89 14
rect 95 4 97 14
rect 141 4 143 24
<< ptransistor >>
rect -1 55 1 75
rect 7 55 9 75
rect 15 55 17 75
rect 21 55 23 75
rect 29 55 31 75
rect 35 55 37 75
rect 43 55 45 75
rect 59 55 61 75
rect 64 55 66 75
rect 74 65 76 75
rect 79 65 81 75
rect 87 55 89 75
rect 95 55 97 75
rect 140 36 142 75
rect 149 36 151 75
<< ndiffusion >>
rect -2 4 -1 14
rect 1 6 2 14
rect 6 6 7 14
rect 1 4 7 6
rect 9 4 10 14
rect 14 4 15 14
rect 17 4 20 14
rect 22 13 29 14
rect 22 6 24 13
rect 28 6 29 13
rect 22 4 29 6
rect 31 4 34 14
rect 36 13 43 14
rect 36 4 37 13
rect 41 4 43 13
rect 45 13 50 14
rect 45 6 46 13
rect 45 4 50 6
rect 54 13 59 14
rect 58 4 59 13
rect 61 4 64 14
rect 66 13 74 14
rect 66 6 68 13
rect 72 6 74 13
rect 66 4 74 6
rect 76 4 79 14
rect 81 4 82 14
rect 86 4 87 14
rect 89 6 90 14
rect 94 6 95 14
rect 89 4 95 6
rect 97 4 98 14
rect 102 4 103 14
rect 137 4 141 24
rect 143 4 147 24
<< pdiffusion >>
rect -2 55 -1 75
rect 1 73 7 75
rect 1 55 2 73
rect 6 55 7 73
rect 9 55 10 75
rect 14 55 15 75
rect 17 55 21 75
rect 23 73 29 75
rect 23 55 24 73
rect 28 55 29 73
rect 31 55 35 75
rect 37 74 43 75
rect 37 55 38 74
rect 42 55 43 74
rect 45 73 50 75
rect 45 55 46 73
rect 54 74 59 75
rect 58 55 59 74
rect 61 55 64 75
rect 66 73 74 75
rect 66 55 68 73
rect 72 65 74 73
rect 76 65 79 75
rect 81 74 87 75
rect 81 65 82 74
rect 72 55 73 65
rect 86 55 87 74
rect 89 73 95 75
rect 89 55 90 73
rect 94 55 95 73
rect 97 74 102 75
rect 97 55 98 74
rect 134 36 140 75
rect 142 36 149 75
rect 151 36 158 75
<< ndcontact >>
rect -6 4 -2 14
rect 2 6 6 14
rect 10 4 14 14
rect 24 6 28 13
rect 37 4 41 13
rect 46 6 50 13
rect 54 4 58 13
rect 68 6 72 13
rect 82 4 86 14
rect 90 6 94 14
rect 98 4 102 14
<< pdcontact >>
rect -6 55 -2 75
rect 2 55 6 73
rect 10 55 14 75
rect 24 55 28 73
rect 38 55 42 74
rect 46 55 50 73
rect 54 55 58 74
rect 68 55 72 73
rect 82 55 86 74
rect 90 55 94 73
rect 98 55 102 74
<< polysilicon >>
rect -1 75 1 77
rect 7 75 9 77
rect 15 75 17 77
rect 21 75 23 77
rect 29 75 31 77
rect 35 75 37 77
rect 43 75 45 77
rect 59 75 61 77
rect 64 75 66 77
rect 74 75 76 77
rect 79 75 81 77
rect 87 75 89 77
rect 95 75 97 77
rect 140 75 142 77
rect 149 75 151 77
rect -1 54 1 55
rect 7 54 9 55
rect -1 52 9 54
rect 7 24 9 52
rect 15 38 17 55
rect 21 38 23 55
rect 29 45 31 55
rect 27 41 31 45
rect 14 34 18 38
rect 21 34 25 38
rect 7 20 12 24
rect 7 18 9 20
rect -1 16 9 18
rect -1 14 1 16
rect 7 14 9 16
rect 15 14 17 34
rect 29 29 31 41
rect 35 38 37 55
rect 43 52 45 55
rect 59 54 61 55
rect 41 48 45 52
rect 35 34 39 38
rect 20 27 31 29
rect 20 14 22 27
rect 27 20 31 24
rect 29 14 31 20
rect 34 20 39 24
rect 34 14 36 20
rect 43 14 45 48
rect 49 52 61 54
rect 49 38 51 52
rect 64 45 66 55
rect 61 41 66 45
rect 49 34 53 38
rect 49 17 51 34
rect 64 32 66 41
rect 55 27 59 31
rect 64 30 71 32
rect 57 25 59 27
rect 57 23 66 25
rect 49 15 61 17
rect 59 14 61 15
rect 64 14 66 23
rect 69 17 71 30
rect 74 31 76 65
rect 79 38 81 65
rect 87 54 89 55
rect 95 54 97 55
rect 87 52 97 54
rect 87 45 89 52
rect 83 41 89 45
rect 79 34 83 38
rect 74 27 78 31
rect 79 20 83 24
rect 69 15 76 17
rect 74 14 76 15
rect 79 14 81 20
rect 87 17 89 41
rect 140 34 142 36
rect 149 34 151 36
rect 141 24 143 30
rect 87 15 97 17
rect 87 14 89 15
rect 95 14 97 15
rect -1 2 1 4
rect 7 2 9 4
rect 15 2 17 4
rect 20 2 22 4
rect 29 2 31 4
rect 34 2 36 4
rect 43 2 45 4
rect 59 2 61 4
rect 64 2 66 4
rect 74 2 76 4
rect 79 2 81 4
rect 87 2 89 4
rect 95 2 97 4
rect 141 2 143 4
<< genericcontact >>
rect 42 49 44 51
rect 28 42 30 44
rect 62 42 64 44
rect 84 42 86 44
rect 15 35 17 37
rect 22 35 24 37
rect 36 35 38 37
rect 50 35 52 37
rect 80 35 82 37
rect 56 28 58 30
rect 75 28 77 30
rect 9 21 11 23
rect 28 21 30 23
rect 36 21 38 23
rect 80 21 82 23
<< metal1 >>
rect -6 76 102 79
rect 120 76 171 79
rect -6 75 -2 76
rect 10 75 14 76
rect 38 74 42 76
rect 54 74 58 76
rect 82 74 86 76
rect 98 74 102 76
rect 120 62 131 66
rect 161 62 171 66
rect 120 55 131 59
rect 161 55 171 59
rect 2 45 6 55
rect 24 48 45 52
rect 2 41 65 45
rect 68 41 87 45
rect 2 39 6 41
rect 2 16 5 39
rect 10 34 18 38
rect 21 34 31 38
rect 35 34 53 38
rect 79 37 83 38
rect 90 37 94 55
rect 120 48 131 52
rect 161 48 171 52
rect 120 41 131 45
rect 161 41 171 45
rect 79 34 94 37
rect 120 34 131 38
rect 161 34 171 38
rect 27 31 31 34
rect 27 27 78 31
rect 27 24 31 27
rect 90 24 94 34
rect 120 27 131 31
rect 161 27 171 31
rect 8 20 31 24
rect 35 20 49 24
rect 79 20 94 24
rect 120 20 129 24
rect 160 20 171 24
rect 2 14 6 16
rect 46 14 49 20
rect 90 14 94 20
rect -6 3 -2 4
rect 24 13 28 14
rect 37 13 42 14
rect 10 3 14 4
rect 41 4 42 13
rect 46 13 50 14
rect 54 13 58 14
rect 37 3 42 4
rect 68 13 72 14
rect 54 3 58 4
rect 82 3 86 4
rect 120 13 129 17
rect 160 13 171 17
rect 120 6 129 10
rect 160 6 171 10
rect 98 3 102 4
rect -12 0 102 3
rect 120 0 171 3
<< metal2 >>
rect 24 9 28 68
rect 46 6 50 63
rect 68 8 72 63
<< gv1 >>
rect 25 59 27 61
rect 47 58 49 60
rect 69 58 71 60
rect 25 49 27 51
rect 69 42 71 44
rect 47 35 49 37
rect 25 10 27 12
rect 47 8 49 10
rect 69 9 71 11
<< labels >>
rlabel ndiffusion s 18 8 18 8 2 x5
rlabel ndiffusion s 32 8 32 8 2 x6
rlabel ndiffusion s 62 7 62 7 2 x7
rlabel ndiffusion s 77 7 77 7 2 x8
rlabel ndiffusion s 2 8 2 8 2 x5
rlabel metal1 120 0 120 0 2 Gnd
port 3 ne
rlabel nwell 120 30 120 30 2 Vdd
rlabel metal1 s 34 28 34 28 2 CLK
port 3 ne
rlabel metal1 s 12 36 12 36 2 D
port 2 ne
rlabel metal1 91 40 91 40 2 Q
port 1 ne
rlabel metal1 12 42 12 42 2 NCLK
rlabel metal1 s 35 49 35 49 2 MAS
rlabel metal1 s 78 43 78 43 2 SLV
rlabel metal1 120 76 120 76 2 Vdd
port 2 ne
rlabel metal1 s 40 36 40 36 2 n1
rlabel pdiffusion s 19 65 19 65 2 x1
rlabel pdiffusion s 32 65 32 65 2 x2
rlabel pdiffusion s 62 65 62 65 2 x3
rlabel pdiffusion s 77 69 77 69 2 x4
rlabel metal1 11 76 11 76 2 Vdd
port 2 ne
rlabel nwell -7 43 -7 43 2 Vdd
<< end >>
