magic
tech amic5n
timestamp 1608317707
<< nwell >>
rect -90 870 2250 2430
<< nselect >>
rect 0 60 2160 750
<< pselect >>
rect 30 990 2130 2310
<< ntransistor >>
rect 210 120 270 690
rect 450 120 510 690
rect 690 120 750 690
rect 930 120 990 690
rect 1170 120 1230 690
rect 1410 120 1470 690
rect 1650 120 1710 690
rect 1890 120 1950 690
<< ptransistor >>
rect 240 1050 300 2250
rect 450 1050 510 2250
rect 690 1050 750 2250
rect 900 1050 960 2250
rect 1200 1050 1260 2250
rect 1410 1050 1470 2250
rect 1650 1050 1710 2250
rect 1860 1050 1920 2250
<< ndiffusion >>
rect 60 120 210 690
rect 270 120 450 690
rect 510 120 690 690
rect 750 120 930 690
rect 990 120 1170 690
rect 1230 120 1410 690
rect 1470 120 1650 690
rect 1710 120 1890 690
rect 1950 120 2100 690
<< pdiffusion >>
rect 90 1050 240 2250
rect 300 1050 450 2250
rect 510 1050 690 2250
rect 750 1050 900 2250
rect 960 1050 1200 2250
rect 1260 1050 1410 2250
rect 1470 1050 1650 2250
rect 1710 1050 1860 2250
rect 1920 1050 2070 2250
<< polysilicon >>
rect 240 2250 300 2310
rect 450 2250 510 2310
rect 690 2250 750 2310
rect 900 2250 960 2310
rect 1200 2250 1260 2310
rect 1410 2250 1470 2310
rect 1650 2250 1710 2310
rect 1860 2250 1920 2310
rect 240 960 300 1050
rect 60 780 300 960
rect 450 960 510 1050
rect 690 960 750 1050
rect 450 780 750 960
rect 900 960 960 1050
rect 1200 960 1260 1050
rect 900 780 1260 960
rect 1410 960 1470 1050
rect 1650 960 1710 1050
rect 1410 780 1710 960
rect 1860 960 1920 1050
rect 1860 780 2100 960
rect 210 690 270 780
rect 450 690 510 780
rect 690 690 750 780
rect 930 690 990 780
rect 1170 690 1230 780
rect 1410 690 1470 780
rect 1650 690 1710 780
rect 1890 690 1950 780
rect 210 60 270 120
rect 450 60 510 120
rect 690 60 750 120
rect 930 60 990 120
rect 1170 60 1230 120
rect 1410 60 1470 120
rect 1650 60 1710 120
rect 1890 60 1950 120
<< pdcontact >>
rect 125 2165 175 2215
<< pdcontact >>
rect 1055 2165 1105 2215
<< pdcontact >>
rect 1985 2165 2035 2215
<< pdcontact >>
rect 575 2105 625 2155
<< pdcontact >>
rect 1535 2105 1585 2155
<< pdcontact >>
rect 125 1985 175 2035
<< pdcontact >>
rect 575 1955 625 2005
<< pdcontact >>
rect 1055 1985 1105 2035
<< pdcontact >>
rect 1535 1955 1585 2005
<< pdcontact >>
rect 1985 1985 2035 2035
<< pdcontact >>
rect 125 1835 175 1885
<< pdcontact >>
rect 1055 1835 1105 1885
<< pdcontact >>
rect 1985 1835 2035 1885
<< pdcontact >>
rect 575 1775 625 1825
<< pdcontact >>
rect 1535 1775 1585 1825
<< pdcontact >>
rect 125 1685 175 1735
<< pdcontact >>
rect 1055 1685 1105 1735
<< pdcontact >>
rect 1985 1685 2035 1735
<< pdcontact >>
rect 575 1595 625 1645
<< pdcontact >>
rect 1535 1595 1585 1645
<< pdcontact >>
rect 125 1535 175 1585
<< pdcontact >>
rect 1055 1535 1105 1585
<< pdcontact >>
rect 1985 1535 2035 1585
<< pdcontact >>
rect 125 1385 175 1435
<< pdcontact >>
rect 575 1415 625 1465
<< pdcontact >>
rect 1055 1385 1105 1435
<< pdcontact >>
rect 1535 1415 1585 1465
<< pdcontact >>
rect 1985 1385 2035 1435
<< pdcontact >>
rect 125 1235 175 1285
<< pdcontact >>
rect 575 1235 625 1285
<< pdcontact >>
rect 1055 1235 1105 1285
<< pdcontact >>
rect 1535 1235 1585 1285
<< pdcontact >>
rect 1985 1235 2035 1285
<< pdcontact >>
rect 125 1085 175 1135
<< pdcontact >>
rect 575 1085 625 1135
<< pdcontact >>
rect 1055 1085 1105 1135
<< pdcontact >>
rect 1535 1085 1585 1135
<< pdcontact >>
rect 1985 1085 2035 1135
<< polycontact >>
rect 125 845 175 895
<< polycontact >>
rect 575 845 625 895
<< polycontact >>
rect 1055 845 1105 895
<< polycontact >>
rect 1535 845 1585 895
<< polycontact >>
rect 1985 845 2035 895
<< ndcontact >>
rect 95 605 145 655
<< ndcontact >>
rect 335 605 385 655
<< ndcontact >>
rect 575 605 625 655
<< ndcontact >>
rect 815 605 865 655
<< ndcontact >>
rect 1055 605 1105 655
<< ndcontact >>
rect 1295 605 1345 655
<< ndcontact >>
rect 1535 605 1585 655
<< ndcontact >>
rect 1775 605 1825 655
<< ndcontact >>
rect 2015 605 2065 655
<< ndcontact >>
rect 95 455 145 505
<< ndcontact >>
rect 575 455 625 505
<< ndcontact >>
rect 1055 455 1105 505
<< ndcontact >>
rect 1535 455 1585 505
<< ndcontact >>
rect 2015 455 2065 505
<< ndcontact >>
rect 335 395 385 445
<< ndcontact >>
rect 815 395 865 445
<< ndcontact >>
rect 1295 395 1345 445
<< ndcontact >>
rect 1775 395 1825 445
<< ndcontact >>
rect 95 305 145 355
<< ndcontact >>
rect 575 305 625 355
<< ndcontact >>
rect 1055 305 1105 355
<< ndcontact >>
rect 1535 305 1585 355
<< ndcontact >>
rect 2015 305 2065 355
<< ndcontact >>
rect 335 215 385 265
<< ndcontact >>
rect 815 215 865 265
<< ndcontact >>
rect 1295 215 1345 265
<< ndcontact >>
rect 1775 215 1825 265
<< ndcontact >>
rect 95 155 145 205
<< ndcontact >>
rect 575 155 625 205
<< ndcontact >>
rect 1055 155 1105 205
<< ndcontact >>
rect 1535 155 1585 205
<< ndcontact >>
rect 2015 155 2065 205
<< metal1 >>
rect 0 2280 2160 2370
rect 90 1050 210 2280
rect 540 1200 660 2190
rect 300 1050 900 1200
rect 1020 1050 1140 2280
rect 1500 1200 1620 2190
rect 1260 1050 1860 1200
rect 1950 1050 2070 2280
rect 90 810 210 930
rect 60 90 180 690
rect 300 180 420 1050
rect 510 810 690 930
rect 540 90 660 690
rect 780 180 900 1050
rect 1020 810 1140 930
rect 1020 90 1140 690
rect 1260 180 1380 1050
rect 1470 810 1650 930
rect 1500 90 1620 690
rect 1740 180 1860 1050
rect 1950 810 2070 930
rect 1980 90 2100 690
rect 0 0 2160 90
<< metal2 >>
rect 540 1230 1620 1350
rect 540 1020 1620 1140
rect 90 720 210 930
rect 540 810 660 1020
rect 1020 720 1140 930
rect 1500 810 1620 1020
rect 1950 720 2070 930
rect 90 600 2070 720
<< via1 >>
rect 575 1265 625 1315
rect 1535 1265 1585 1315
rect 125 845 175 895
rect 575 845 625 895
rect 1055 845 1105 895
rect 1535 845 1585 895
rect 1985 845 2035 895
<< labels >>
flabel metal1 s 30 30 30 30 2 FreeSans 400 0 0 0 vss
port 5 ne
flabel metal1 s 30 2310 30 2310 2 FreeSans 400 0 0 0 vdd
port 4 ne
flabel metal1 s 570 870 570 870 2 FreeSans 400 0 0 0 b
port 3 ne
flabel metal1 s 150 870 150 870 2 FreeSans 400 0 0 0 a
port 2 ne
flabel metal1 s 360 780 360 780 2 FreeSans 400 0 0 0 z
port 1 ne
flabel nwell  0 930 0 930 2 FreeSans 400 0 0 0 vdd
flabel ndiffusion s 330 1260 330 1260 2 FreeSans 400 0 0 0 x1
flabel ndiffusion s 780 1260 780 1260 2 FreeSans 400 0 0 0 x2
flabel ndiffusion s 1290 1260 1290 1260 2 FreeSans 400 0 0 0 x3
flabel ndiffusion s 1740 1260 1740 1260 2 FreeSans 400 0 0 0 x4
<< checkpaint >>
rect -100 -10 2260 2440
<< end >>
