magic
tech amic5n
timestamp 1608317708
<< metal1 >>
rect 0 0 3000000 3000000
<< labels >>
flabel metal1 s 12300 12300 12300 12300 2 FreeSans 400 0 0 0 node_a
<< checkpaint >>
rect -10 -10 3000010 3000010
<< end >>
