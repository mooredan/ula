magic
tech amic5n
timestamp 1624549694
<< nwell >>
rect -130 550 280 1495
<< nselect >>
rect -10 0 160 430
<< pselect >>
rect -10 670 160 1440
<< metal1 >>
rect 0 1395 150 1485
rect 0 -45 150 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 1 ne
flabel metal1 s 20 1415 20 1415 2 FreeSans 400 0 0 0 vdd
port 0 ne
flabel nwell 95 600 95 600 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
<< end >>
