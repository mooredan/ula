magic
tech scmos
timestamp 1570494029
<< error_s >>
rect 35 230 39 231
rect 35 228 36 230
rect 38 228 39 230
rect 35 227 39 228
rect 47 230 51 231
rect 47 228 48 230
rect 50 228 51 230
rect 47 227 51 228
rect 59 230 63 231
rect 59 228 60 230
rect 62 228 63 230
rect 59 227 63 228
rect 71 230 75 231
rect 71 228 72 230
rect 74 228 75 230
rect 71 227 75 228
rect 83 230 87 231
rect 83 228 84 230
rect 86 228 87 230
rect 83 227 87 228
rect 95 230 99 231
rect 95 228 96 230
rect 98 228 99 230
rect 95 227 99 228
rect 107 230 111 231
rect 107 228 108 230
rect 110 228 111 230
rect 107 227 111 228
rect 119 230 123 231
rect 119 228 120 230
rect 122 228 123 230
rect 119 227 123 228
rect 131 230 135 231
rect 131 228 132 230
rect 134 228 135 230
rect 131 227 135 228
rect 143 230 147 231
rect 143 228 144 230
rect 146 228 147 230
rect 143 227 147 228
rect 155 230 159 231
rect 155 228 156 230
rect 158 228 159 230
rect 155 227 159 228
rect 167 230 171 231
rect 167 228 168 230
rect 170 228 171 230
rect 167 227 171 228
rect 179 230 183 231
rect 179 228 180 230
rect 182 228 183 230
rect 179 227 183 228
rect 191 230 195 231
rect 191 228 192 230
rect 194 228 195 230
rect 191 227 195 228
rect 203 230 207 231
rect 203 228 204 230
rect 206 228 207 230
rect 203 227 207 228
rect 215 230 219 231
rect 215 228 216 230
rect 218 228 219 230
rect 215 227 219 228
rect 227 230 231 231
rect 227 228 228 230
rect 230 228 231 230
rect 227 227 231 228
rect 29 224 33 225
rect 29 222 30 224
rect 32 222 33 224
rect 29 221 33 222
rect 41 224 45 225
rect 41 222 42 224
rect 44 222 45 224
rect 41 221 45 222
rect 53 224 57 225
rect 53 222 54 224
rect 56 222 57 224
rect 53 221 57 222
rect 65 224 69 225
rect 65 222 66 224
rect 68 222 69 224
rect 65 221 69 222
rect 77 224 81 225
rect 77 222 78 224
rect 80 222 81 224
rect 77 221 81 222
rect 89 224 93 225
rect 89 222 90 224
rect 92 222 93 224
rect 89 221 93 222
rect 101 224 105 225
rect 101 222 102 224
rect 104 222 105 224
rect 101 221 105 222
rect 113 224 117 225
rect 113 222 114 224
rect 116 222 117 224
rect 113 221 117 222
rect 125 224 129 225
rect 125 222 126 224
rect 128 222 129 224
rect 125 221 129 222
rect 137 224 141 225
rect 137 222 138 224
rect 140 222 141 224
rect 137 221 141 222
rect 149 224 153 225
rect 149 222 150 224
rect 152 222 153 224
rect 149 221 153 222
rect 161 224 165 225
rect 161 222 162 224
rect 164 222 165 224
rect 161 221 165 222
rect 173 224 177 225
rect 173 222 174 224
rect 176 222 177 224
rect 173 221 177 222
rect 185 224 189 225
rect 185 222 186 224
rect 188 222 189 224
rect 185 221 189 222
rect 197 224 201 225
rect 197 222 198 224
rect 200 222 201 224
rect 197 221 201 222
rect 209 224 213 225
rect 209 222 210 224
rect 212 222 213 224
rect 209 221 213 222
rect 221 224 225 225
rect 221 222 222 224
rect 224 222 225 224
rect 221 221 225 222
rect 35 218 39 219
rect 35 216 36 218
rect 38 216 39 218
rect 35 215 39 216
rect 47 218 51 219
rect 47 216 48 218
rect 50 216 51 218
rect 47 215 51 216
rect 59 218 63 219
rect 59 216 60 218
rect 62 216 63 218
rect 59 215 63 216
rect 71 218 75 219
rect 71 216 72 218
rect 74 216 75 218
rect 71 215 75 216
rect 83 218 87 219
rect 83 216 84 218
rect 86 216 87 218
rect 83 215 87 216
rect 95 218 99 219
rect 95 216 96 218
rect 98 216 99 218
rect 95 215 99 216
rect 107 218 111 219
rect 107 216 108 218
rect 110 216 111 218
rect 107 215 111 216
rect 119 218 123 219
rect 119 216 120 218
rect 122 216 123 218
rect 119 215 123 216
rect 131 218 135 219
rect 131 216 132 218
rect 134 216 135 218
rect 131 215 135 216
rect 143 218 147 219
rect 143 216 144 218
rect 146 216 147 218
rect 143 215 147 216
rect 155 218 159 219
rect 155 216 156 218
rect 158 216 159 218
rect 155 215 159 216
rect 167 218 171 219
rect 167 216 168 218
rect 170 216 171 218
rect 167 215 171 216
rect 179 218 183 219
rect 179 216 180 218
rect 182 216 183 218
rect 179 215 183 216
rect 191 218 195 219
rect 191 216 192 218
rect 194 216 195 218
rect 191 215 195 216
rect 203 218 207 219
rect 203 216 204 218
rect 206 216 207 218
rect 203 215 207 216
rect 215 218 219 219
rect 215 216 216 218
rect 218 216 219 218
rect 215 215 219 216
rect 227 218 231 219
rect 227 216 228 218
rect 230 216 231 218
rect 227 215 231 216
rect 29 212 33 213
rect 29 210 30 212
rect 32 210 33 212
rect 29 209 33 210
rect 41 212 45 213
rect 41 210 42 212
rect 44 210 45 212
rect 41 209 45 210
rect 53 212 57 213
rect 53 210 54 212
rect 56 210 57 212
rect 53 209 57 210
rect 65 212 69 213
rect 65 210 66 212
rect 68 210 69 212
rect 65 209 69 210
rect 77 212 81 213
rect 77 210 78 212
rect 80 210 81 212
rect 77 209 81 210
rect 89 212 93 213
rect 89 210 90 212
rect 92 210 93 212
rect 89 209 93 210
rect 101 212 105 213
rect 101 210 102 212
rect 104 210 105 212
rect 101 209 105 210
rect 113 212 117 213
rect 113 210 114 212
rect 116 210 117 212
rect 113 209 117 210
rect 125 212 129 213
rect 125 210 126 212
rect 128 210 129 212
rect 125 209 129 210
rect 137 212 141 213
rect 137 210 138 212
rect 140 210 141 212
rect 137 209 141 210
rect 149 212 153 213
rect 149 210 150 212
rect 152 210 153 212
rect 149 209 153 210
rect 161 212 165 213
rect 161 210 162 212
rect 164 210 165 212
rect 161 209 165 210
rect 173 212 177 213
rect 173 210 174 212
rect 176 210 177 212
rect 173 209 177 210
rect 185 212 189 213
rect 185 210 186 212
rect 188 210 189 212
rect 185 209 189 210
rect 197 212 201 213
rect 197 210 198 212
rect 200 210 201 212
rect 197 209 201 210
rect 209 212 213 213
rect 209 210 210 212
rect 212 210 213 212
rect 209 209 213 210
rect 221 212 225 213
rect 221 210 222 212
rect 224 210 225 212
rect 221 209 225 210
rect 35 206 39 207
rect 35 204 36 206
rect 38 204 39 206
rect 35 203 39 204
rect 47 206 51 207
rect 47 204 48 206
rect 50 204 51 206
rect 47 203 51 204
rect 59 206 63 207
rect 59 204 60 206
rect 62 204 63 206
rect 59 203 63 204
rect 71 206 75 207
rect 71 204 72 206
rect 74 204 75 206
rect 71 203 75 204
rect 83 206 87 207
rect 83 204 84 206
rect 86 204 87 206
rect 83 203 87 204
rect 95 206 99 207
rect 95 204 96 206
rect 98 204 99 206
rect 95 203 99 204
rect 107 206 111 207
rect 107 204 108 206
rect 110 204 111 206
rect 107 203 111 204
rect 119 206 123 207
rect 119 204 120 206
rect 122 204 123 206
rect 119 203 123 204
rect 131 206 135 207
rect 131 204 132 206
rect 134 204 135 206
rect 131 203 135 204
rect 143 206 147 207
rect 143 204 144 206
rect 146 204 147 206
rect 143 203 147 204
rect 155 206 159 207
rect 155 204 156 206
rect 158 204 159 206
rect 155 203 159 204
rect 167 206 171 207
rect 167 204 168 206
rect 170 204 171 206
rect 167 203 171 204
rect 179 206 183 207
rect 179 204 180 206
rect 182 204 183 206
rect 179 203 183 204
rect 191 206 195 207
rect 191 204 192 206
rect 194 204 195 206
rect 191 203 195 204
rect 203 206 207 207
rect 203 204 204 206
rect 206 204 207 206
rect 203 203 207 204
rect 215 206 219 207
rect 215 204 216 206
rect 218 204 219 206
rect 215 203 219 204
rect 227 206 231 207
rect 227 204 228 206
rect 230 204 231 206
rect 227 203 231 204
rect 29 200 33 201
rect 29 198 30 200
rect 32 198 33 200
rect 29 197 33 198
rect 41 200 45 201
rect 41 198 42 200
rect 44 198 45 200
rect 41 197 45 198
rect 53 200 57 201
rect 53 198 54 200
rect 56 198 57 200
rect 53 197 57 198
rect 65 200 69 201
rect 65 198 66 200
rect 68 198 69 200
rect 65 197 69 198
rect 77 200 81 201
rect 77 198 78 200
rect 80 198 81 200
rect 77 197 81 198
rect 89 200 93 201
rect 89 198 90 200
rect 92 198 93 200
rect 89 197 93 198
rect 101 200 105 201
rect 101 198 102 200
rect 104 198 105 200
rect 101 197 105 198
rect 113 200 117 201
rect 113 198 114 200
rect 116 198 117 200
rect 113 197 117 198
rect 125 200 129 201
rect 125 198 126 200
rect 128 198 129 200
rect 125 197 129 198
rect 137 200 141 201
rect 137 198 138 200
rect 140 198 141 200
rect 137 197 141 198
rect 149 200 153 201
rect 149 198 150 200
rect 152 198 153 200
rect 149 197 153 198
rect 161 200 165 201
rect 161 198 162 200
rect 164 198 165 200
rect 161 197 165 198
rect 173 200 177 201
rect 173 198 174 200
rect 176 198 177 200
rect 173 197 177 198
rect 185 200 189 201
rect 185 198 186 200
rect 188 198 189 200
rect 185 197 189 198
rect 197 200 201 201
rect 197 198 198 200
rect 200 198 201 200
rect 197 197 201 198
rect 209 200 213 201
rect 209 198 210 200
rect 212 198 213 200
rect 209 197 213 198
rect 221 200 225 201
rect 221 198 222 200
rect 224 198 225 200
rect 221 197 225 198
rect 35 194 39 195
rect 35 192 36 194
rect 38 192 39 194
rect 35 191 39 192
rect 47 194 51 195
rect 47 192 48 194
rect 50 192 51 194
rect 47 191 51 192
rect 59 194 63 195
rect 59 192 60 194
rect 62 192 63 194
rect 59 191 63 192
rect 71 194 75 195
rect 71 192 72 194
rect 74 192 75 194
rect 71 191 75 192
rect 83 194 87 195
rect 83 192 84 194
rect 86 192 87 194
rect 83 191 87 192
rect 95 194 99 195
rect 95 192 96 194
rect 98 192 99 194
rect 95 191 99 192
rect 107 194 111 195
rect 107 192 108 194
rect 110 192 111 194
rect 107 191 111 192
rect 119 194 123 195
rect 119 192 120 194
rect 122 192 123 194
rect 119 191 123 192
rect 131 194 135 195
rect 131 192 132 194
rect 134 192 135 194
rect 131 191 135 192
rect 143 194 147 195
rect 143 192 144 194
rect 146 192 147 194
rect 143 191 147 192
rect 155 194 159 195
rect 155 192 156 194
rect 158 192 159 194
rect 155 191 159 192
rect 167 194 171 195
rect 167 192 168 194
rect 170 192 171 194
rect 167 191 171 192
rect 179 194 183 195
rect 179 192 180 194
rect 182 192 183 194
rect 179 191 183 192
rect 191 194 195 195
rect 191 192 192 194
rect 194 192 195 194
rect 191 191 195 192
rect 203 194 207 195
rect 203 192 204 194
rect 206 192 207 194
rect 203 191 207 192
rect 215 194 219 195
rect 215 192 216 194
rect 218 192 219 194
rect 215 191 219 192
rect 227 194 231 195
rect 227 192 228 194
rect 230 192 231 194
rect 227 191 231 192
rect 29 188 33 189
rect 29 186 30 188
rect 32 186 33 188
rect 29 185 33 186
rect 41 188 45 189
rect 41 186 42 188
rect 44 186 45 188
rect 41 185 45 186
rect 53 188 57 189
rect 53 186 54 188
rect 56 186 57 188
rect 53 185 57 186
rect 65 188 69 189
rect 65 186 66 188
rect 68 186 69 188
rect 65 185 69 186
rect 77 188 81 189
rect 77 186 78 188
rect 80 186 81 188
rect 77 185 81 186
rect 89 188 93 189
rect 89 186 90 188
rect 92 186 93 188
rect 89 185 93 186
rect 101 188 105 189
rect 101 186 102 188
rect 104 186 105 188
rect 101 185 105 186
rect 113 188 117 189
rect 113 186 114 188
rect 116 186 117 188
rect 113 185 117 186
rect 125 188 129 189
rect 125 186 126 188
rect 128 186 129 188
rect 125 185 129 186
rect 137 188 141 189
rect 137 186 138 188
rect 140 186 141 188
rect 137 185 141 186
rect 149 188 153 189
rect 149 186 150 188
rect 152 186 153 188
rect 149 185 153 186
rect 161 188 165 189
rect 161 186 162 188
rect 164 186 165 188
rect 161 185 165 186
rect 173 188 177 189
rect 173 186 174 188
rect 176 186 177 188
rect 173 185 177 186
rect 185 188 189 189
rect 185 186 186 188
rect 188 186 189 188
rect 185 185 189 186
rect 197 188 201 189
rect 197 186 198 188
rect 200 186 201 188
rect 197 185 201 186
rect 209 188 213 189
rect 209 186 210 188
rect 212 186 213 188
rect 209 185 213 186
rect 221 188 225 189
rect 221 186 222 188
rect 224 186 225 188
rect 221 185 225 186
rect 35 182 39 183
rect 35 180 36 182
rect 38 180 39 182
rect 35 179 39 180
rect 47 182 51 183
rect 47 180 48 182
rect 50 180 51 182
rect 47 179 51 180
rect 59 182 63 183
rect 59 180 60 182
rect 62 180 63 182
rect 59 179 63 180
rect 71 182 75 183
rect 71 180 72 182
rect 74 180 75 182
rect 71 179 75 180
rect 83 182 87 183
rect 83 180 84 182
rect 86 180 87 182
rect 83 179 87 180
rect 95 182 99 183
rect 95 180 96 182
rect 98 180 99 182
rect 95 179 99 180
rect 107 182 111 183
rect 107 180 108 182
rect 110 180 111 182
rect 107 179 111 180
rect 119 182 123 183
rect 119 180 120 182
rect 122 180 123 182
rect 119 179 123 180
rect 131 182 135 183
rect 131 180 132 182
rect 134 180 135 182
rect 131 179 135 180
rect 143 182 147 183
rect 143 180 144 182
rect 146 180 147 182
rect 143 179 147 180
rect 155 182 159 183
rect 155 180 156 182
rect 158 180 159 182
rect 155 179 159 180
rect 167 182 171 183
rect 167 180 168 182
rect 170 180 171 182
rect 167 179 171 180
rect 179 182 183 183
rect 179 180 180 182
rect 182 180 183 182
rect 179 179 183 180
rect 191 182 195 183
rect 191 180 192 182
rect 194 180 195 182
rect 191 179 195 180
rect 203 182 207 183
rect 203 180 204 182
rect 206 180 207 182
rect 203 179 207 180
rect 215 182 219 183
rect 215 180 216 182
rect 218 180 219 182
rect 215 179 219 180
rect 227 182 231 183
rect 227 180 228 182
rect 230 180 231 182
rect 227 179 231 180
rect 29 176 33 177
rect 29 174 30 176
rect 32 174 33 176
rect 29 173 33 174
rect 41 176 45 177
rect 41 174 42 176
rect 44 174 45 176
rect 41 173 45 174
rect 53 176 57 177
rect 53 174 54 176
rect 56 174 57 176
rect 53 173 57 174
rect 65 176 69 177
rect 65 174 66 176
rect 68 174 69 176
rect 65 173 69 174
rect 77 176 81 177
rect 77 174 78 176
rect 80 174 81 176
rect 77 173 81 174
rect 89 176 93 177
rect 89 174 90 176
rect 92 174 93 176
rect 89 173 93 174
rect 101 176 105 177
rect 101 174 102 176
rect 104 174 105 176
rect 101 173 105 174
rect 113 176 117 177
rect 113 174 114 176
rect 116 174 117 176
rect 113 173 117 174
rect 125 176 129 177
rect 125 174 126 176
rect 128 174 129 176
rect 125 173 129 174
rect 137 176 141 177
rect 137 174 138 176
rect 140 174 141 176
rect 137 173 141 174
rect 149 176 153 177
rect 149 174 150 176
rect 152 174 153 176
rect 149 173 153 174
rect 161 176 165 177
rect 161 174 162 176
rect 164 174 165 176
rect 161 173 165 174
rect 173 176 177 177
rect 173 174 174 176
rect 176 174 177 176
rect 173 173 177 174
rect 185 176 189 177
rect 185 174 186 176
rect 188 174 189 176
rect 185 173 189 174
rect 197 176 201 177
rect 197 174 198 176
rect 200 174 201 176
rect 197 173 201 174
rect 209 176 213 177
rect 209 174 210 176
rect 212 174 213 176
rect 209 173 213 174
rect 221 176 225 177
rect 221 174 222 176
rect 224 174 225 176
rect 221 173 225 174
rect 35 170 39 171
rect 35 168 36 170
rect 38 168 39 170
rect 35 167 39 168
rect 47 170 51 171
rect 47 168 48 170
rect 50 168 51 170
rect 47 167 51 168
rect 59 170 63 171
rect 59 168 60 170
rect 62 168 63 170
rect 59 167 63 168
rect 71 170 75 171
rect 71 168 72 170
rect 74 168 75 170
rect 71 167 75 168
rect 83 170 87 171
rect 83 168 84 170
rect 86 168 87 170
rect 83 167 87 168
rect 95 170 99 171
rect 95 168 96 170
rect 98 168 99 170
rect 95 167 99 168
rect 107 170 111 171
rect 107 168 108 170
rect 110 168 111 170
rect 107 167 111 168
rect 119 170 123 171
rect 119 168 120 170
rect 122 168 123 170
rect 119 167 123 168
rect 131 170 135 171
rect 131 168 132 170
rect 134 168 135 170
rect 131 167 135 168
rect 143 170 147 171
rect 143 168 144 170
rect 146 168 147 170
rect 143 167 147 168
rect 155 170 159 171
rect 155 168 156 170
rect 158 168 159 170
rect 155 167 159 168
rect 167 170 171 171
rect 167 168 168 170
rect 170 168 171 170
rect 167 167 171 168
rect 179 170 183 171
rect 179 168 180 170
rect 182 168 183 170
rect 179 167 183 168
rect 191 170 195 171
rect 191 168 192 170
rect 194 168 195 170
rect 191 167 195 168
rect 203 170 207 171
rect 203 168 204 170
rect 206 168 207 170
rect 203 167 207 168
rect 215 170 219 171
rect 215 168 216 170
rect 218 168 219 170
rect 215 167 219 168
rect 227 170 231 171
rect 227 168 228 170
rect 230 168 231 170
rect 227 167 231 168
rect 29 164 33 165
rect 29 162 30 164
rect 32 162 33 164
rect 29 161 33 162
rect 41 164 45 165
rect 41 162 42 164
rect 44 162 45 164
rect 41 161 45 162
rect 53 164 57 165
rect 53 162 54 164
rect 56 162 57 164
rect 53 161 57 162
rect 65 164 69 165
rect 65 162 66 164
rect 68 162 69 164
rect 65 161 69 162
rect 77 164 81 165
rect 77 162 78 164
rect 80 162 81 164
rect 77 161 81 162
rect 89 164 93 165
rect 89 162 90 164
rect 92 162 93 164
rect 89 161 93 162
rect 101 164 105 165
rect 101 162 102 164
rect 104 162 105 164
rect 101 161 105 162
rect 113 164 117 165
rect 113 162 114 164
rect 116 162 117 164
rect 113 161 117 162
rect 125 164 129 165
rect 125 162 126 164
rect 128 162 129 164
rect 125 161 129 162
rect 137 164 141 165
rect 137 162 138 164
rect 140 162 141 164
rect 137 161 141 162
rect 149 164 153 165
rect 149 162 150 164
rect 152 162 153 164
rect 149 161 153 162
rect 161 164 165 165
rect 161 162 162 164
rect 164 162 165 164
rect 161 161 165 162
rect 173 164 177 165
rect 173 162 174 164
rect 176 162 177 164
rect 173 161 177 162
rect 185 164 189 165
rect 185 162 186 164
rect 188 162 189 164
rect 185 161 189 162
rect 197 164 201 165
rect 197 162 198 164
rect 200 162 201 164
rect 197 161 201 162
rect 209 164 213 165
rect 209 162 210 164
rect 212 162 213 164
rect 209 161 213 162
rect 221 164 225 165
rect 221 162 222 164
rect 224 162 225 164
rect 221 161 225 162
rect 35 158 39 159
rect 35 156 36 158
rect 38 156 39 158
rect 35 155 39 156
rect 47 158 51 159
rect 47 156 48 158
rect 50 156 51 158
rect 47 155 51 156
rect 59 158 63 159
rect 59 156 60 158
rect 62 156 63 158
rect 59 155 63 156
rect 71 158 75 159
rect 71 156 72 158
rect 74 156 75 158
rect 71 155 75 156
rect 83 158 87 159
rect 83 156 84 158
rect 86 156 87 158
rect 83 155 87 156
rect 95 158 99 159
rect 95 156 96 158
rect 98 156 99 158
rect 95 155 99 156
rect 107 158 111 159
rect 107 156 108 158
rect 110 156 111 158
rect 107 155 111 156
rect 119 158 123 159
rect 119 156 120 158
rect 122 156 123 158
rect 119 155 123 156
rect 131 158 135 159
rect 131 156 132 158
rect 134 156 135 158
rect 131 155 135 156
rect 143 158 147 159
rect 143 156 144 158
rect 146 156 147 158
rect 143 155 147 156
rect 155 158 159 159
rect 155 156 156 158
rect 158 156 159 158
rect 155 155 159 156
rect 167 158 171 159
rect 167 156 168 158
rect 170 156 171 158
rect 167 155 171 156
rect 179 158 183 159
rect 179 156 180 158
rect 182 156 183 158
rect 179 155 183 156
rect 191 158 195 159
rect 191 156 192 158
rect 194 156 195 158
rect 191 155 195 156
rect 203 158 207 159
rect 203 156 204 158
rect 206 156 207 158
rect 203 155 207 156
rect 215 158 219 159
rect 215 156 216 158
rect 218 156 219 158
rect 215 155 219 156
rect 227 158 231 159
rect 227 156 228 158
rect 230 156 231 158
rect 227 155 231 156
rect 29 152 33 153
rect 29 150 30 152
rect 32 150 33 152
rect 29 149 33 150
rect 41 152 45 153
rect 41 150 42 152
rect 44 150 45 152
rect 41 149 45 150
rect 53 152 57 153
rect 53 150 54 152
rect 56 150 57 152
rect 53 149 57 150
rect 65 152 69 153
rect 65 150 66 152
rect 68 150 69 152
rect 65 149 69 150
rect 77 152 81 153
rect 77 150 78 152
rect 80 150 81 152
rect 77 149 81 150
rect 89 152 93 153
rect 89 150 90 152
rect 92 150 93 152
rect 89 149 93 150
rect 101 152 105 153
rect 101 150 102 152
rect 104 150 105 152
rect 101 149 105 150
rect 113 152 117 153
rect 113 150 114 152
rect 116 150 117 152
rect 113 149 117 150
rect 125 152 129 153
rect 125 150 126 152
rect 128 150 129 152
rect 125 149 129 150
rect 137 152 141 153
rect 137 150 138 152
rect 140 150 141 152
rect 137 149 141 150
rect 149 152 153 153
rect 149 150 150 152
rect 152 150 153 152
rect 149 149 153 150
rect 161 152 165 153
rect 161 150 162 152
rect 164 150 165 152
rect 161 149 165 150
rect 173 152 177 153
rect 173 150 174 152
rect 176 150 177 152
rect 173 149 177 150
rect 185 152 189 153
rect 185 150 186 152
rect 188 150 189 152
rect 185 149 189 150
rect 197 152 201 153
rect 197 150 198 152
rect 200 150 201 152
rect 197 149 201 150
rect 209 152 213 153
rect 209 150 210 152
rect 212 150 213 152
rect 209 149 213 150
rect 221 152 225 153
rect 221 150 222 152
rect 224 150 225 152
rect 221 149 225 150
rect 35 146 39 147
rect 35 144 36 146
rect 38 144 39 146
rect 35 143 39 144
rect 47 146 51 147
rect 47 144 48 146
rect 50 144 51 146
rect 47 143 51 144
rect 59 146 63 147
rect 59 144 60 146
rect 62 144 63 146
rect 59 143 63 144
rect 71 146 75 147
rect 71 144 72 146
rect 74 144 75 146
rect 71 143 75 144
rect 83 146 87 147
rect 83 144 84 146
rect 86 144 87 146
rect 83 143 87 144
rect 95 146 99 147
rect 95 144 96 146
rect 98 144 99 146
rect 95 143 99 144
rect 107 146 111 147
rect 107 144 108 146
rect 110 144 111 146
rect 107 143 111 144
rect 119 146 123 147
rect 119 144 120 146
rect 122 144 123 146
rect 119 143 123 144
rect 131 146 135 147
rect 131 144 132 146
rect 134 144 135 146
rect 131 143 135 144
rect 143 146 147 147
rect 143 144 144 146
rect 146 144 147 146
rect 143 143 147 144
rect 155 146 159 147
rect 155 144 156 146
rect 158 144 159 146
rect 155 143 159 144
rect 167 146 171 147
rect 167 144 168 146
rect 170 144 171 146
rect 167 143 171 144
rect 179 146 183 147
rect 179 144 180 146
rect 182 144 183 146
rect 179 143 183 144
rect 191 146 195 147
rect 191 144 192 146
rect 194 144 195 146
rect 191 143 195 144
rect 203 146 207 147
rect 203 144 204 146
rect 206 144 207 146
rect 203 143 207 144
rect 215 146 219 147
rect 215 144 216 146
rect 218 144 219 146
rect 215 143 219 144
rect 227 146 231 147
rect 227 144 228 146
rect 230 144 231 146
rect 227 143 231 144
rect 29 140 33 141
rect 29 138 30 140
rect 32 138 33 140
rect 29 137 33 138
rect 41 140 45 141
rect 41 138 42 140
rect 44 138 45 140
rect 41 137 45 138
rect 53 140 57 141
rect 53 138 54 140
rect 56 138 57 140
rect 53 137 57 138
rect 65 140 69 141
rect 65 138 66 140
rect 68 138 69 140
rect 65 137 69 138
rect 77 140 81 141
rect 77 138 78 140
rect 80 138 81 140
rect 77 137 81 138
rect 89 140 93 141
rect 89 138 90 140
rect 92 138 93 140
rect 89 137 93 138
rect 101 140 105 141
rect 101 138 102 140
rect 104 138 105 140
rect 101 137 105 138
rect 113 140 117 141
rect 113 138 114 140
rect 116 138 117 140
rect 113 137 117 138
rect 125 140 129 141
rect 125 138 126 140
rect 128 138 129 140
rect 125 137 129 138
rect 137 140 141 141
rect 137 138 138 140
rect 140 138 141 140
rect 137 137 141 138
rect 149 140 153 141
rect 149 138 150 140
rect 152 138 153 140
rect 149 137 153 138
rect 161 140 165 141
rect 161 138 162 140
rect 164 138 165 140
rect 161 137 165 138
rect 173 140 177 141
rect 173 138 174 140
rect 176 138 177 140
rect 173 137 177 138
rect 185 140 189 141
rect 185 138 186 140
rect 188 138 189 140
rect 185 137 189 138
rect 197 140 201 141
rect 197 138 198 140
rect 200 138 201 140
rect 197 137 201 138
rect 209 140 213 141
rect 209 138 210 140
rect 212 138 213 140
rect 209 137 213 138
rect 221 140 225 141
rect 221 138 222 140
rect 224 138 225 140
rect 221 137 225 138
rect 35 134 39 135
rect 35 132 36 134
rect 38 132 39 134
rect 35 131 39 132
rect 47 134 51 135
rect 47 132 48 134
rect 50 132 51 134
rect 47 131 51 132
rect 59 134 63 135
rect 59 132 60 134
rect 62 132 63 134
rect 59 131 63 132
rect 71 134 75 135
rect 71 132 72 134
rect 74 132 75 134
rect 71 131 75 132
rect 83 134 87 135
rect 83 132 84 134
rect 86 132 87 134
rect 83 131 87 132
rect 95 134 99 135
rect 95 132 96 134
rect 98 132 99 134
rect 95 131 99 132
rect 107 134 111 135
rect 107 132 108 134
rect 110 132 111 134
rect 107 131 111 132
rect 119 134 123 135
rect 119 132 120 134
rect 122 132 123 134
rect 119 131 123 132
rect 131 134 135 135
rect 131 132 132 134
rect 134 132 135 134
rect 131 131 135 132
rect 143 134 147 135
rect 143 132 144 134
rect 146 132 147 134
rect 143 131 147 132
rect 155 134 159 135
rect 155 132 156 134
rect 158 132 159 134
rect 155 131 159 132
rect 167 134 171 135
rect 167 132 168 134
rect 170 132 171 134
rect 167 131 171 132
rect 179 134 183 135
rect 179 132 180 134
rect 182 132 183 134
rect 179 131 183 132
rect 191 134 195 135
rect 191 132 192 134
rect 194 132 195 134
rect 191 131 195 132
rect 203 134 207 135
rect 203 132 204 134
rect 206 132 207 134
rect 203 131 207 132
rect 215 134 219 135
rect 215 132 216 134
rect 218 132 219 134
rect 215 131 219 132
rect 227 134 231 135
rect 227 132 228 134
rect 230 132 231 134
rect 227 131 231 132
rect 29 128 33 129
rect 29 126 30 128
rect 32 126 33 128
rect 29 125 33 126
rect 41 128 45 129
rect 41 126 42 128
rect 44 126 45 128
rect 41 125 45 126
rect 53 128 57 129
rect 53 126 54 128
rect 56 126 57 128
rect 53 125 57 126
rect 65 128 69 129
rect 65 126 66 128
rect 68 126 69 128
rect 65 125 69 126
rect 77 128 81 129
rect 77 126 78 128
rect 80 126 81 128
rect 77 125 81 126
rect 89 128 93 129
rect 89 126 90 128
rect 92 126 93 128
rect 89 125 93 126
rect 101 128 105 129
rect 101 126 102 128
rect 104 126 105 128
rect 101 125 105 126
rect 113 128 117 129
rect 113 126 114 128
rect 116 126 117 128
rect 113 125 117 126
rect 125 128 129 129
rect 125 126 126 128
rect 128 126 129 128
rect 125 125 129 126
rect 137 128 141 129
rect 137 126 138 128
rect 140 126 141 128
rect 137 125 141 126
rect 149 128 153 129
rect 149 126 150 128
rect 152 126 153 128
rect 149 125 153 126
rect 161 128 165 129
rect 161 126 162 128
rect 164 126 165 128
rect 161 125 165 126
rect 173 128 177 129
rect 173 126 174 128
rect 176 126 177 128
rect 173 125 177 126
rect 185 128 189 129
rect 185 126 186 128
rect 188 126 189 128
rect 185 125 189 126
rect 197 128 201 129
rect 197 126 198 128
rect 200 126 201 128
rect 197 125 201 126
rect 209 128 213 129
rect 209 126 210 128
rect 212 126 213 128
rect 209 125 213 126
rect 221 128 225 129
rect 221 126 222 128
rect 224 126 225 128
rect 221 125 225 126
rect 35 122 39 123
rect 35 120 36 122
rect 38 120 39 122
rect 35 119 39 120
rect 47 122 51 123
rect 47 120 48 122
rect 50 120 51 122
rect 47 119 51 120
rect 59 122 63 123
rect 59 120 60 122
rect 62 120 63 122
rect 59 119 63 120
rect 71 122 75 123
rect 71 120 72 122
rect 74 120 75 122
rect 71 119 75 120
rect 83 122 87 123
rect 83 120 84 122
rect 86 120 87 122
rect 83 119 87 120
rect 95 122 99 123
rect 95 120 96 122
rect 98 120 99 122
rect 95 119 99 120
rect 107 122 111 123
rect 107 120 108 122
rect 110 120 111 122
rect 107 119 111 120
rect 119 122 123 123
rect 119 120 120 122
rect 122 120 123 122
rect 119 119 123 120
rect 131 122 135 123
rect 131 120 132 122
rect 134 120 135 122
rect 131 119 135 120
rect 143 122 147 123
rect 143 120 144 122
rect 146 120 147 122
rect 143 119 147 120
rect 155 122 159 123
rect 155 120 156 122
rect 158 120 159 122
rect 155 119 159 120
rect 167 122 171 123
rect 167 120 168 122
rect 170 120 171 122
rect 167 119 171 120
rect 179 122 183 123
rect 179 120 180 122
rect 182 120 183 122
rect 179 119 183 120
rect 191 122 195 123
rect 191 120 192 122
rect 194 120 195 122
rect 191 119 195 120
rect 203 122 207 123
rect 203 120 204 122
rect 206 120 207 122
rect 203 119 207 120
rect 215 122 219 123
rect 215 120 216 122
rect 218 120 219 122
rect 215 119 219 120
rect 227 122 231 123
rect 227 120 228 122
rect 230 120 231 122
rect 227 119 231 120
rect 29 116 33 117
rect 29 114 30 116
rect 32 114 33 116
rect 29 113 33 114
rect 41 116 45 117
rect 41 114 42 116
rect 44 114 45 116
rect 41 113 45 114
rect 53 116 57 117
rect 53 114 54 116
rect 56 114 57 116
rect 53 113 57 114
rect 65 116 69 117
rect 65 114 66 116
rect 68 114 69 116
rect 65 113 69 114
rect 77 116 81 117
rect 77 114 78 116
rect 80 114 81 116
rect 77 113 81 114
rect 89 116 93 117
rect 89 114 90 116
rect 92 114 93 116
rect 89 113 93 114
rect 101 116 105 117
rect 101 114 102 116
rect 104 114 105 116
rect 101 113 105 114
rect 113 116 117 117
rect 113 114 114 116
rect 116 114 117 116
rect 113 113 117 114
rect 125 116 129 117
rect 125 114 126 116
rect 128 114 129 116
rect 125 113 129 114
rect 137 116 141 117
rect 137 114 138 116
rect 140 114 141 116
rect 137 113 141 114
rect 149 116 153 117
rect 149 114 150 116
rect 152 114 153 116
rect 149 113 153 114
rect 161 116 165 117
rect 161 114 162 116
rect 164 114 165 116
rect 161 113 165 114
rect 173 116 177 117
rect 173 114 174 116
rect 176 114 177 116
rect 173 113 177 114
rect 185 116 189 117
rect 185 114 186 116
rect 188 114 189 116
rect 185 113 189 114
rect 197 116 201 117
rect 197 114 198 116
rect 200 114 201 116
rect 197 113 201 114
rect 209 116 213 117
rect 209 114 210 116
rect 212 114 213 116
rect 209 113 213 114
rect 221 116 225 117
rect 221 114 222 116
rect 224 114 225 116
rect 221 113 225 114
rect 35 110 39 111
rect 35 108 36 110
rect 38 108 39 110
rect 35 107 39 108
rect 47 110 51 111
rect 47 108 48 110
rect 50 108 51 110
rect 47 107 51 108
rect 59 110 63 111
rect 59 108 60 110
rect 62 108 63 110
rect 59 107 63 108
rect 71 110 75 111
rect 71 108 72 110
rect 74 108 75 110
rect 71 107 75 108
rect 83 110 87 111
rect 83 108 84 110
rect 86 108 87 110
rect 83 107 87 108
rect 95 110 99 111
rect 95 108 96 110
rect 98 108 99 110
rect 95 107 99 108
rect 107 110 111 111
rect 107 108 108 110
rect 110 108 111 110
rect 107 107 111 108
rect 119 110 123 111
rect 119 108 120 110
rect 122 108 123 110
rect 119 107 123 108
rect 131 110 135 111
rect 131 108 132 110
rect 134 108 135 110
rect 131 107 135 108
rect 143 110 147 111
rect 143 108 144 110
rect 146 108 147 110
rect 143 107 147 108
rect 155 110 159 111
rect 155 108 156 110
rect 158 108 159 110
rect 155 107 159 108
rect 167 110 171 111
rect 167 108 168 110
rect 170 108 171 110
rect 167 107 171 108
rect 179 110 183 111
rect 179 108 180 110
rect 182 108 183 110
rect 179 107 183 108
rect 191 110 195 111
rect 191 108 192 110
rect 194 108 195 110
rect 191 107 195 108
rect 203 110 207 111
rect 203 108 204 110
rect 206 108 207 110
rect 203 107 207 108
rect 215 110 219 111
rect 215 108 216 110
rect 218 108 219 110
rect 215 107 219 108
rect 227 110 231 111
rect 227 108 228 110
rect 230 108 231 110
rect 227 107 231 108
rect 29 104 33 105
rect 29 102 30 104
rect 32 102 33 104
rect 29 101 33 102
rect 41 104 45 105
rect 41 102 42 104
rect 44 102 45 104
rect 41 101 45 102
rect 53 104 57 105
rect 53 102 54 104
rect 56 102 57 104
rect 53 101 57 102
rect 65 104 69 105
rect 65 102 66 104
rect 68 102 69 104
rect 65 101 69 102
rect 77 104 81 105
rect 77 102 78 104
rect 80 102 81 104
rect 77 101 81 102
rect 89 104 93 105
rect 89 102 90 104
rect 92 102 93 104
rect 89 101 93 102
rect 101 104 105 105
rect 101 102 102 104
rect 104 102 105 104
rect 101 101 105 102
rect 113 104 117 105
rect 113 102 114 104
rect 116 102 117 104
rect 113 101 117 102
rect 125 104 129 105
rect 125 102 126 104
rect 128 102 129 104
rect 125 101 129 102
rect 137 104 141 105
rect 137 102 138 104
rect 140 102 141 104
rect 137 101 141 102
rect 149 104 153 105
rect 149 102 150 104
rect 152 102 153 104
rect 149 101 153 102
rect 161 104 165 105
rect 161 102 162 104
rect 164 102 165 104
rect 161 101 165 102
rect 173 104 177 105
rect 173 102 174 104
rect 176 102 177 104
rect 173 101 177 102
rect 185 104 189 105
rect 185 102 186 104
rect 188 102 189 104
rect 185 101 189 102
rect 197 104 201 105
rect 197 102 198 104
rect 200 102 201 104
rect 197 101 201 102
rect 209 104 213 105
rect 209 102 210 104
rect 212 102 213 104
rect 209 101 213 102
rect 221 104 225 105
rect 221 102 222 104
rect 224 102 225 104
rect 221 101 225 102
rect 35 98 39 99
rect 35 96 36 98
rect 38 96 39 98
rect 35 95 39 96
rect 47 98 51 99
rect 47 96 48 98
rect 50 96 51 98
rect 47 95 51 96
rect 59 98 63 99
rect 59 96 60 98
rect 62 96 63 98
rect 59 95 63 96
rect 71 98 75 99
rect 71 96 72 98
rect 74 96 75 98
rect 71 95 75 96
rect 83 98 87 99
rect 83 96 84 98
rect 86 96 87 98
rect 83 95 87 96
rect 95 98 99 99
rect 95 96 96 98
rect 98 96 99 98
rect 95 95 99 96
rect 107 98 111 99
rect 107 96 108 98
rect 110 96 111 98
rect 107 95 111 96
rect 119 98 123 99
rect 119 96 120 98
rect 122 96 123 98
rect 119 95 123 96
rect 131 98 135 99
rect 131 96 132 98
rect 134 96 135 98
rect 131 95 135 96
rect 143 98 147 99
rect 143 96 144 98
rect 146 96 147 98
rect 143 95 147 96
rect 155 98 159 99
rect 155 96 156 98
rect 158 96 159 98
rect 155 95 159 96
rect 167 98 171 99
rect 167 96 168 98
rect 170 96 171 98
rect 167 95 171 96
rect 179 98 183 99
rect 179 96 180 98
rect 182 96 183 98
rect 179 95 183 96
rect 191 98 195 99
rect 191 96 192 98
rect 194 96 195 98
rect 191 95 195 96
rect 203 98 207 99
rect 203 96 204 98
rect 206 96 207 98
rect 203 95 207 96
rect 215 98 219 99
rect 215 96 216 98
rect 218 96 219 98
rect 215 95 219 96
rect 227 98 231 99
rect 227 96 228 98
rect 230 96 231 98
rect 227 95 231 96
rect 29 92 33 93
rect 29 90 30 92
rect 32 90 33 92
rect 29 89 33 90
rect 41 92 45 93
rect 41 90 42 92
rect 44 90 45 92
rect 41 89 45 90
rect 53 92 57 93
rect 53 90 54 92
rect 56 90 57 92
rect 53 89 57 90
rect 65 92 69 93
rect 65 90 66 92
rect 68 90 69 92
rect 65 89 69 90
rect 77 92 81 93
rect 77 90 78 92
rect 80 90 81 92
rect 77 89 81 90
rect 89 92 93 93
rect 89 90 90 92
rect 92 90 93 92
rect 89 89 93 90
rect 101 92 105 93
rect 101 90 102 92
rect 104 90 105 92
rect 101 89 105 90
rect 113 92 117 93
rect 113 90 114 92
rect 116 90 117 92
rect 113 89 117 90
rect 125 92 129 93
rect 125 90 126 92
rect 128 90 129 92
rect 125 89 129 90
rect 137 92 141 93
rect 137 90 138 92
rect 140 90 141 92
rect 137 89 141 90
rect 149 92 153 93
rect 149 90 150 92
rect 152 90 153 92
rect 149 89 153 90
rect 161 92 165 93
rect 161 90 162 92
rect 164 90 165 92
rect 161 89 165 90
rect 173 92 177 93
rect 173 90 174 92
rect 176 90 177 92
rect 173 89 177 90
rect 185 92 189 93
rect 185 90 186 92
rect 188 90 189 92
rect 185 89 189 90
rect 197 92 201 93
rect 197 90 198 92
rect 200 90 201 92
rect 197 89 201 90
rect 209 92 213 93
rect 209 90 210 92
rect 212 90 213 92
rect 209 89 213 90
rect 221 92 225 93
rect 221 90 222 92
rect 224 90 225 92
rect 221 89 225 90
rect 35 86 39 87
rect 35 84 36 86
rect 38 84 39 86
rect 35 83 39 84
rect 47 86 51 87
rect 47 84 48 86
rect 50 84 51 86
rect 47 83 51 84
rect 59 86 63 87
rect 59 84 60 86
rect 62 84 63 86
rect 59 83 63 84
rect 71 86 75 87
rect 71 84 72 86
rect 74 84 75 86
rect 71 83 75 84
rect 83 86 87 87
rect 83 84 84 86
rect 86 84 87 86
rect 83 83 87 84
rect 95 86 99 87
rect 95 84 96 86
rect 98 84 99 86
rect 95 83 99 84
rect 107 86 111 87
rect 107 84 108 86
rect 110 84 111 86
rect 107 83 111 84
rect 119 86 123 87
rect 119 84 120 86
rect 122 84 123 86
rect 119 83 123 84
rect 131 86 135 87
rect 131 84 132 86
rect 134 84 135 86
rect 131 83 135 84
rect 143 86 147 87
rect 143 84 144 86
rect 146 84 147 86
rect 143 83 147 84
rect 155 86 159 87
rect 155 84 156 86
rect 158 84 159 86
rect 155 83 159 84
rect 167 86 171 87
rect 167 84 168 86
rect 170 84 171 86
rect 167 83 171 84
rect 179 86 183 87
rect 179 84 180 86
rect 182 84 183 86
rect 179 83 183 84
rect 191 86 195 87
rect 191 84 192 86
rect 194 84 195 86
rect 191 83 195 84
rect 203 86 207 87
rect 203 84 204 86
rect 206 84 207 86
rect 203 83 207 84
rect 215 86 219 87
rect 215 84 216 86
rect 218 84 219 86
rect 215 83 219 84
rect 227 86 231 87
rect 227 84 228 86
rect 230 84 231 86
rect 227 83 231 84
rect 29 80 33 81
rect 29 78 30 80
rect 32 78 33 80
rect 29 77 33 78
rect 41 80 45 81
rect 41 78 42 80
rect 44 78 45 80
rect 41 77 45 78
rect 53 80 57 81
rect 53 78 54 80
rect 56 78 57 80
rect 53 77 57 78
rect 65 80 69 81
rect 65 78 66 80
rect 68 78 69 80
rect 65 77 69 78
rect 77 80 81 81
rect 77 78 78 80
rect 80 78 81 80
rect 77 77 81 78
rect 89 80 93 81
rect 89 78 90 80
rect 92 78 93 80
rect 89 77 93 78
rect 101 80 105 81
rect 101 78 102 80
rect 104 78 105 80
rect 101 77 105 78
rect 113 80 117 81
rect 113 78 114 80
rect 116 78 117 80
rect 113 77 117 78
rect 125 80 129 81
rect 125 78 126 80
rect 128 78 129 80
rect 125 77 129 78
rect 137 80 141 81
rect 137 78 138 80
rect 140 78 141 80
rect 137 77 141 78
rect 149 80 153 81
rect 149 78 150 80
rect 152 78 153 80
rect 149 77 153 78
rect 161 80 165 81
rect 161 78 162 80
rect 164 78 165 80
rect 161 77 165 78
rect 173 80 177 81
rect 173 78 174 80
rect 176 78 177 80
rect 173 77 177 78
rect 185 80 189 81
rect 185 78 186 80
rect 188 78 189 80
rect 185 77 189 78
rect 197 80 201 81
rect 197 78 198 80
rect 200 78 201 80
rect 197 77 201 78
rect 209 80 213 81
rect 209 78 210 80
rect 212 78 213 80
rect 209 77 213 78
rect 221 80 225 81
rect 221 78 222 80
rect 224 78 225 80
rect 221 77 225 78
rect 35 74 39 75
rect 35 72 36 74
rect 38 72 39 74
rect 35 71 39 72
rect 47 74 51 75
rect 47 72 48 74
rect 50 72 51 74
rect 47 71 51 72
rect 59 74 63 75
rect 59 72 60 74
rect 62 72 63 74
rect 59 71 63 72
rect 71 74 75 75
rect 71 72 72 74
rect 74 72 75 74
rect 71 71 75 72
rect 83 74 87 75
rect 83 72 84 74
rect 86 72 87 74
rect 83 71 87 72
rect 95 74 99 75
rect 95 72 96 74
rect 98 72 99 74
rect 95 71 99 72
rect 107 74 111 75
rect 107 72 108 74
rect 110 72 111 74
rect 107 71 111 72
rect 119 74 123 75
rect 119 72 120 74
rect 122 72 123 74
rect 119 71 123 72
rect 131 74 135 75
rect 131 72 132 74
rect 134 72 135 74
rect 131 71 135 72
rect 143 74 147 75
rect 143 72 144 74
rect 146 72 147 74
rect 143 71 147 72
rect 155 74 159 75
rect 155 72 156 74
rect 158 72 159 74
rect 155 71 159 72
rect 167 74 171 75
rect 167 72 168 74
rect 170 72 171 74
rect 167 71 171 72
rect 179 74 183 75
rect 179 72 180 74
rect 182 72 183 74
rect 179 71 183 72
rect 191 74 195 75
rect 191 72 192 74
rect 194 72 195 74
rect 191 71 195 72
rect 203 74 207 75
rect 203 72 204 74
rect 206 72 207 74
rect 203 71 207 72
rect 215 74 219 75
rect 215 72 216 74
rect 218 72 219 74
rect 215 71 219 72
rect 227 74 231 75
rect 227 72 228 74
rect 230 72 231 74
rect 227 71 231 72
rect 29 68 33 69
rect 29 66 30 68
rect 32 66 33 68
rect 29 65 33 66
rect 41 68 45 69
rect 41 66 42 68
rect 44 66 45 68
rect 41 65 45 66
rect 53 68 57 69
rect 53 66 54 68
rect 56 66 57 68
rect 53 65 57 66
rect 65 68 69 69
rect 65 66 66 68
rect 68 66 69 68
rect 65 65 69 66
rect 77 68 81 69
rect 77 66 78 68
rect 80 66 81 68
rect 77 65 81 66
rect 89 68 93 69
rect 89 66 90 68
rect 92 66 93 68
rect 89 65 93 66
rect 101 68 105 69
rect 101 66 102 68
rect 104 66 105 68
rect 101 65 105 66
rect 113 68 117 69
rect 113 66 114 68
rect 116 66 117 68
rect 113 65 117 66
rect 125 68 129 69
rect 125 66 126 68
rect 128 66 129 68
rect 125 65 129 66
rect 137 68 141 69
rect 137 66 138 68
rect 140 66 141 68
rect 137 65 141 66
rect 149 68 153 69
rect 149 66 150 68
rect 152 66 153 68
rect 149 65 153 66
rect 161 68 165 69
rect 161 66 162 68
rect 164 66 165 68
rect 161 65 165 66
rect 173 68 177 69
rect 173 66 174 68
rect 176 66 177 68
rect 173 65 177 66
rect 185 68 189 69
rect 185 66 186 68
rect 188 66 189 68
rect 185 65 189 66
rect 197 68 201 69
rect 197 66 198 68
rect 200 66 201 68
rect 197 65 201 66
rect 209 68 213 69
rect 209 66 210 68
rect 212 66 213 68
rect 209 65 213 66
rect 221 68 225 69
rect 221 66 222 68
rect 224 66 225 68
rect 221 65 225 66
rect 35 62 39 63
rect 35 60 36 62
rect 38 60 39 62
rect 35 59 39 60
rect 47 62 51 63
rect 47 60 48 62
rect 50 60 51 62
rect 47 59 51 60
rect 59 62 63 63
rect 59 60 60 62
rect 62 60 63 62
rect 59 59 63 60
rect 71 62 75 63
rect 71 60 72 62
rect 74 60 75 62
rect 71 59 75 60
rect 83 62 87 63
rect 83 60 84 62
rect 86 60 87 62
rect 83 59 87 60
rect 95 62 99 63
rect 95 60 96 62
rect 98 60 99 62
rect 95 59 99 60
rect 107 62 111 63
rect 107 60 108 62
rect 110 60 111 62
rect 107 59 111 60
rect 119 62 123 63
rect 119 60 120 62
rect 122 60 123 62
rect 119 59 123 60
rect 131 62 135 63
rect 131 60 132 62
rect 134 60 135 62
rect 131 59 135 60
rect 143 62 147 63
rect 143 60 144 62
rect 146 60 147 62
rect 143 59 147 60
rect 155 62 159 63
rect 155 60 156 62
rect 158 60 159 62
rect 155 59 159 60
rect 167 62 171 63
rect 167 60 168 62
rect 170 60 171 62
rect 167 59 171 60
rect 179 62 183 63
rect 179 60 180 62
rect 182 60 183 62
rect 179 59 183 60
rect 191 62 195 63
rect 191 60 192 62
rect 194 60 195 62
rect 191 59 195 60
rect 203 62 207 63
rect 203 60 204 62
rect 206 60 207 62
rect 203 59 207 60
rect 215 62 219 63
rect 215 60 216 62
rect 218 60 219 62
rect 215 59 219 60
rect 227 62 231 63
rect 227 60 228 62
rect 230 60 231 62
rect 227 59 231 60
rect 29 56 33 57
rect 29 54 30 56
rect 32 54 33 56
rect 29 53 33 54
rect 41 56 45 57
rect 41 54 42 56
rect 44 54 45 56
rect 41 53 45 54
rect 53 56 57 57
rect 53 54 54 56
rect 56 54 57 56
rect 53 53 57 54
rect 65 56 69 57
rect 65 54 66 56
rect 68 54 69 56
rect 65 53 69 54
rect 77 56 81 57
rect 77 54 78 56
rect 80 54 81 56
rect 77 53 81 54
rect 89 56 93 57
rect 89 54 90 56
rect 92 54 93 56
rect 89 53 93 54
rect 101 56 105 57
rect 101 54 102 56
rect 104 54 105 56
rect 101 53 105 54
rect 113 56 117 57
rect 113 54 114 56
rect 116 54 117 56
rect 113 53 117 54
rect 125 56 129 57
rect 125 54 126 56
rect 128 54 129 56
rect 125 53 129 54
rect 137 56 141 57
rect 137 54 138 56
rect 140 54 141 56
rect 137 53 141 54
rect 149 56 153 57
rect 149 54 150 56
rect 152 54 153 56
rect 149 53 153 54
rect 161 56 165 57
rect 161 54 162 56
rect 164 54 165 56
rect 161 53 165 54
rect 173 56 177 57
rect 173 54 174 56
rect 176 54 177 56
rect 173 53 177 54
rect 185 56 189 57
rect 185 54 186 56
rect 188 54 189 56
rect 185 53 189 54
rect 197 56 201 57
rect 197 54 198 56
rect 200 54 201 56
rect 197 53 201 54
rect 209 56 213 57
rect 209 54 210 56
rect 212 54 213 56
rect 209 53 213 54
rect 221 56 225 57
rect 221 54 222 56
rect 224 54 225 56
rect 221 53 225 54
rect 35 50 39 51
rect 35 48 36 50
rect 38 48 39 50
rect 35 47 39 48
rect 47 50 51 51
rect 47 48 48 50
rect 50 48 51 50
rect 47 47 51 48
rect 59 50 63 51
rect 59 48 60 50
rect 62 48 63 50
rect 59 47 63 48
rect 71 50 75 51
rect 71 48 72 50
rect 74 48 75 50
rect 71 47 75 48
rect 83 50 87 51
rect 83 48 84 50
rect 86 48 87 50
rect 83 47 87 48
rect 95 50 99 51
rect 95 48 96 50
rect 98 48 99 50
rect 95 47 99 48
rect 107 50 111 51
rect 107 48 108 50
rect 110 48 111 50
rect 107 47 111 48
rect 119 50 123 51
rect 119 48 120 50
rect 122 48 123 50
rect 119 47 123 48
rect 131 50 135 51
rect 131 48 132 50
rect 134 48 135 50
rect 131 47 135 48
rect 143 50 147 51
rect 143 48 144 50
rect 146 48 147 50
rect 143 47 147 48
rect 155 50 159 51
rect 155 48 156 50
rect 158 48 159 50
rect 155 47 159 48
rect 167 50 171 51
rect 167 48 168 50
rect 170 48 171 50
rect 167 47 171 48
rect 179 50 183 51
rect 179 48 180 50
rect 182 48 183 50
rect 179 47 183 48
rect 191 50 195 51
rect 191 48 192 50
rect 194 48 195 50
rect 191 47 195 48
rect 203 50 207 51
rect 203 48 204 50
rect 206 48 207 50
rect 203 47 207 48
rect 215 50 219 51
rect 215 48 216 50
rect 218 48 219 50
rect 215 47 219 48
rect 227 50 231 51
rect 227 48 228 50
rect 230 48 231 50
rect 227 47 231 48
rect 29 44 33 45
rect 29 42 30 44
rect 32 42 33 44
rect 29 41 33 42
rect 41 44 45 45
rect 41 42 42 44
rect 44 42 45 44
rect 41 41 45 42
rect 53 44 57 45
rect 53 42 54 44
rect 56 42 57 44
rect 53 41 57 42
rect 65 44 69 45
rect 65 42 66 44
rect 68 42 69 44
rect 65 41 69 42
rect 77 44 81 45
rect 77 42 78 44
rect 80 42 81 44
rect 77 41 81 42
rect 89 44 93 45
rect 89 42 90 44
rect 92 42 93 44
rect 89 41 93 42
rect 101 44 105 45
rect 101 42 102 44
rect 104 42 105 44
rect 101 41 105 42
rect 113 44 117 45
rect 113 42 114 44
rect 116 42 117 44
rect 113 41 117 42
rect 125 44 129 45
rect 125 42 126 44
rect 128 42 129 44
rect 125 41 129 42
rect 137 44 141 45
rect 137 42 138 44
rect 140 42 141 44
rect 137 41 141 42
rect 149 44 153 45
rect 149 42 150 44
rect 152 42 153 44
rect 149 41 153 42
rect 161 44 165 45
rect 161 42 162 44
rect 164 42 165 44
rect 161 41 165 42
rect 173 44 177 45
rect 173 42 174 44
rect 176 42 177 44
rect 173 41 177 42
rect 185 44 189 45
rect 185 42 186 44
rect 188 42 189 44
rect 185 41 189 42
rect 197 44 201 45
rect 197 42 198 44
rect 200 42 201 44
rect 197 41 201 42
rect 209 44 213 45
rect 209 42 210 44
rect 212 42 213 44
rect 209 41 213 42
rect 221 44 225 45
rect 221 42 222 44
rect 224 42 225 44
rect 221 41 225 42
rect 35 38 39 39
rect 35 36 36 38
rect 38 36 39 38
rect 35 35 39 36
rect 47 38 51 39
rect 47 36 48 38
rect 50 36 51 38
rect 47 35 51 36
rect 59 38 63 39
rect 59 36 60 38
rect 62 36 63 38
rect 59 35 63 36
rect 71 38 75 39
rect 71 36 72 38
rect 74 36 75 38
rect 71 35 75 36
rect 83 38 87 39
rect 83 36 84 38
rect 86 36 87 38
rect 83 35 87 36
rect 95 38 99 39
rect 95 36 96 38
rect 98 36 99 38
rect 95 35 99 36
rect 107 38 111 39
rect 107 36 108 38
rect 110 36 111 38
rect 107 35 111 36
rect 119 38 123 39
rect 119 36 120 38
rect 122 36 123 38
rect 119 35 123 36
rect 131 38 135 39
rect 131 36 132 38
rect 134 36 135 38
rect 131 35 135 36
rect 143 38 147 39
rect 143 36 144 38
rect 146 36 147 38
rect 143 35 147 36
rect 155 38 159 39
rect 155 36 156 38
rect 158 36 159 38
rect 155 35 159 36
rect 167 38 171 39
rect 167 36 168 38
rect 170 36 171 38
rect 167 35 171 36
rect 179 38 183 39
rect 179 36 180 38
rect 182 36 183 38
rect 179 35 183 36
rect 191 38 195 39
rect 191 36 192 38
rect 194 36 195 38
rect 191 35 195 36
rect 203 38 207 39
rect 203 36 204 38
rect 206 36 207 38
rect 203 35 207 36
rect 215 38 219 39
rect 215 36 216 38
rect 218 36 219 38
rect 215 35 219 36
rect 227 38 231 39
rect 227 36 228 38
rect 230 36 231 38
rect 227 35 231 36
rect 29 32 33 33
rect 29 30 30 32
rect 32 30 33 32
rect 29 29 33 30
rect 41 32 45 33
rect 41 30 42 32
rect 44 30 45 32
rect 41 29 45 30
rect 53 32 57 33
rect 53 30 54 32
rect 56 30 57 32
rect 53 29 57 30
rect 65 32 69 33
rect 65 30 66 32
rect 68 30 69 32
rect 65 29 69 30
rect 77 32 81 33
rect 77 30 78 32
rect 80 30 81 32
rect 77 29 81 30
rect 89 32 93 33
rect 89 30 90 32
rect 92 30 93 32
rect 89 29 93 30
rect 101 32 105 33
rect 101 30 102 32
rect 104 30 105 32
rect 101 29 105 30
rect 113 32 117 33
rect 113 30 114 32
rect 116 30 117 32
rect 113 29 117 30
rect 125 32 129 33
rect 125 30 126 32
rect 128 30 129 32
rect 125 29 129 30
rect 137 32 141 33
rect 137 30 138 32
rect 140 30 141 32
rect 137 29 141 30
rect 149 32 153 33
rect 149 30 150 32
rect 152 30 153 32
rect 149 29 153 30
rect 161 32 165 33
rect 161 30 162 32
rect 164 30 165 32
rect 161 29 165 30
rect 173 32 177 33
rect 173 30 174 32
rect 176 30 177 32
rect 173 29 177 30
rect 185 32 189 33
rect 185 30 186 32
rect 188 30 189 32
rect 185 29 189 30
rect 197 32 201 33
rect 197 30 198 32
rect 200 30 201 32
rect 197 29 201 30
rect 209 32 213 33
rect 209 30 210 32
rect 212 30 213 32
rect 209 29 213 30
rect 221 32 225 33
rect 221 30 222 32
rect 224 30 225 32
rect 221 29 225 30
<< nwell >>
rect 0 0 260 260
<< metal1 >>
rect 0 257 260 260
rect 0 3 3 257
rect 257 3 260 257
rect 0 0 260 3
<< metal2 >>
rect 0 257 260 260
rect 0 3 3 257
rect 257 3 260 257
rect 0 0 260 3
<< pad >>
rect 3 3 257 257
use PadBoxX  PadBoxX_0
timestamp 1570494029
transform 1 0 30 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_1
timestamp 1570494029
transform 1 0 42 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_2
timestamp 1570494029
transform 1 0 54 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_3
timestamp 1570494029
transform 1 0 66 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_4
timestamp 1570494029
transform 1 0 78 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_5
timestamp 1570494029
transform 1 0 90 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_6
timestamp 1570494029
transform 1 0 102 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_7
timestamp 1570494029
transform 1 0 114 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_8
timestamp 1570494029
transform 1 0 126 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_9
timestamp 1570494029
transform 1 0 138 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_10
timestamp 1570494029
transform 1 0 150 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_11
timestamp 1570494029
transform 1 0 162 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_12
timestamp 1570494029
transform 1 0 174 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_13
timestamp 1570494029
transform 1 0 186 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_14
timestamp 1570494029
transform 1 0 198 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_15
timestamp 1570494029
transform 1 0 210 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_16
timestamp 1570494029
transform 1 0 222 0 1 222
box -1 -1 10 10
use PadBoxX  PadBoxX_17
timestamp 1570494029
transform 1 0 30 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_18
timestamp 1570494029
transform 1 0 42 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_19
timestamp 1570494029
transform 1 0 54 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_20
timestamp 1570494029
transform 1 0 66 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_21
timestamp 1570494029
transform 1 0 78 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_22
timestamp 1570494029
transform 1 0 90 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_23
timestamp 1570494029
transform 1 0 102 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_24
timestamp 1570494029
transform 1 0 114 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_25
timestamp 1570494029
transform 1 0 126 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_26
timestamp 1570494029
transform 1 0 138 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_27
timestamp 1570494029
transform 1 0 150 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_28
timestamp 1570494029
transform 1 0 162 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_29
timestamp 1570494029
transform 1 0 174 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_30
timestamp 1570494029
transform 1 0 186 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_31
timestamp 1570494029
transform 1 0 198 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_32
timestamp 1570494029
transform 1 0 210 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_33
timestamp 1570494029
transform 1 0 222 0 1 210
box -1 -1 10 10
use PadBoxX  PadBoxX_34
timestamp 1570494029
transform 1 0 30 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_35
timestamp 1570494029
transform 1 0 42 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_36
timestamp 1570494029
transform 1 0 54 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_37
timestamp 1570494029
transform 1 0 66 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_38
timestamp 1570494029
transform 1 0 78 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_39
timestamp 1570494029
transform 1 0 90 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_40
timestamp 1570494029
transform 1 0 102 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_41
timestamp 1570494029
transform 1 0 114 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_42
timestamp 1570494029
transform 1 0 126 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_43
timestamp 1570494029
transform 1 0 138 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_44
timestamp 1570494029
transform 1 0 150 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_45
timestamp 1570494029
transform 1 0 162 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_46
timestamp 1570494029
transform 1 0 174 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_47
timestamp 1570494029
transform 1 0 186 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_48
timestamp 1570494029
transform 1 0 198 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_49
timestamp 1570494029
transform 1 0 210 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_50
timestamp 1570494029
transform 1 0 222 0 1 198
box -1 -1 10 10
use PadBoxX  PadBoxX_51
timestamp 1570494029
transform 1 0 30 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_52
timestamp 1570494029
transform 1 0 42 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_53
timestamp 1570494029
transform 1 0 54 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_54
timestamp 1570494029
transform 1 0 66 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_55
timestamp 1570494029
transform 1 0 78 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_56
timestamp 1570494029
transform 1 0 90 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_57
timestamp 1570494029
transform 1 0 102 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_58
timestamp 1570494029
transform 1 0 114 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_59
timestamp 1570494029
transform 1 0 126 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_60
timestamp 1570494029
transform 1 0 138 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_61
timestamp 1570494029
transform 1 0 150 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_62
timestamp 1570494029
transform 1 0 162 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_63
timestamp 1570494029
transform 1 0 174 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_64
timestamp 1570494029
transform 1 0 186 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_65
timestamp 1570494029
transform 1 0 198 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_66
timestamp 1570494029
transform 1 0 210 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_67
timestamp 1570494029
transform 1 0 222 0 1 186
box -1 -1 10 10
use PadBoxX  PadBoxX_68
timestamp 1570494029
transform 1 0 30 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_69
timestamp 1570494029
transform 1 0 42 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_70
timestamp 1570494029
transform 1 0 54 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_71
timestamp 1570494029
transform 1 0 66 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_72
timestamp 1570494029
transform 1 0 78 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_73
timestamp 1570494029
transform 1 0 90 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_74
timestamp 1570494029
transform 1 0 102 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_75
timestamp 1570494029
transform 1 0 114 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_76
timestamp 1570494029
transform 1 0 126 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_77
timestamp 1570494029
transform 1 0 138 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_78
timestamp 1570494029
transform 1 0 150 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_79
timestamp 1570494029
transform 1 0 162 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_80
timestamp 1570494029
transform 1 0 174 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_81
timestamp 1570494029
transform 1 0 186 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_82
timestamp 1570494029
transform 1 0 198 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_83
timestamp 1570494029
transform 1 0 210 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_84
timestamp 1570494029
transform 1 0 222 0 1 174
box -1 -1 10 10
use PadBoxX  PadBoxX_85
timestamp 1570494029
transform 1 0 30 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_86
timestamp 1570494029
transform 1 0 42 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_87
timestamp 1570494029
transform 1 0 54 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_88
timestamp 1570494029
transform 1 0 66 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_89
timestamp 1570494029
transform 1 0 78 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_90
timestamp 1570494029
transform 1 0 90 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_91
timestamp 1570494029
transform 1 0 102 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_92
timestamp 1570494029
transform 1 0 114 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_93
timestamp 1570494029
transform 1 0 126 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_94
timestamp 1570494029
transform 1 0 138 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_95
timestamp 1570494029
transform 1 0 150 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_96
timestamp 1570494029
transform 1 0 162 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_97
timestamp 1570494029
transform 1 0 174 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_98
timestamp 1570494029
transform 1 0 186 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_99
timestamp 1570494029
transform 1 0 198 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_100
timestamp 1570494029
transform 1 0 210 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_101
timestamp 1570494029
transform 1 0 222 0 1 162
box -1 -1 10 10
use PadBoxX  PadBoxX_102
timestamp 1570494029
transform 1 0 30 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_103
timestamp 1570494029
transform 1 0 42 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_104
timestamp 1570494029
transform 1 0 54 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_105
timestamp 1570494029
transform 1 0 66 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_106
timestamp 1570494029
transform 1 0 78 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_107
timestamp 1570494029
transform 1 0 90 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_108
timestamp 1570494029
transform 1 0 102 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_109
timestamp 1570494029
transform 1 0 114 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_110
timestamp 1570494029
transform 1 0 126 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_111
timestamp 1570494029
transform 1 0 138 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_112
timestamp 1570494029
transform 1 0 150 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_113
timestamp 1570494029
transform 1 0 162 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_114
timestamp 1570494029
transform 1 0 174 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_115
timestamp 1570494029
transform 1 0 186 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_116
timestamp 1570494029
transform 1 0 198 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_117
timestamp 1570494029
transform 1 0 210 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_118
timestamp 1570494029
transform 1 0 222 0 1 150
box -1 -1 10 10
use PadBoxX  PadBoxX_119
timestamp 1570494029
transform 1 0 30 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_120
timestamp 1570494029
transform 1 0 42 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_121
timestamp 1570494029
transform 1 0 54 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_122
timestamp 1570494029
transform 1 0 66 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_123
timestamp 1570494029
transform 1 0 78 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_124
timestamp 1570494029
transform 1 0 90 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_125
timestamp 1570494029
transform 1 0 102 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_126
timestamp 1570494029
transform 1 0 114 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_127
timestamp 1570494029
transform 1 0 126 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_128
timestamp 1570494029
transform 1 0 138 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_129
timestamp 1570494029
transform 1 0 150 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_130
timestamp 1570494029
transform 1 0 162 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_131
timestamp 1570494029
transform 1 0 174 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_132
timestamp 1570494029
transform 1 0 186 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_133
timestamp 1570494029
transform 1 0 198 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_134
timestamp 1570494029
transform 1 0 210 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_135
timestamp 1570494029
transform 1 0 222 0 1 138
box -1 -1 10 10
use PadBoxX  PadBoxX_136
timestamp 1570494029
transform 1 0 30 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_137
timestamp 1570494029
transform 1 0 42 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_138
timestamp 1570494029
transform 1 0 54 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_139
timestamp 1570494029
transform 1 0 66 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_140
timestamp 1570494029
transform 1 0 78 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_141
timestamp 1570494029
transform 1 0 90 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_142
timestamp 1570494029
transform 1 0 102 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_143
timestamp 1570494029
transform 1 0 114 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_144
timestamp 1570494029
transform 1 0 126 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_145
timestamp 1570494029
transform 1 0 138 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_146
timestamp 1570494029
transform 1 0 150 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_147
timestamp 1570494029
transform 1 0 162 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_148
timestamp 1570494029
transform 1 0 174 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_149
timestamp 1570494029
transform 1 0 186 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_150
timestamp 1570494029
transform 1 0 198 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_151
timestamp 1570494029
transform 1 0 210 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_152
timestamp 1570494029
transform 1 0 222 0 1 126
box -1 -1 10 10
use PadBoxX  PadBoxX_153
timestamp 1570494029
transform 1 0 30 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_154
timestamp 1570494029
transform 1 0 42 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_155
timestamp 1570494029
transform 1 0 54 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_156
timestamp 1570494029
transform 1 0 66 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_157
timestamp 1570494029
transform 1 0 78 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_158
timestamp 1570494029
transform 1 0 90 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_159
timestamp 1570494029
transform 1 0 102 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_160
timestamp 1570494029
transform 1 0 114 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_161
timestamp 1570494029
transform 1 0 126 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_162
timestamp 1570494029
transform 1 0 138 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_163
timestamp 1570494029
transform 1 0 150 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_164
timestamp 1570494029
transform 1 0 162 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_165
timestamp 1570494029
transform 1 0 174 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_166
timestamp 1570494029
transform 1 0 186 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_167
timestamp 1570494029
transform 1 0 198 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_168
timestamp 1570494029
transform 1 0 210 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_169
timestamp 1570494029
transform 1 0 222 0 1 114
box -1 -1 10 10
use PadBoxX  PadBoxX_170
timestamp 1570494029
transform 1 0 30 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_171
timestamp 1570494029
transform 1 0 42 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_172
timestamp 1570494029
transform 1 0 54 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_173
timestamp 1570494029
transform 1 0 66 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_174
timestamp 1570494029
transform 1 0 78 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_175
timestamp 1570494029
transform 1 0 90 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_176
timestamp 1570494029
transform 1 0 102 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_177
timestamp 1570494029
transform 1 0 114 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_178
timestamp 1570494029
transform 1 0 126 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_179
timestamp 1570494029
transform 1 0 138 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_180
timestamp 1570494029
transform 1 0 150 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_181
timestamp 1570494029
transform 1 0 162 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_182
timestamp 1570494029
transform 1 0 174 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_183
timestamp 1570494029
transform 1 0 186 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_184
timestamp 1570494029
transform 1 0 198 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_185
timestamp 1570494029
transform 1 0 210 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_186
timestamp 1570494029
transform 1 0 222 0 1 102
box -1 -1 10 10
use PadBoxX  PadBoxX_187
timestamp 1570494029
transform 1 0 30 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_188
timestamp 1570494029
transform 1 0 42 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_189
timestamp 1570494029
transform 1 0 54 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_190
timestamp 1570494029
transform 1 0 66 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_191
timestamp 1570494029
transform 1 0 78 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_192
timestamp 1570494029
transform 1 0 90 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_193
timestamp 1570494029
transform 1 0 102 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_194
timestamp 1570494029
transform 1 0 114 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_195
timestamp 1570494029
transform 1 0 126 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_196
timestamp 1570494029
transform 1 0 138 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_197
timestamp 1570494029
transform 1 0 150 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_198
timestamp 1570494029
transform 1 0 162 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_199
timestamp 1570494029
transform 1 0 174 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_200
timestamp 1570494029
transform 1 0 186 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_201
timestamp 1570494029
transform 1 0 198 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_202
timestamp 1570494029
transform 1 0 210 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_203
timestamp 1570494029
transform 1 0 222 0 1 90
box -1 -1 10 10
use PadBoxX  PadBoxX_204
timestamp 1570494029
transform 1 0 30 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_205
timestamp 1570494029
transform 1 0 42 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_206
timestamp 1570494029
transform 1 0 54 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_207
timestamp 1570494029
transform 1 0 66 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_208
timestamp 1570494029
transform 1 0 78 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_209
timestamp 1570494029
transform 1 0 90 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_210
timestamp 1570494029
transform 1 0 102 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_211
timestamp 1570494029
transform 1 0 114 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_212
timestamp 1570494029
transform 1 0 126 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_213
timestamp 1570494029
transform 1 0 138 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_214
timestamp 1570494029
transform 1 0 150 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_215
timestamp 1570494029
transform 1 0 162 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_216
timestamp 1570494029
transform 1 0 174 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_217
timestamp 1570494029
transform 1 0 186 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_218
timestamp 1570494029
transform 1 0 198 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_219
timestamp 1570494029
transform 1 0 210 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_220
timestamp 1570494029
transform 1 0 222 0 1 78
box -1 -1 10 10
use PadBoxX  PadBoxX_221
timestamp 1570494029
transform 1 0 30 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_222
timestamp 1570494029
transform 1 0 42 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_223
timestamp 1570494029
transform 1 0 54 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_224
timestamp 1570494029
transform 1 0 66 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_225
timestamp 1570494029
transform 1 0 78 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_226
timestamp 1570494029
transform 1 0 90 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_227
timestamp 1570494029
transform 1 0 102 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_228
timestamp 1570494029
transform 1 0 114 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_229
timestamp 1570494029
transform 1 0 126 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_230
timestamp 1570494029
transform 1 0 138 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_231
timestamp 1570494029
transform 1 0 150 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_232
timestamp 1570494029
transform 1 0 162 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_233
timestamp 1570494029
transform 1 0 174 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_234
timestamp 1570494029
transform 1 0 186 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_235
timestamp 1570494029
transform 1 0 198 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_236
timestamp 1570494029
transform 1 0 210 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_237
timestamp 1570494029
transform 1 0 222 0 1 66
box -1 -1 10 10
use PadBoxX  PadBoxX_238
timestamp 1570494029
transform 1 0 30 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_239
timestamp 1570494029
transform 1 0 42 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_240
timestamp 1570494029
transform 1 0 54 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_241
timestamp 1570494029
transform 1 0 66 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_242
timestamp 1570494029
transform 1 0 78 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_243
timestamp 1570494029
transform 1 0 90 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_244
timestamp 1570494029
transform 1 0 102 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_245
timestamp 1570494029
transform 1 0 114 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_246
timestamp 1570494029
transform 1 0 126 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_247
timestamp 1570494029
transform 1 0 138 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_248
timestamp 1570494029
transform 1 0 150 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_249
timestamp 1570494029
transform 1 0 162 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_250
timestamp 1570494029
transform 1 0 174 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_251
timestamp 1570494029
transform 1 0 186 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_252
timestamp 1570494029
transform 1 0 198 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_253
timestamp 1570494029
transform 1 0 210 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_254
timestamp 1570494029
transform 1 0 222 0 1 54
box -1 -1 10 10
use PadBoxX  PadBoxX_255
timestamp 1570494029
transform 1 0 30 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_256
timestamp 1570494029
transform 1 0 42 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_257
timestamp 1570494029
transform 1 0 54 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_258
timestamp 1570494029
transform 1 0 66 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_259
timestamp 1570494029
transform 1 0 78 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_260
timestamp 1570494029
transform 1 0 90 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_261
timestamp 1570494029
transform 1 0 102 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_262
timestamp 1570494029
transform 1 0 114 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_263
timestamp 1570494029
transform 1 0 126 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_264
timestamp 1570494029
transform 1 0 138 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_265
timestamp 1570494029
transform 1 0 150 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_266
timestamp 1570494029
transform 1 0 162 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_267
timestamp 1570494029
transform 1 0 174 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_268
timestamp 1570494029
transform 1 0 186 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_269
timestamp 1570494029
transform 1 0 198 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_270
timestamp 1570494029
transform 1 0 210 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_271
timestamp 1570494029
transform 1 0 222 0 1 42
box -1 -1 10 10
use PadBoxX  PadBoxX_272
timestamp 1570494029
transform 1 0 30 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_273
timestamp 1570494029
transform 1 0 42 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_274
timestamp 1570494029
transform 1 0 54 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_275
timestamp 1570494029
transform 1 0 66 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_276
timestamp 1570494029
transform 1 0 78 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_277
timestamp 1570494029
transform 1 0 90 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_278
timestamp 1570494029
transform 1 0 102 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_279
timestamp 1570494029
transform 1 0 114 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_280
timestamp 1570494029
transform 1 0 126 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_281
timestamp 1570494029
transform 1 0 138 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_282
timestamp 1570494029
transform 1 0 150 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_283
timestamp 1570494029
transform 1 0 162 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_284
timestamp 1570494029
transform 1 0 174 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_285
timestamp 1570494029
transform 1 0 186 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_286
timestamp 1570494029
transform 1 0 198 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_287
timestamp 1570494029
transform 1 0 210 0 1 30
box -1 -1 10 10
use PadBoxX  PadBoxX_288
timestamp 1570494029
transform 1 0 222 0 1 30
box -1 -1 10 10
<< properties >>
string path 0.000 0.000 1170.000 0.000 1170.000 1170.000 0.000 1170.000 0.000 0.000 
<< end >>
