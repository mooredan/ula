`celldefine
module decap8 ();
endmodule
`endcelldefine
