`celldefine
module buf_c (z, a);
  output z;
  input  a;

  buf G1 (z, a);
endmodule
`endcelldefine
