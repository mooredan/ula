magic
tech scmos
magscale 1 2
timestamp 1570494029
<< error_p >>
rect 12 1328 14 1330
rect 586 1328 588 1330
rect 10 1326 12 1328
rect 588 1326 590 1328
rect 74 1290 76 1292
rect 104 1290 106 1292
rect 134 1290 136 1292
rect 164 1290 166 1292
rect 194 1290 196 1292
rect 224 1290 226 1292
rect 254 1290 256 1292
rect 284 1290 286 1292
rect 314 1290 316 1292
rect 344 1290 346 1292
rect 374 1290 376 1292
rect 404 1290 406 1292
rect 434 1290 436 1292
rect 464 1290 466 1292
rect 494 1290 496 1292
rect 524 1290 526 1292
rect 76 1288 78 1290
rect 82 1288 84 1290
rect 106 1288 108 1290
rect 112 1288 114 1290
rect 136 1288 138 1290
rect 142 1288 144 1290
rect 166 1288 168 1290
rect 172 1288 174 1290
rect 196 1288 198 1290
rect 202 1288 204 1290
rect 226 1288 228 1290
rect 232 1288 234 1290
rect 256 1288 258 1290
rect 262 1288 264 1290
rect 286 1288 288 1290
rect 292 1288 294 1290
rect 316 1288 318 1290
rect 322 1288 324 1290
rect 346 1288 348 1290
rect 352 1288 354 1290
rect 376 1288 378 1290
rect 382 1288 384 1290
rect 406 1288 408 1290
rect 412 1288 414 1290
rect 436 1288 438 1290
rect 442 1288 444 1290
rect 466 1288 468 1290
rect 472 1288 474 1290
rect 496 1288 498 1290
rect 502 1288 504 1290
rect 526 1288 528 1290
rect 532 1288 534 1290
rect 84 1286 86 1288
rect 114 1286 116 1288
rect 144 1286 146 1288
rect 174 1286 176 1288
rect 204 1286 206 1288
rect 234 1286 236 1288
rect 264 1286 266 1288
rect 294 1286 296 1288
rect 324 1286 326 1288
rect 354 1286 356 1288
rect 384 1286 386 1288
rect 414 1286 416 1288
rect 444 1286 446 1288
rect 474 1286 476 1288
rect 504 1286 506 1288
rect 534 1286 536 1288
rect 84 1280 86 1282
rect 114 1280 116 1282
rect 144 1280 146 1282
rect 174 1280 176 1282
rect 204 1280 206 1282
rect 234 1280 236 1282
rect 264 1280 266 1282
rect 294 1280 296 1282
rect 324 1280 326 1282
rect 354 1280 356 1282
rect 384 1280 386 1282
rect 414 1280 416 1282
rect 444 1280 446 1282
rect 474 1280 476 1282
rect 504 1280 506 1282
rect 534 1280 536 1282
rect 76 1278 78 1280
rect 82 1278 84 1280
rect 106 1278 108 1280
rect 112 1278 114 1280
rect 136 1278 138 1280
rect 142 1278 144 1280
rect 166 1278 168 1280
rect 172 1278 174 1280
rect 196 1278 198 1280
rect 202 1278 204 1280
rect 226 1278 228 1280
rect 232 1278 234 1280
rect 256 1278 258 1280
rect 262 1278 264 1280
rect 286 1278 288 1280
rect 292 1278 294 1280
rect 316 1278 318 1280
rect 322 1278 324 1280
rect 346 1278 348 1280
rect 352 1278 354 1280
rect 376 1278 378 1280
rect 382 1278 384 1280
rect 406 1278 408 1280
rect 412 1278 414 1280
rect 436 1278 438 1280
rect 442 1278 444 1280
rect 466 1278 468 1280
rect 472 1278 474 1280
rect 496 1278 498 1280
rect 502 1278 504 1280
rect 526 1278 528 1280
rect 532 1278 534 1280
rect 74 1276 76 1278
rect 104 1276 106 1278
rect 134 1276 136 1278
rect 164 1276 166 1278
rect 194 1276 196 1278
rect 224 1276 226 1278
rect 254 1276 256 1278
rect 284 1276 286 1278
rect 314 1276 316 1278
rect 344 1276 346 1278
rect 374 1276 376 1278
rect 404 1276 406 1278
rect 434 1276 436 1278
rect 464 1276 466 1278
rect 494 1276 496 1278
rect 524 1276 526 1278
rect 74 1270 76 1272
rect 104 1270 106 1272
rect 134 1270 136 1272
rect 164 1270 166 1272
rect 194 1270 196 1272
rect 224 1270 226 1272
rect 254 1270 256 1272
rect 284 1270 286 1272
rect 314 1270 316 1272
rect 344 1270 346 1272
rect 374 1270 376 1272
rect 404 1270 406 1272
rect 434 1270 436 1272
rect 464 1270 466 1272
rect 494 1270 496 1272
rect 524 1270 526 1272
rect 76 1268 78 1270
rect 82 1268 84 1270
rect 106 1268 108 1270
rect 112 1268 114 1270
rect 136 1268 138 1270
rect 142 1268 144 1270
rect 166 1268 168 1270
rect 172 1268 174 1270
rect 196 1268 198 1270
rect 202 1268 204 1270
rect 226 1268 228 1270
rect 232 1268 234 1270
rect 256 1268 258 1270
rect 262 1268 264 1270
rect 286 1268 288 1270
rect 292 1268 294 1270
rect 316 1268 318 1270
rect 322 1268 324 1270
rect 346 1268 348 1270
rect 352 1268 354 1270
rect 376 1268 378 1270
rect 382 1268 384 1270
rect 406 1268 408 1270
rect 412 1268 414 1270
rect 436 1268 438 1270
rect 442 1268 444 1270
rect 466 1268 468 1270
rect 472 1268 474 1270
rect 496 1268 498 1270
rect 502 1268 504 1270
rect 526 1268 528 1270
rect 532 1268 534 1270
rect 84 1266 86 1268
rect 114 1266 116 1268
rect 144 1266 146 1268
rect 174 1266 176 1268
rect 204 1266 206 1268
rect 234 1266 236 1268
rect 264 1266 266 1268
rect 294 1266 296 1268
rect 324 1266 326 1268
rect 354 1266 356 1268
rect 384 1266 386 1268
rect 414 1266 416 1268
rect 444 1266 446 1268
rect 474 1266 476 1268
rect 504 1266 506 1268
rect 534 1266 536 1268
rect 84 1260 86 1262
rect 114 1260 116 1262
rect 144 1260 146 1262
rect 174 1260 176 1262
rect 204 1260 206 1262
rect 234 1260 236 1262
rect 264 1260 266 1262
rect 294 1260 296 1262
rect 324 1260 326 1262
rect 354 1260 356 1262
rect 384 1260 386 1262
rect 414 1260 416 1262
rect 444 1260 446 1262
rect 474 1260 476 1262
rect 504 1260 506 1262
rect 534 1260 536 1262
rect 76 1258 78 1260
rect 82 1258 84 1260
rect 106 1258 108 1260
rect 112 1258 114 1260
rect 136 1258 138 1260
rect 142 1258 144 1260
rect 166 1258 168 1260
rect 172 1258 174 1260
rect 196 1258 198 1260
rect 202 1258 204 1260
rect 226 1258 228 1260
rect 232 1258 234 1260
rect 256 1258 258 1260
rect 262 1258 264 1260
rect 286 1258 288 1260
rect 292 1258 294 1260
rect 316 1258 318 1260
rect 322 1258 324 1260
rect 346 1258 348 1260
rect 352 1258 354 1260
rect 376 1258 378 1260
rect 382 1258 384 1260
rect 406 1258 408 1260
rect 412 1258 414 1260
rect 436 1258 438 1260
rect 442 1258 444 1260
rect 466 1258 468 1260
rect 472 1258 474 1260
rect 496 1258 498 1260
rect 502 1258 504 1260
rect 526 1258 528 1260
rect 532 1258 534 1260
rect 74 1256 76 1258
rect 104 1256 106 1258
rect 134 1256 136 1258
rect 164 1256 166 1258
rect 194 1256 196 1258
rect 224 1256 226 1258
rect 254 1256 256 1258
rect 284 1256 286 1258
rect 314 1256 316 1258
rect 344 1256 346 1258
rect 374 1256 376 1258
rect 404 1256 406 1258
rect 434 1256 436 1258
rect 464 1256 466 1258
rect 494 1256 496 1258
rect 524 1256 526 1258
rect 74 1250 76 1252
rect 104 1250 106 1252
rect 134 1250 136 1252
rect 164 1250 166 1252
rect 194 1250 196 1252
rect 224 1250 226 1252
rect 254 1250 256 1252
rect 284 1250 286 1252
rect 314 1250 316 1252
rect 344 1250 346 1252
rect 374 1250 376 1252
rect 404 1250 406 1252
rect 434 1250 436 1252
rect 464 1250 466 1252
rect 494 1250 496 1252
rect 524 1250 526 1252
rect 76 1248 78 1250
rect 82 1248 84 1250
rect 106 1248 108 1250
rect 112 1248 114 1250
rect 136 1248 138 1250
rect 142 1248 144 1250
rect 166 1248 168 1250
rect 172 1248 174 1250
rect 196 1248 198 1250
rect 202 1248 204 1250
rect 226 1248 228 1250
rect 232 1248 234 1250
rect 256 1248 258 1250
rect 262 1248 264 1250
rect 286 1248 288 1250
rect 292 1248 294 1250
rect 316 1248 318 1250
rect 322 1248 324 1250
rect 346 1248 348 1250
rect 352 1248 354 1250
rect 376 1248 378 1250
rect 382 1248 384 1250
rect 406 1248 408 1250
rect 412 1248 414 1250
rect 436 1248 438 1250
rect 442 1248 444 1250
rect 466 1248 468 1250
rect 472 1248 474 1250
rect 496 1248 498 1250
rect 502 1248 504 1250
rect 526 1248 528 1250
rect 532 1248 534 1250
rect 84 1246 86 1248
rect 114 1246 116 1248
rect 144 1246 146 1248
rect 174 1246 176 1248
rect 204 1246 206 1248
rect 234 1246 236 1248
rect 264 1246 266 1248
rect 294 1246 296 1248
rect 324 1246 326 1248
rect 354 1246 356 1248
rect 384 1246 386 1248
rect 414 1246 416 1248
rect 444 1246 446 1248
rect 474 1246 476 1248
rect 504 1246 506 1248
rect 534 1246 536 1248
rect 84 1240 86 1242
rect 114 1240 116 1242
rect 144 1240 146 1242
rect 174 1240 176 1242
rect 204 1240 206 1242
rect 234 1240 236 1242
rect 264 1240 266 1242
rect 294 1240 296 1242
rect 324 1240 326 1242
rect 354 1240 356 1242
rect 384 1240 386 1242
rect 414 1240 416 1242
rect 444 1240 446 1242
rect 474 1240 476 1242
rect 504 1240 506 1242
rect 534 1240 536 1242
rect 76 1238 78 1240
rect 82 1238 84 1240
rect 106 1238 108 1240
rect 112 1238 114 1240
rect 136 1238 138 1240
rect 142 1238 144 1240
rect 166 1238 168 1240
rect 172 1238 174 1240
rect 196 1238 198 1240
rect 202 1238 204 1240
rect 226 1238 228 1240
rect 232 1238 234 1240
rect 256 1238 258 1240
rect 262 1238 264 1240
rect 286 1238 288 1240
rect 292 1238 294 1240
rect 316 1238 318 1240
rect 322 1238 324 1240
rect 346 1238 348 1240
rect 352 1238 354 1240
rect 376 1238 378 1240
rect 382 1238 384 1240
rect 406 1238 408 1240
rect 412 1238 414 1240
rect 436 1238 438 1240
rect 442 1238 444 1240
rect 466 1238 468 1240
rect 472 1238 474 1240
rect 496 1238 498 1240
rect 502 1238 504 1240
rect 526 1238 528 1240
rect 532 1238 534 1240
rect 74 1236 76 1238
rect 104 1236 106 1238
rect 134 1236 136 1238
rect 164 1236 166 1238
rect 194 1236 196 1238
rect 224 1236 226 1238
rect 254 1236 256 1238
rect 284 1236 286 1238
rect 314 1236 316 1238
rect 344 1236 346 1238
rect 374 1236 376 1238
rect 404 1236 406 1238
rect 434 1236 436 1238
rect 464 1236 466 1238
rect 494 1236 496 1238
rect 524 1236 526 1238
rect 74 1230 76 1232
rect 104 1230 106 1232
rect 134 1230 136 1232
rect 164 1230 166 1232
rect 194 1230 196 1232
rect 224 1230 226 1232
rect 254 1230 256 1232
rect 284 1230 286 1232
rect 314 1230 316 1232
rect 344 1230 346 1232
rect 374 1230 376 1232
rect 404 1230 406 1232
rect 434 1230 436 1232
rect 464 1230 466 1232
rect 494 1230 496 1232
rect 524 1230 526 1232
rect 76 1228 78 1230
rect 82 1228 84 1230
rect 106 1228 108 1230
rect 112 1228 114 1230
rect 136 1228 138 1230
rect 142 1228 144 1230
rect 166 1228 168 1230
rect 172 1228 174 1230
rect 196 1228 198 1230
rect 202 1228 204 1230
rect 226 1228 228 1230
rect 232 1228 234 1230
rect 256 1228 258 1230
rect 262 1228 264 1230
rect 286 1228 288 1230
rect 292 1228 294 1230
rect 316 1228 318 1230
rect 322 1228 324 1230
rect 346 1228 348 1230
rect 352 1228 354 1230
rect 376 1228 378 1230
rect 382 1228 384 1230
rect 406 1228 408 1230
rect 412 1228 414 1230
rect 436 1228 438 1230
rect 442 1228 444 1230
rect 466 1228 468 1230
rect 472 1228 474 1230
rect 496 1228 498 1230
rect 502 1228 504 1230
rect 526 1228 528 1230
rect 532 1228 534 1230
rect 84 1226 86 1228
rect 114 1226 116 1228
rect 144 1226 146 1228
rect 174 1226 176 1228
rect 204 1226 206 1228
rect 234 1226 236 1228
rect 264 1226 266 1228
rect 294 1226 296 1228
rect 324 1226 326 1228
rect 354 1226 356 1228
rect 384 1226 386 1228
rect 414 1226 416 1228
rect 444 1226 446 1228
rect 474 1226 476 1228
rect 504 1226 506 1228
rect 534 1226 536 1228
rect 84 1220 86 1222
rect 114 1220 116 1222
rect 144 1220 146 1222
rect 174 1220 176 1222
rect 204 1220 206 1222
rect 234 1220 236 1222
rect 264 1220 266 1222
rect 294 1220 296 1222
rect 324 1220 326 1222
rect 354 1220 356 1222
rect 384 1220 386 1222
rect 414 1220 416 1222
rect 444 1220 446 1222
rect 474 1220 476 1222
rect 504 1220 506 1222
rect 534 1220 536 1222
rect 76 1218 78 1220
rect 82 1218 84 1220
rect 106 1218 108 1220
rect 112 1218 114 1220
rect 136 1218 138 1220
rect 142 1218 144 1220
rect 166 1218 168 1220
rect 172 1218 174 1220
rect 196 1218 198 1220
rect 202 1218 204 1220
rect 226 1218 228 1220
rect 232 1218 234 1220
rect 256 1218 258 1220
rect 262 1218 264 1220
rect 286 1218 288 1220
rect 292 1218 294 1220
rect 316 1218 318 1220
rect 322 1218 324 1220
rect 346 1218 348 1220
rect 352 1218 354 1220
rect 376 1218 378 1220
rect 382 1218 384 1220
rect 406 1218 408 1220
rect 412 1218 414 1220
rect 436 1218 438 1220
rect 442 1218 444 1220
rect 466 1218 468 1220
rect 472 1218 474 1220
rect 496 1218 498 1220
rect 502 1218 504 1220
rect 526 1218 528 1220
rect 532 1218 534 1220
rect 74 1216 76 1218
rect 104 1216 106 1218
rect 134 1216 136 1218
rect 164 1216 166 1218
rect 194 1216 196 1218
rect 224 1216 226 1218
rect 254 1216 256 1218
rect 284 1216 286 1218
rect 314 1216 316 1218
rect 344 1216 346 1218
rect 374 1216 376 1218
rect 404 1216 406 1218
rect 434 1216 436 1218
rect 464 1216 466 1218
rect 494 1216 496 1218
rect 524 1216 526 1218
rect 74 1210 76 1212
rect 104 1210 106 1212
rect 134 1210 136 1212
rect 164 1210 166 1212
rect 194 1210 196 1212
rect 224 1210 226 1212
rect 254 1210 256 1212
rect 284 1210 286 1212
rect 314 1210 316 1212
rect 344 1210 346 1212
rect 374 1210 376 1212
rect 404 1210 406 1212
rect 434 1210 436 1212
rect 464 1210 466 1212
rect 494 1210 496 1212
rect 524 1210 526 1212
rect 76 1208 78 1210
rect 82 1208 84 1210
rect 106 1208 108 1210
rect 112 1208 114 1210
rect 136 1208 138 1210
rect 142 1208 144 1210
rect 166 1208 168 1210
rect 172 1208 174 1210
rect 196 1208 198 1210
rect 202 1208 204 1210
rect 226 1208 228 1210
rect 232 1208 234 1210
rect 256 1208 258 1210
rect 262 1208 264 1210
rect 286 1208 288 1210
rect 292 1208 294 1210
rect 316 1208 318 1210
rect 322 1208 324 1210
rect 346 1208 348 1210
rect 352 1208 354 1210
rect 376 1208 378 1210
rect 382 1208 384 1210
rect 406 1208 408 1210
rect 412 1208 414 1210
rect 436 1208 438 1210
rect 442 1208 444 1210
rect 466 1208 468 1210
rect 472 1208 474 1210
rect 496 1208 498 1210
rect 502 1208 504 1210
rect 526 1208 528 1210
rect 532 1208 534 1210
rect 84 1206 86 1208
rect 114 1206 116 1208
rect 144 1206 146 1208
rect 174 1206 176 1208
rect 204 1206 206 1208
rect 234 1206 236 1208
rect 264 1206 266 1208
rect 294 1206 296 1208
rect 324 1206 326 1208
rect 354 1206 356 1208
rect 384 1206 386 1208
rect 414 1206 416 1208
rect 444 1206 446 1208
rect 474 1206 476 1208
rect 504 1206 506 1208
rect 534 1206 536 1208
rect 84 1200 86 1202
rect 114 1200 116 1202
rect 144 1200 146 1202
rect 174 1200 176 1202
rect 204 1200 206 1202
rect 234 1200 236 1202
rect 264 1200 266 1202
rect 294 1200 296 1202
rect 324 1200 326 1202
rect 354 1200 356 1202
rect 384 1200 386 1202
rect 414 1200 416 1202
rect 444 1200 446 1202
rect 474 1200 476 1202
rect 504 1200 506 1202
rect 534 1200 536 1202
rect 76 1198 78 1200
rect 82 1198 84 1200
rect 106 1198 108 1200
rect 112 1198 114 1200
rect 136 1198 138 1200
rect 142 1198 144 1200
rect 166 1198 168 1200
rect 172 1198 174 1200
rect 196 1198 198 1200
rect 202 1198 204 1200
rect 226 1198 228 1200
rect 232 1198 234 1200
rect 256 1198 258 1200
rect 262 1198 264 1200
rect 286 1198 288 1200
rect 292 1198 294 1200
rect 316 1198 318 1200
rect 322 1198 324 1200
rect 346 1198 348 1200
rect 352 1198 354 1200
rect 376 1198 378 1200
rect 382 1198 384 1200
rect 406 1198 408 1200
rect 412 1198 414 1200
rect 436 1198 438 1200
rect 442 1198 444 1200
rect 466 1198 468 1200
rect 472 1198 474 1200
rect 496 1198 498 1200
rect 502 1198 504 1200
rect 526 1198 528 1200
rect 532 1198 534 1200
rect 74 1196 76 1198
rect 104 1196 106 1198
rect 134 1196 136 1198
rect 164 1196 166 1198
rect 194 1196 196 1198
rect 224 1196 226 1198
rect 254 1196 256 1198
rect 284 1196 286 1198
rect 314 1196 316 1198
rect 344 1196 346 1198
rect 374 1196 376 1198
rect 404 1196 406 1198
rect 434 1196 436 1198
rect 464 1196 466 1198
rect 494 1196 496 1198
rect 524 1196 526 1198
rect 74 1190 76 1192
rect 524 1190 526 1192
rect 76 1188 78 1190
rect 82 1188 84 1190
rect 526 1188 528 1190
rect 532 1188 534 1190
rect 84 1186 86 1188
rect 534 1186 536 1188
rect 84 1180 86 1182
rect 534 1180 536 1182
rect 76 1178 78 1180
rect 82 1178 84 1180
rect 526 1178 528 1180
rect 532 1178 534 1180
rect 74 1176 76 1178
rect 524 1176 526 1178
rect 74 1170 76 1172
rect 104 1170 106 1172
rect 134 1170 136 1172
rect 164 1170 166 1172
rect 194 1170 196 1172
rect 224 1170 226 1172
rect 254 1170 256 1172
rect 284 1170 286 1172
rect 314 1170 316 1172
rect 344 1170 346 1172
rect 374 1170 376 1172
rect 404 1170 406 1172
rect 434 1170 436 1172
rect 464 1170 466 1172
rect 494 1170 496 1172
rect 524 1170 526 1172
rect 76 1168 78 1170
rect 82 1168 84 1170
rect 106 1168 108 1170
rect 112 1168 114 1170
rect 136 1168 138 1170
rect 142 1168 144 1170
rect 166 1168 168 1170
rect 172 1168 174 1170
rect 196 1168 198 1170
rect 202 1168 204 1170
rect 226 1168 228 1170
rect 232 1168 234 1170
rect 256 1168 258 1170
rect 262 1168 264 1170
rect 286 1168 288 1170
rect 292 1168 294 1170
rect 316 1168 318 1170
rect 322 1168 324 1170
rect 346 1168 348 1170
rect 352 1168 354 1170
rect 376 1168 378 1170
rect 382 1168 384 1170
rect 406 1168 408 1170
rect 412 1168 414 1170
rect 436 1168 438 1170
rect 442 1168 444 1170
rect 466 1168 468 1170
rect 472 1168 474 1170
rect 496 1168 498 1170
rect 502 1168 504 1170
rect 526 1168 528 1170
rect 532 1168 534 1170
rect 84 1166 86 1168
rect 114 1166 116 1168
rect 144 1166 146 1168
rect 174 1166 176 1168
rect 204 1166 206 1168
rect 234 1166 236 1168
rect 264 1166 266 1168
rect 294 1166 296 1168
rect 324 1166 326 1168
rect 354 1166 356 1168
rect 384 1166 386 1168
rect 414 1166 416 1168
rect 444 1166 446 1168
rect 474 1166 476 1168
rect 504 1166 506 1168
rect 534 1166 536 1168
rect 84 1160 86 1162
rect 114 1160 116 1162
rect 144 1160 146 1162
rect 174 1160 176 1162
rect 204 1160 206 1162
rect 234 1160 236 1162
rect 264 1160 266 1162
rect 294 1160 296 1162
rect 324 1160 326 1162
rect 354 1160 356 1162
rect 384 1160 386 1162
rect 414 1160 416 1162
rect 444 1160 446 1162
rect 474 1160 476 1162
rect 504 1160 506 1162
rect 534 1160 536 1162
rect 76 1158 78 1160
rect 82 1158 84 1160
rect 106 1158 108 1160
rect 112 1158 114 1160
rect 136 1158 138 1160
rect 142 1158 144 1160
rect 166 1158 168 1160
rect 172 1158 174 1160
rect 196 1158 198 1160
rect 202 1158 204 1160
rect 226 1158 228 1160
rect 232 1158 234 1160
rect 256 1158 258 1160
rect 262 1158 264 1160
rect 286 1158 288 1160
rect 292 1158 294 1160
rect 316 1158 318 1160
rect 322 1158 324 1160
rect 346 1158 348 1160
rect 352 1158 354 1160
rect 376 1158 378 1160
rect 382 1158 384 1160
rect 406 1158 408 1160
rect 412 1158 414 1160
rect 436 1158 438 1160
rect 442 1158 444 1160
rect 466 1158 468 1160
rect 472 1158 474 1160
rect 496 1158 498 1160
rect 502 1158 504 1160
rect 526 1158 528 1160
rect 532 1158 534 1160
rect 74 1156 76 1158
rect 104 1156 106 1158
rect 134 1156 136 1158
rect 164 1156 166 1158
rect 194 1156 196 1158
rect 224 1156 226 1158
rect 254 1156 256 1158
rect 284 1156 286 1158
rect 314 1156 316 1158
rect 344 1156 346 1158
rect 374 1156 376 1158
rect 404 1156 406 1158
rect 434 1156 436 1158
rect 464 1156 466 1158
rect 494 1156 496 1158
rect 524 1156 526 1158
rect 74 1150 76 1152
rect 104 1150 106 1152
rect 134 1150 136 1152
rect 164 1150 166 1152
rect 194 1150 196 1152
rect 224 1150 226 1152
rect 254 1150 256 1152
rect 284 1150 286 1152
rect 314 1150 316 1152
rect 344 1150 346 1152
rect 374 1150 376 1152
rect 404 1150 406 1152
rect 434 1150 436 1152
rect 464 1150 466 1152
rect 494 1150 496 1152
rect 524 1150 526 1152
rect 76 1148 78 1150
rect 82 1148 84 1150
rect 106 1148 108 1150
rect 112 1148 114 1150
rect 136 1148 138 1150
rect 142 1148 144 1150
rect 166 1148 168 1150
rect 172 1148 174 1150
rect 196 1148 198 1150
rect 202 1148 204 1150
rect 226 1148 228 1150
rect 232 1148 234 1150
rect 256 1148 258 1150
rect 262 1148 264 1150
rect 286 1148 288 1150
rect 292 1148 294 1150
rect 316 1148 318 1150
rect 322 1148 324 1150
rect 346 1148 348 1150
rect 352 1148 354 1150
rect 376 1148 378 1150
rect 382 1148 384 1150
rect 406 1148 408 1150
rect 412 1148 414 1150
rect 436 1148 438 1150
rect 442 1148 444 1150
rect 466 1148 468 1150
rect 472 1148 474 1150
rect 496 1148 498 1150
rect 502 1148 504 1150
rect 526 1148 528 1150
rect 532 1148 534 1150
rect 84 1146 86 1148
rect 114 1146 116 1148
rect 144 1146 146 1148
rect 174 1146 176 1148
rect 204 1146 206 1148
rect 234 1146 236 1148
rect 264 1146 266 1148
rect 294 1146 296 1148
rect 324 1146 326 1148
rect 354 1146 356 1148
rect 384 1146 386 1148
rect 414 1146 416 1148
rect 444 1146 446 1148
rect 474 1146 476 1148
rect 504 1146 506 1148
rect 534 1146 536 1148
rect 84 1140 86 1142
rect 114 1140 116 1142
rect 144 1140 146 1142
rect 174 1140 176 1142
rect 204 1140 206 1142
rect 234 1140 236 1142
rect 264 1140 266 1142
rect 294 1140 296 1142
rect 324 1140 326 1142
rect 354 1140 356 1142
rect 384 1140 386 1142
rect 414 1140 416 1142
rect 444 1140 446 1142
rect 474 1140 476 1142
rect 504 1140 506 1142
rect 534 1140 536 1142
rect 76 1138 78 1140
rect 82 1138 84 1140
rect 106 1138 108 1140
rect 112 1138 114 1140
rect 136 1138 138 1140
rect 142 1138 144 1140
rect 166 1138 168 1140
rect 172 1138 174 1140
rect 196 1138 198 1140
rect 202 1138 204 1140
rect 226 1138 228 1140
rect 232 1138 234 1140
rect 256 1138 258 1140
rect 262 1138 264 1140
rect 286 1138 288 1140
rect 292 1138 294 1140
rect 316 1138 318 1140
rect 322 1138 324 1140
rect 346 1138 348 1140
rect 352 1138 354 1140
rect 376 1138 378 1140
rect 382 1138 384 1140
rect 406 1138 408 1140
rect 412 1138 414 1140
rect 436 1138 438 1140
rect 442 1138 444 1140
rect 466 1138 468 1140
rect 472 1138 474 1140
rect 496 1138 498 1140
rect 502 1138 504 1140
rect 526 1138 528 1140
rect 532 1138 534 1140
rect 74 1136 76 1138
rect 104 1136 106 1138
rect 134 1136 136 1138
rect 164 1136 166 1138
rect 194 1136 196 1138
rect 224 1136 226 1138
rect 254 1136 256 1138
rect 284 1136 286 1138
rect 314 1136 316 1138
rect 344 1136 346 1138
rect 374 1136 376 1138
rect 404 1136 406 1138
rect 434 1136 436 1138
rect 464 1136 466 1138
rect 494 1136 496 1138
rect 524 1136 526 1138
rect 74 1130 76 1132
rect 104 1130 106 1132
rect 134 1130 136 1132
rect 164 1130 166 1132
rect 194 1130 196 1132
rect 224 1130 226 1132
rect 254 1130 256 1132
rect 284 1130 286 1132
rect 314 1130 316 1132
rect 344 1130 346 1132
rect 374 1130 376 1132
rect 404 1130 406 1132
rect 434 1130 436 1132
rect 464 1130 466 1132
rect 494 1130 496 1132
rect 524 1130 526 1132
rect 76 1128 78 1130
rect 82 1128 84 1130
rect 106 1128 108 1130
rect 112 1128 114 1130
rect 136 1128 138 1130
rect 142 1128 144 1130
rect 166 1128 168 1130
rect 172 1128 174 1130
rect 196 1128 198 1130
rect 202 1128 204 1130
rect 226 1128 228 1130
rect 232 1128 234 1130
rect 256 1128 258 1130
rect 262 1128 264 1130
rect 286 1128 288 1130
rect 292 1128 294 1130
rect 316 1128 318 1130
rect 322 1128 324 1130
rect 346 1128 348 1130
rect 352 1128 354 1130
rect 376 1128 378 1130
rect 382 1128 384 1130
rect 406 1128 408 1130
rect 412 1128 414 1130
rect 436 1128 438 1130
rect 442 1128 444 1130
rect 466 1128 468 1130
rect 472 1128 474 1130
rect 496 1128 498 1130
rect 502 1128 504 1130
rect 526 1128 528 1130
rect 532 1128 534 1130
rect 84 1126 86 1128
rect 114 1126 116 1128
rect 144 1126 146 1128
rect 174 1126 176 1128
rect 204 1126 206 1128
rect 234 1126 236 1128
rect 264 1126 266 1128
rect 294 1126 296 1128
rect 324 1126 326 1128
rect 354 1126 356 1128
rect 384 1126 386 1128
rect 414 1126 416 1128
rect 444 1126 446 1128
rect 474 1126 476 1128
rect 504 1126 506 1128
rect 534 1126 536 1128
rect 84 1120 86 1122
rect 504 1120 506 1122
rect 534 1120 536 1122
rect 86 1118 88 1120
rect 506 1118 508 1120
rect 532 1118 534 1120
rect 86 1108 88 1110
rect 506 1108 508 1110
rect 532 1108 534 1110
rect 84 1106 86 1108
rect 504 1106 506 1108
rect 534 1106 536 1108
rect 84 1100 86 1102
rect 114 1100 116 1102
rect 144 1100 146 1102
rect 174 1100 176 1102
rect 204 1100 206 1102
rect 234 1100 236 1102
rect 264 1100 266 1102
rect 294 1100 296 1102
rect 324 1100 326 1102
rect 354 1100 356 1102
rect 384 1100 386 1102
rect 414 1100 416 1102
rect 444 1100 446 1102
rect 474 1100 476 1102
rect 504 1100 506 1102
rect 534 1100 536 1102
rect 76 1098 78 1100
rect 82 1098 84 1100
rect 106 1098 108 1100
rect 112 1098 114 1100
rect 136 1098 138 1100
rect 142 1098 144 1100
rect 166 1098 168 1100
rect 172 1098 174 1100
rect 196 1098 198 1100
rect 202 1098 204 1100
rect 226 1098 228 1100
rect 232 1098 234 1100
rect 256 1098 258 1100
rect 262 1098 264 1100
rect 286 1098 288 1100
rect 292 1098 294 1100
rect 316 1098 318 1100
rect 322 1098 324 1100
rect 346 1098 348 1100
rect 352 1098 354 1100
rect 376 1098 378 1100
rect 382 1098 384 1100
rect 406 1098 408 1100
rect 412 1098 414 1100
rect 436 1098 438 1100
rect 442 1098 444 1100
rect 466 1098 468 1100
rect 472 1098 474 1100
rect 496 1098 498 1100
rect 502 1098 504 1100
rect 526 1098 528 1100
rect 532 1098 534 1100
rect 74 1096 76 1098
rect 104 1096 106 1098
rect 134 1096 136 1098
rect 164 1096 166 1098
rect 194 1096 196 1098
rect 224 1096 226 1098
rect 254 1096 256 1098
rect 284 1096 286 1098
rect 314 1096 316 1098
rect 344 1096 346 1098
rect 374 1096 376 1098
rect 404 1096 406 1098
rect 434 1096 436 1098
rect 464 1096 466 1098
rect 494 1096 496 1098
rect 524 1096 526 1098
rect 74 1090 76 1092
rect 104 1090 106 1092
rect 134 1090 136 1092
rect 164 1090 166 1092
rect 194 1090 196 1092
rect 224 1090 226 1092
rect 254 1090 256 1092
rect 284 1090 286 1092
rect 314 1090 316 1092
rect 344 1090 346 1092
rect 374 1090 376 1092
rect 404 1090 406 1092
rect 434 1090 436 1092
rect 464 1090 466 1092
rect 494 1090 496 1092
rect 524 1090 526 1092
rect 76 1088 78 1090
rect 82 1088 84 1090
rect 106 1088 108 1090
rect 112 1088 114 1090
rect 136 1088 138 1090
rect 142 1088 144 1090
rect 166 1088 168 1090
rect 172 1088 174 1090
rect 196 1088 198 1090
rect 202 1088 204 1090
rect 226 1088 228 1090
rect 232 1088 234 1090
rect 256 1088 258 1090
rect 262 1088 264 1090
rect 286 1088 288 1090
rect 292 1088 294 1090
rect 316 1088 318 1090
rect 322 1088 324 1090
rect 346 1088 348 1090
rect 352 1088 354 1090
rect 376 1088 378 1090
rect 382 1088 384 1090
rect 406 1088 408 1090
rect 412 1088 414 1090
rect 436 1088 438 1090
rect 442 1088 444 1090
rect 466 1088 468 1090
rect 472 1088 474 1090
rect 496 1088 498 1090
rect 502 1088 504 1090
rect 526 1088 528 1090
rect 532 1088 534 1090
rect 84 1086 86 1088
rect 114 1086 116 1088
rect 144 1086 146 1088
rect 174 1086 176 1088
rect 204 1086 206 1088
rect 234 1086 236 1088
rect 264 1086 266 1088
rect 294 1086 296 1088
rect 324 1086 326 1088
rect 354 1086 356 1088
rect 384 1086 386 1088
rect 414 1086 416 1088
rect 444 1086 446 1088
rect 474 1086 476 1088
rect 504 1086 506 1088
rect 534 1086 536 1088
rect 84 1080 86 1082
rect 114 1080 116 1082
rect 144 1080 146 1082
rect 174 1080 176 1082
rect 204 1080 206 1082
rect 234 1080 236 1082
rect 264 1080 266 1082
rect 294 1080 296 1082
rect 324 1080 326 1082
rect 354 1080 356 1082
rect 384 1080 386 1082
rect 414 1080 416 1082
rect 444 1080 446 1082
rect 474 1080 476 1082
rect 504 1080 506 1082
rect 534 1080 536 1082
rect 76 1078 78 1080
rect 82 1078 84 1080
rect 106 1078 108 1080
rect 112 1078 114 1080
rect 136 1078 138 1080
rect 142 1078 144 1080
rect 166 1078 168 1080
rect 172 1078 174 1080
rect 196 1078 198 1080
rect 202 1078 204 1080
rect 226 1078 228 1080
rect 232 1078 234 1080
rect 256 1078 258 1080
rect 262 1078 264 1080
rect 286 1078 288 1080
rect 292 1078 294 1080
rect 316 1078 318 1080
rect 322 1078 324 1080
rect 346 1078 348 1080
rect 352 1078 354 1080
rect 376 1078 378 1080
rect 382 1078 384 1080
rect 406 1078 408 1080
rect 412 1078 414 1080
rect 436 1078 438 1080
rect 442 1078 444 1080
rect 466 1078 468 1080
rect 472 1078 474 1080
rect 496 1078 498 1080
rect 502 1078 504 1080
rect 526 1078 528 1080
rect 532 1078 534 1080
rect 74 1076 76 1078
rect 104 1076 106 1078
rect 134 1076 136 1078
rect 164 1076 166 1078
rect 194 1076 196 1078
rect 224 1076 226 1078
rect 254 1076 256 1078
rect 284 1076 286 1078
rect 314 1076 316 1078
rect 344 1076 346 1078
rect 374 1076 376 1078
rect 404 1076 406 1078
rect 434 1076 436 1078
rect 464 1076 466 1078
rect 494 1076 496 1078
rect 524 1076 526 1078
rect 74 1070 76 1072
rect 104 1070 106 1072
rect 134 1070 136 1072
rect 164 1070 166 1072
rect 194 1070 196 1072
rect 224 1070 226 1072
rect 254 1070 256 1072
rect 284 1070 286 1072
rect 314 1070 316 1072
rect 344 1070 346 1072
rect 374 1070 376 1072
rect 404 1070 406 1072
rect 434 1070 436 1072
rect 464 1070 466 1072
rect 494 1070 496 1072
rect 524 1070 526 1072
rect 76 1068 78 1070
rect 82 1068 84 1070
rect 106 1068 108 1070
rect 112 1068 114 1070
rect 136 1068 138 1070
rect 142 1068 144 1070
rect 166 1068 168 1070
rect 172 1068 174 1070
rect 196 1068 198 1070
rect 202 1068 204 1070
rect 226 1068 228 1070
rect 232 1068 234 1070
rect 256 1068 258 1070
rect 262 1068 264 1070
rect 286 1068 288 1070
rect 292 1068 294 1070
rect 316 1068 318 1070
rect 322 1068 324 1070
rect 346 1068 348 1070
rect 352 1068 354 1070
rect 376 1068 378 1070
rect 382 1068 384 1070
rect 406 1068 408 1070
rect 412 1068 414 1070
rect 436 1068 438 1070
rect 442 1068 444 1070
rect 466 1068 468 1070
rect 472 1068 474 1070
rect 496 1068 498 1070
rect 502 1068 504 1070
rect 526 1068 528 1070
rect 532 1068 534 1070
rect 84 1066 86 1068
rect 114 1066 116 1068
rect 144 1066 146 1068
rect 174 1066 176 1068
rect 204 1066 206 1068
rect 234 1066 236 1068
rect 264 1066 266 1068
rect 294 1066 296 1068
rect 324 1066 326 1068
rect 354 1066 356 1068
rect 384 1066 386 1068
rect 414 1066 416 1068
rect 444 1066 446 1068
rect 474 1066 476 1068
rect 504 1066 506 1068
rect 534 1066 536 1068
rect 84 1060 86 1062
rect 114 1060 116 1062
rect 144 1060 146 1062
rect 174 1060 176 1062
rect 204 1060 206 1062
rect 234 1060 236 1062
rect 264 1060 266 1062
rect 294 1060 296 1062
rect 324 1060 326 1062
rect 354 1060 356 1062
rect 384 1060 386 1062
rect 414 1060 416 1062
rect 444 1060 446 1062
rect 474 1060 476 1062
rect 504 1060 506 1062
rect 534 1060 536 1062
rect 76 1058 78 1060
rect 82 1058 84 1060
rect 106 1058 108 1060
rect 112 1058 114 1060
rect 136 1058 138 1060
rect 142 1058 144 1060
rect 166 1058 168 1060
rect 172 1058 174 1060
rect 196 1058 198 1060
rect 202 1058 204 1060
rect 226 1058 228 1060
rect 232 1058 234 1060
rect 256 1058 258 1060
rect 262 1058 264 1060
rect 286 1058 288 1060
rect 292 1058 294 1060
rect 316 1058 318 1060
rect 322 1058 324 1060
rect 346 1058 348 1060
rect 352 1058 354 1060
rect 376 1058 378 1060
rect 382 1058 384 1060
rect 406 1058 408 1060
rect 412 1058 414 1060
rect 436 1058 438 1060
rect 442 1058 444 1060
rect 466 1058 468 1060
rect 472 1058 474 1060
rect 496 1058 498 1060
rect 502 1058 504 1060
rect 526 1058 528 1060
rect 532 1058 534 1060
rect 74 1056 76 1058
rect 104 1056 106 1058
rect 134 1056 136 1058
rect 164 1056 166 1058
rect 194 1056 196 1058
rect 224 1056 226 1058
rect 254 1056 256 1058
rect 284 1056 286 1058
rect 314 1056 316 1058
rect 344 1056 346 1058
rect 374 1056 376 1058
rect 404 1056 406 1058
rect 434 1056 436 1058
rect 464 1056 466 1058
rect 494 1056 496 1058
rect 524 1056 526 1058
rect 74 1050 76 1052
rect 104 1050 106 1052
rect 134 1050 136 1052
rect 164 1050 166 1052
rect 194 1050 196 1052
rect 224 1050 226 1052
rect 254 1050 256 1052
rect 284 1050 286 1052
rect 314 1050 316 1052
rect 344 1050 346 1052
rect 374 1050 376 1052
rect 404 1050 406 1052
rect 434 1050 436 1052
rect 464 1050 466 1052
rect 494 1050 496 1052
rect 524 1050 526 1052
rect 76 1048 78 1050
rect 82 1048 84 1050
rect 106 1048 108 1050
rect 112 1048 114 1050
rect 136 1048 138 1050
rect 142 1048 144 1050
rect 166 1048 168 1050
rect 172 1048 174 1050
rect 196 1048 198 1050
rect 202 1048 204 1050
rect 226 1048 228 1050
rect 232 1048 234 1050
rect 256 1048 258 1050
rect 262 1048 264 1050
rect 286 1048 288 1050
rect 292 1048 294 1050
rect 316 1048 318 1050
rect 322 1048 324 1050
rect 346 1048 348 1050
rect 352 1048 354 1050
rect 376 1048 378 1050
rect 382 1048 384 1050
rect 406 1048 408 1050
rect 412 1048 414 1050
rect 436 1048 438 1050
rect 442 1048 444 1050
rect 466 1048 468 1050
rect 472 1048 474 1050
rect 496 1048 498 1050
rect 502 1048 504 1050
rect 526 1048 528 1050
rect 532 1048 534 1050
rect 84 1046 86 1048
rect 114 1046 116 1048
rect 144 1046 146 1048
rect 174 1046 176 1048
rect 204 1046 206 1048
rect 234 1046 236 1048
rect 264 1046 266 1048
rect 294 1046 296 1048
rect 324 1046 326 1048
rect 354 1046 356 1048
rect 384 1046 386 1048
rect 414 1046 416 1048
rect 444 1046 446 1048
rect 474 1046 476 1048
rect 504 1046 506 1048
rect 534 1046 536 1048
rect 84 1040 86 1042
rect 504 1040 506 1042
rect 534 1040 536 1042
rect 76 1038 78 1040
rect 82 1038 84 1040
rect 506 1038 508 1040
rect 532 1038 534 1040
rect 74 1036 76 1038
rect 74 1030 76 1032
rect 76 1028 78 1030
rect 82 1028 84 1030
rect 506 1028 508 1030
rect 532 1028 534 1030
rect 84 1026 86 1028
rect 504 1026 506 1028
rect 534 1026 536 1028
rect 84 1020 86 1022
rect 114 1020 116 1022
rect 144 1020 146 1022
rect 174 1020 176 1022
rect 204 1020 206 1022
rect 234 1020 236 1022
rect 264 1020 266 1022
rect 294 1020 296 1022
rect 324 1020 326 1022
rect 354 1020 356 1022
rect 384 1020 386 1022
rect 414 1020 416 1022
rect 444 1020 446 1022
rect 474 1020 476 1022
rect 504 1020 506 1022
rect 534 1020 536 1022
rect 76 1018 78 1020
rect 82 1018 84 1020
rect 106 1018 108 1020
rect 112 1018 114 1020
rect 136 1018 138 1020
rect 142 1018 144 1020
rect 166 1018 168 1020
rect 172 1018 174 1020
rect 196 1018 198 1020
rect 202 1018 204 1020
rect 226 1018 228 1020
rect 232 1018 234 1020
rect 256 1018 258 1020
rect 262 1018 264 1020
rect 286 1018 288 1020
rect 292 1018 294 1020
rect 316 1018 318 1020
rect 322 1018 324 1020
rect 346 1018 348 1020
rect 352 1018 354 1020
rect 376 1018 378 1020
rect 382 1018 384 1020
rect 406 1018 408 1020
rect 412 1018 414 1020
rect 436 1018 438 1020
rect 442 1018 444 1020
rect 466 1018 468 1020
rect 472 1018 474 1020
rect 496 1018 498 1020
rect 502 1018 504 1020
rect 526 1018 528 1020
rect 532 1018 534 1020
rect 74 1016 76 1018
rect 104 1016 106 1018
rect 134 1016 136 1018
rect 164 1016 166 1018
rect 194 1016 196 1018
rect 224 1016 226 1018
rect 254 1016 256 1018
rect 284 1016 286 1018
rect 314 1016 316 1018
rect 344 1016 346 1018
rect 374 1016 376 1018
rect 404 1016 406 1018
rect 434 1016 436 1018
rect 464 1016 466 1018
rect 494 1016 496 1018
rect 524 1016 526 1018
rect 74 1010 76 1012
rect 104 1010 106 1012
rect 134 1010 136 1012
rect 164 1010 166 1012
rect 194 1010 196 1012
rect 224 1010 226 1012
rect 254 1010 256 1012
rect 284 1010 286 1012
rect 314 1010 316 1012
rect 344 1010 346 1012
rect 374 1010 376 1012
rect 404 1010 406 1012
rect 434 1010 436 1012
rect 464 1010 466 1012
rect 494 1010 496 1012
rect 524 1010 526 1012
rect 76 1008 78 1010
rect 82 1008 84 1010
rect 106 1008 108 1010
rect 112 1008 114 1010
rect 136 1008 138 1010
rect 142 1008 144 1010
rect 166 1008 168 1010
rect 172 1008 174 1010
rect 196 1008 198 1010
rect 202 1008 204 1010
rect 226 1008 228 1010
rect 232 1008 234 1010
rect 256 1008 258 1010
rect 262 1008 264 1010
rect 286 1008 288 1010
rect 292 1008 294 1010
rect 316 1008 318 1010
rect 322 1008 324 1010
rect 346 1008 348 1010
rect 352 1008 354 1010
rect 376 1008 378 1010
rect 382 1008 384 1010
rect 406 1008 408 1010
rect 412 1008 414 1010
rect 436 1008 438 1010
rect 442 1008 444 1010
rect 466 1008 468 1010
rect 472 1008 474 1010
rect 496 1008 498 1010
rect 502 1008 504 1010
rect 526 1008 528 1010
rect 532 1008 534 1010
rect 84 1006 86 1008
rect 114 1006 116 1008
rect 144 1006 146 1008
rect 174 1006 176 1008
rect 204 1006 206 1008
rect 234 1006 236 1008
rect 264 1006 266 1008
rect 294 1006 296 1008
rect 324 1006 326 1008
rect 354 1006 356 1008
rect 384 1006 386 1008
rect 414 1006 416 1008
rect 444 1006 446 1008
rect 474 1006 476 1008
rect 504 1006 506 1008
rect 534 1006 536 1008
rect 84 1000 86 1002
rect 114 1000 116 1002
rect 144 1000 146 1002
rect 174 1000 176 1002
rect 204 1000 206 1002
rect 234 1000 236 1002
rect 264 1000 266 1002
rect 294 1000 296 1002
rect 324 1000 326 1002
rect 354 1000 356 1002
rect 384 1000 386 1002
rect 414 1000 416 1002
rect 444 1000 446 1002
rect 474 1000 476 1002
rect 504 1000 506 1002
rect 534 1000 536 1002
rect 76 998 78 1000
rect 82 998 84 1000
rect 106 998 108 1000
rect 112 998 114 1000
rect 136 998 138 1000
rect 142 998 144 1000
rect 166 998 168 1000
rect 172 998 174 1000
rect 196 998 198 1000
rect 202 998 204 1000
rect 226 998 228 1000
rect 232 998 234 1000
rect 256 998 258 1000
rect 262 998 264 1000
rect 286 998 288 1000
rect 292 998 294 1000
rect 316 998 318 1000
rect 322 998 324 1000
rect 346 998 348 1000
rect 352 998 354 1000
rect 376 998 378 1000
rect 382 998 384 1000
rect 406 998 408 1000
rect 412 998 414 1000
rect 436 998 438 1000
rect 442 998 444 1000
rect 466 998 468 1000
rect 472 998 474 1000
rect 496 998 498 1000
rect 502 998 504 1000
rect 526 998 528 1000
rect 532 998 534 1000
rect 74 996 76 998
rect 104 996 106 998
rect 134 996 136 998
rect 164 996 166 998
rect 194 996 196 998
rect 224 996 226 998
rect 254 996 256 998
rect 284 996 286 998
rect 314 996 316 998
rect 344 996 346 998
rect 374 996 376 998
rect 404 996 406 998
rect 434 996 436 998
rect 464 996 466 998
rect 494 996 496 998
rect 524 996 526 998
rect 74 990 76 992
rect 104 990 106 992
rect 134 990 136 992
rect 164 990 166 992
rect 194 990 196 992
rect 224 990 226 992
rect 254 990 256 992
rect 284 990 286 992
rect 314 990 316 992
rect 344 990 346 992
rect 374 990 376 992
rect 404 990 406 992
rect 434 990 436 992
rect 464 990 466 992
rect 494 990 496 992
rect 524 990 526 992
rect 76 988 78 990
rect 82 988 84 990
rect 106 988 108 990
rect 112 988 114 990
rect 136 988 138 990
rect 142 988 144 990
rect 166 988 168 990
rect 172 988 174 990
rect 196 988 198 990
rect 202 988 204 990
rect 226 988 228 990
rect 232 988 234 990
rect 256 988 258 990
rect 262 988 264 990
rect 286 988 288 990
rect 292 988 294 990
rect 316 988 318 990
rect 322 988 324 990
rect 346 988 348 990
rect 352 988 354 990
rect 376 988 378 990
rect 382 988 384 990
rect 406 988 408 990
rect 412 988 414 990
rect 436 988 438 990
rect 442 988 444 990
rect 466 988 468 990
rect 472 988 474 990
rect 496 988 498 990
rect 502 988 504 990
rect 526 988 528 990
rect 532 988 534 990
rect 84 986 86 988
rect 114 986 116 988
rect 144 986 146 988
rect 174 986 176 988
rect 204 986 206 988
rect 234 986 236 988
rect 264 986 266 988
rect 294 986 296 988
rect 324 986 326 988
rect 354 986 356 988
rect 384 986 386 988
rect 414 986 416 988
rect 444 986 446 988
rect 474 986 476 988
rect 504 986 506 988
rect 534 986 536 988
rect 84 980 86 982
rect 114 980 116 982
rect 144 980 146 982
rect 174 980 176 982
rect 204 980 206 982
rect 234 980 236 982
rect 264 980 266 982
rect 294 980 296 982
rect 324 980 326 982
rect 354 980 356 982
rect 384 980 386 982
rect 414 980 416 982
rect 444 980 446 982
rect 474 980 476 982
rect 504 980 506 982
rect 534 980 536 982
rect 76 978 78 980
rect 82 978 84 980
rect 106 978 108 980
rect 112 978 114 980
rect 136 978 138 980
rect 142 978 144 980
rect 166 978 168 980
rect 172 978 174 980
rect 196 978 198 980
rect 202 978 204 980
rect 226 978 228 980
rect 232 978 234 980
rect 256 978 258 980
rect 262 978 264 980
rect 286 978 288 980
rect 292 978 294 980
rect 316 978 318 980
rect 322 978 324 980
rect 346 978 348 980
rect 352 978 354 980
rect 376 978 378 980
rect 382 978 384 980
rect 406 978 408 980
rect 412 978 414 980
rect 436 978 438 980
rect 442 978 444 980
rect 466 978 468 980
rect 472 978 474 980
rect 496 978 498 980
rect 502 978 504 980
rect 526 978 528 980
rect 532 978 534 980
rect 74 976 76 978
rect 104 976 106 978
rect 134 976 136 978
rect 164 976 166 978
rect 194 976 196 978
rect 224 976 226 978
rect 254 976 256 978
rect 284 976 286 978
rect 314 976 316 978
rect 344 976 346 978
rect 374 976 376 978
rect 404 976 406 978
rect 434 976 436 978
rect 464 976 466 978
rect 494 976 496 978
rect 524 976 526 978
rect 74 950 76 952
rect 104 950 106 952
rect 134 950 136 952
rect 164 950 166 952
rect 194 950 196 952
rect 224 950 226 952
rect 254 950 256 952
rect 284 950 286 952
rect 314 950 316 952
rect 344 950 346 952
rect 374 950 376 952
rect 404 950 406 952
rect 434 950 436 952
rect 464 950 466 952
rect 494 950 496 952
rect 524 950 526 952
rect 76 948 78 950
rect 82 948 84 950
rect 106 948 108 950
rect 112 948 114 950
rect 136 948 138 950
rect 142 948 144 950
rect 166 948 168 950
rect 172 948 174 950
rect 196 948 198 950
rect 202 948 204 950
rect 226 948 228 950
rect 232 948 234 950
rect 256 948 258 950
rect 262 948 264 950
rect 286 948 288 950
rect 292 948 294 950
rect 316 948 318 950
rect 322 948 324 950
rect 346 948 348 950
rect 352 948 354 950
rect 376 948 378 950
rect 382 948 384 950
rect 406 948 408 950
rect 412 948 414 950
rect 436 948 438 950
rect 442 948 444 950
rect 466 948 468 950
rect 472 948 474 950
rect 496 948 498 950
rect 502 948 504 950
rect 526 948 528 950
rect 532 948 534 950
rect 84 946 86 948
rect 114 946 116 948
rect 144 946 146 948
rect 174 946 176 948
rect 204 946 206 948
rect 234 946 236 948
rect 264 946 266 948
rect 294 946 296 948
rect 324 946 326 948
rect 354 946 356 948
rect 384 946 386 948
rect 414 946 416 948
rect 444 946 446 948
rect 474 946 476 948
rect 504 946 506 948
rect 534 946 536 948
rect 84 940 86 942
rect 114 940 116 942
rect 144 940 146 942
rect 174 940 176 942
rect 204 940 206 942
rect 234 940 236 942
rect 264 940 266 942
rect 294 940 296 942
rect 324 940 326 942
rect 354 940 356 942
rect 384 940 386 942
rect 414 940 416 942
rect 444 940 446 942
rect 474 940 476 942
rect 504 940 506 942
rect 534 940 536 942
rect 76 938 78 940
rect 82 938 84 940
rect 106 938 108 940
rect 112 938 114 940
rect 136 938 138 940
rect 142 938 144 940
rect 166 938 168 940
rect 172 938 174 940
rect 196 938 198 940
rect 202 938 204 940
rect 226 938 228 940
rect 232 938 234 940
rect 256 938 258 940
rect 262 938 264 940
rect 286 938 288 940
rect 292 938 294 940
rect 316 938 318 940
rect 322 938 324 940
rect 346 938 348 940
rect 352 938 354 940
rect 376 938 378 940
rect 382 938 384 940
rect 406 938 408 940
rect 412 938 414 940
rect 436 938 438 940
rect 442 938 444 940
rect 466 938 468 940
rect 472 938 474 940
rect 496 938 498 940
rect 502 938 504 940
rect 526 938 528 940
rect 532 938 534 940
rect 74 936 76 938
rect 104 936 106 938
rect 134 936 136 938
rect 164 936 166 938
rect 194 936 196 938
rect 224 936 226 938
rect 254 936 256 938
rect 284 936 286 938
rect 314 936 316 938
rect 344 936 346 938
rect 374 936 376 938
rect 404 936 406 938
rect 434 936 436 938
rect 464 936 466 938
rect 494 936 496 938
rect 524 936 526 938
rect 74 930 76 932
rect 104 930 106 932
rect 134 930 136 932
rect 164 930 166 932
rect 194 930 196 932
rect 224 930 226 932
rect 254 930 256 932
rect 284 930 286 932
rect 314 930 316 932
rect 344 930 346 932
rect 374 930 376 932
rect 404 930 406 932
rect 434 930 436 932
rect 464 930 466 932
rect 494 930 496 932
rect 524 930 526 932
rect 76 928 78 930
rect 82 928 84 930
rect 106 928 108 930
rect 112 928 114 930
rect 136 928 138 930
rect 142 928 144 930
rect 166 928 168 930
rect 172 928 174 930
rect 196 928 198 930
rect 202 928 204 930
rect 226 928 228 930
rect 232 928 234 930
rect 256 928 258 930
rect 262 928 264 930
rect 286 928 288 930
rect 292 928 294 930
rect 316 928 318 930
rect 322 928 324 930
rect 346 928 348 930
rect 352 928 354 930
rect 376 928 378 930
rect 382 928 384 930
rect 406 928 408 930
rect 412 928 414 930
rect 436 928 438 930
rect 442 928 444 930
rect 466 928 468 930
rect 472 928 474 930
rect 496 928 498 930
rect 502 928 504 930
rect 526 928 528 930
rect 532 928 534 930
rect 84 926 86 928
rect 114 926 116 928
rect 144 926 146 928
rect 174 926 176 928
rect 204 926 206 928
rect 234 926 236 928
rect 264 926 266 928
rect 294 926 296 928
rect 324 926 326 928
rect 354 926 356 928
rect 384 926 386 928
rect 414 926 416 928
rect 444 926 446 928
rect 474 926 476 928
rect 504 926 506 928
rect 534 926 536 928
rect 84 920 86 922
rect 114 920 116 922
rect 144 920 146 922
rect 174 920 176 922
rect 204 920 206 922
rect 234 920 236 922
rect 264 920 266 922
rect 294 920 296 922
rect 324 920 326 922
rect 354 920 356 922
rect 384 920 386 922
rect 414 920 416 922
rect 444 920 446 922
rect 474 920 476 922
rect 504 920 506 922
rect 534 920 536 922
rect 76 918 78 920
rect 82 918 84 920
rect 106 918 108 920
rect 112 918 114 920
rect 136 918 138 920
rect 142 918 144 920
rect 166 918 168 920
rect 172 918 174 920
rect 196 918 198 920
rect 202 918 204 920
rect 226 918 228 920
rect 232 918 234 920
rect 256 918 258 920
rect 262 918 264 920
rect 286 918 288 920
rect 292 918 294 920
rect 316 918 318 920
rect 322 918 324 920
rect 346 918 348 920
rect 352 918 354 920
rect 376 918 378 920
rect 382 918 384 920
rect 406 918 408 920
rect 412 918 414 920
rect 436 918 438 920
rect 442 918 444 920
rect 466 918 468 920
rect 472 918 474 920
rect 496 918 498 920
rect 502 918 504 920
rect 526 918 528 920
rect 532 918 534 920
rect 74 916 76 918
rect 104 916 106 918
rect 134 916 136 918
rect 164 916 166 918
rect 194 916 196 918
rect 224 916 226 918
rect 254 916 256 918
rect 284 916 286 918
rect 314 916 316 918
rect 344 916 346 918
rect 374 916 376 918
rect 404 916 406 918
rect 434 916 436 918
rect 464 916 466 918
rect 494 916 496 918
rect 524 916 526 918
rect 74 910 76 912
rect 104 910 106 912
rect 134 910 136 912
rect 164 910 166 912
rect 194 910 196 912
rect 224 910 226 912
rect 254 910 256 912
rect 284 910 286 912
rect 314 910 316 912
rect 344 910 346 912
rect 374 910 376 912
rect 404 910 406 912
rect 434 910 436 912
rect 464 910 466 912
rect 494 910 496 912
rect 524 910 526 912
rect 76 908 78 910
rect 82 908 84 910
rect 106 908 108 910
rect 112 908 114 910
rect 136 908 138 910
rect 142 908 144 910
rect 166 908 168 910
rect 172 908 174 910
rect 196 908 198 910
rect 202 908 204 910
rect 226 908 228 910
rect 232 908 234 910
rect 256 908 258 910
rect 262 908 264 910
rect 286 908 288 910
rect 292 908 294 910
rect 316 908 318 910
rect 322 908 324 910
rect 346 908 348 910
rect 352 908 354 910
rect 376 908 378 910
rect 382 908 384 910
rect 406 908 408 910
rect 412 908 414 910
rect 436 908 438 910
rect 442 908 444 910
rect 466 908 468 910
rect 472 908 474 910
rect 496 908 498 910
rect 502 908 504 910
rect 526 908 528 910
rect 532 908 534 910
rect 84 906 86 908
rect 114 906 116 908
rect 144 906 146 908
rect 174 906 176 908
rect 204 906 206 908
rect 234 906 236 908
rect 264 906 266 908
rect 294 906 296 908
rect 324 906 326 908
rect 354 906 356 908
rect 384 906 386 908
rect 414 906 416 908
rect 444 906 446 908
rect 474 906 476 908
rect 504 906 506 908
rect 534 906 536 908
rect 84 900 86 902
rect 114 900 116 902
rect 144 900 146 902
rect 174 900 176 902
rect 204 900 206 902
rect 234 900 236 902
rect 264 900 266 902
rect 294 900 296 902
rect 324 900 326 902
rect 354 900 356 902
rect 384 900 386 902
rect 414 900 416 902
rect 444 900 446 902
rect 474 900 476 902
rect 504 900 506 902
rect 534 900 536 902
rect 76 898 78 900
rect 82 898 84 900
rect 106 898 108 900
rect 112 898 114 900
rect 136 898 138 900
rect 142 898 144 900
rect 166 898 168 900
rect 172 898 174 900
rect 196 898 198 900
rect 202 898 204 900
rect 226 898 228 900
rect 232 898 234 900
rect 256 898 258 900
rect 262 898 264 900
rect 286 898 288 900
rect 292 898 294 900
rect 316 898 318 900
rect 322 898 324 900
rect 346 898 348 900
rect 352 898 354 900
rect 376 898 378 900
rect 382 898 384 900
rect 406 898 408 900
rect 412 898 414 900
rect 436 898 438 900
rect 442 898 444 900
rect 466 898 468 900
rect 472 898 474 900
rect 496 898 498 900
rect 502 898 504 900
rect 526 898 528 900
rect 532 898 534 900
rect 74 896 76 898
rect 104 896 106 898
rect 134 896 136 898
rect 164 896 166 898
rect 194 896 196 898
rect 224 896 226 898
rect 254 896 256 898
rect 284 896 286 898
rect 314 896 316 898
rect 344 896 346 898
rect 374 896 376 898
rect 404 896 406 898
rect 434 896 436 898
rect 464 896 466 898
rect 494 896 496 898
rect 524 896 526 898
rect 74 890 76 892
rect 104 890 106 892
rect 134 890 136 892
rect 164 890 166 892
rect 194 890 196 892
rect 224 890 226 892
rect 254 890 256 892
rect 284 890 286 892
rect 314 890 316 892
rect 344 890 346 892
rect 374 890 376 892
rect 404 890 406 892
rect 434 890 436 892
rect 464 890 466 892
rect 494 890 496 892
rect 524 890 526 892
rect 76 888 78 890
rect 82 888 84 890
rect 106 888 108 890
rect 112 888 114 890
rect 136 888 138 890
rect 142 888 144 890
rect 166 888 168 890
rect 172 888 174 890
rect 196 888 198 890
rect 202 888 204 890
rect 226 888 228 890
rect 232 888 234 890
rect 256 888 258 890
rect 262 888 264 890
rect 286 888 288 890
rect 292 888 294 890
rect 316 888 318 890
rect 322 888 324 890
rect 346 888 348 890
rect 352 888 354 890
rect 376 888 378 890
rect 382 888 384 890
rect 406 888 408 890
rect 412 888 414 890
rect 436 888 438 890
rect 442 888 444 890
rect 466 888 468 890
rect 472 888 474 890
rect 496 888 498 890
rect 502 888 504 890
rect 526 888 528 890
rect 532 888 534 890
rect 84 886 86 888
rect 114 886 116 888
rect 144 886 146 888
rect 174 886 176 888
rect 204 886 206 888
rect 234 886 236 888
rect 264 886 266 888
rect 294 886 296 888
rect 324 886 326 888
rect 354 886 356 888
rect 384 886 386 888
rect 414 886 416 888
rect 444 886 446 888
rect 474 886 476 888
rect 504 886 506 888
rect 534 886 536 888
rect 56 878 58 880
rect 62 878 64 880
rect 76 878 78 880
rect 92 878 94 880
rect 106 878 108 880
rect 122 878 124 880
rect 136 878 138 880
rect 152 878 154 880
rect 166 878 168 880
rect 182 878 184 880
rect 196 878 198 880
rect 212 878 214 880
rect 226 878 228 880
rect 242 878 244 880
rect 256 878 258 880
rect 272 878 274 880
rect 286 878 288 880
rect 302 878 304 880
rect 316 878 318 880
rect 332 878 334 880
rect 346 878 348 880
rect 362 878 364 880
rect 376 878 378 880
rect 392 878 394 880
rect 406 878 408 880
rect 422 878 424 880
rect 436 878 438 880
rect 452 878 454 880
rect 466 878 468 880
rect 482 878 484 880
rect 496 878 498 880
rect 512 878 514 880
rect 526 878 528 880
rect 542 878 544 880
rect 54 876 56 878
rect 64 876 66 878
rect 74 876 76 878
rect 94 876 96 878
rect 104 876 106 878
rect 124 876 126 878
rect 134 876 136 878
rect 154 876 156 878
rect 164 876 166 878
rect 184 876 186 878
rect 194 876 196 878
rect 214 876 216 878
rect 224 876 226 878
rect 244 876 246 878
rect 254 876 256 878
rect 274 876 276 878
rect 284 876 286 878
rect 304 876 306 878
rect 314 876 316 878
rect 334 876 336 878
rect 344 876 346 878
rect 364 876 366 878
rect 374 876 376 878
rect 394 876 396 878
rect 404 876 406 878
rect 424 876 426 878
rect 434 876 436 878
rect 454 876 456 878
rect 464 876 466 878
rect 484 876 486 878
rect 494 876 496 878
rect 514 876 516 878
rect 524 876 526 878
rect 544 876 546 878
rect 32 828 34 830
rect 62 828 64 830
rect 92 828 94 830
rect 122 828 124 830
rect 152 828 154 830
rect 182 828 184 830
rect 212 828 214 830
rect 284 828 286 830
rect 314 828 316 830
rect 386 828 388 830
rect 416 828 418 830
rect 446 828 448 830
rect 476 828 478 830
rect 506 828 508 830
rect 536 828 538 830
rect 566 828 568 830
rect 34 826 36 828
rect 40 826 42 828
rect 64 826 66 828
rect 70 826 72 828
rect 94 826 96 828
rect 100 826 102 828
rect 124 826 126 828
rect 130 826 132 828
rect 154 826 156 828
rect 160 826 162 828
rect 184 826 186 828
rect 190 826 192 828
rect 214 826 216 828
rect 220 826 222 828
rect 286 826 288 828
rect 292 826 294 828
rect 316 826 318 828
rect 322 826 324 828
rect 378 826 380 828
rect 384 826 386 828
rect 408 826 410 828
rect 414 826 416 828
rect 438 826 440 828
rect 444 826 446 828
rect 468 826 470 828
rect 474 826 476 828
rect 498 826 500 828
rect 504 826 506 828
rect 528 826 530 828
rect 534 826 536 828
rect 558 826 560 828
rect 564 826 566 828
rect 42 824 44 826
rect 72 824 74 826
rect 102 824 104 826
rect 132 824 134 826
rect 162 824 164 826
rect 192 824 194 826
rect 222 824 224 826
rect 294 824 296 826
rect 324 824 326 826
rect 376 824 378 826
rect 406 824 408 826
rect 436 824 438 826
rect 466 824 468 826
rect 496 824 498 826
rect 526 824 528 826
rect 556 824 558 826
rect 42 818 44 820
rect 72 818 74 820
rect 102 818 104 820
rect 132 818 134 820
rect 162 818 164 820
rect 192 818 194 820
rect 222 818 224 820
rect 294 818 296 820
rect 324 818 326 820
rect 376 818 378 820
rect 406 818 408 820
rect 436 818 438 820
rect 466 818 468 820
rect 496 818 498 820
rect 526 818 528 820
rect 556 818 558 820
rect 34 816 36 818
rect 40 816 42 818
rect 64 816 66 818
rect 70 816 72 818
rect 94 816 96 818
rect 100 816 102 818
rect 124 816 126 818
rect 130 816 132 818
rect 154 816 156 818
rect 160 816 162 818
rect 184 816 186 818
rect 190 816 192 818
rect 214 816 216 818
rect 220 816 222 818
rect 286 816 288 818
rect 292 816 294 818
rect 316 816 318 818
rect 322 816 324 818
rect 378 816 380 818
rect 384 816 386 818
rect 408 816 410 818
rect 414 816 416 818
rect 438 816 440 818
rect 444 816 446 818
rect 468 816 470 818
rect 474 816 476 818
rect 498 816 500 818
rect 504 816 506 818
rect 528 816 530 818
rect 534 816 536 818
rect 558 816 560 818
rect 564 816 566 818
rect 32 814 34 816
rect 62 814 64 816
rect 92 814 94 816
rect 122 814 124 816
rect 152 814 154 816
rect 182 814 184 816
rect 212 814 214 816
rect 284 814 286 816
rect 314 814 316 816
rect 386 814 388 816
rect 416 814 418 816
rect 446 814 448 816
rect 476 814 478 816
rect 506 814 508 816
rect 536 814 538 816
rect 566 814 568 816
rect 32 808 34 810
rect 62 808 64 810
rect 92 808 94 810
rect 122 808 124 810
rect 152 808 154 810
rect 182 808 184 810
rect 212 808 214 810
rect 284 808 286 810
rect 314 808 316 810
rect 386 808 388 810
rect 416 808 418 810
rect 446 808 448 810
rect 476 808 478 810
rect 506 808 508 810
rect 536 808 538 810
rect 566 808 568 810
rect 34 806 36 808
rect 40 806 42 808
rect 64 806 66 808
rect 70 806 72 808
rect 94 806 96 808
rect 100 806 102 808
rect 124 806 126 808
rect 130 806 132 808
rect 154 806 156 808
rect 160 806 162 808
rect 184 806 186 808
rect 190 806 192 808
rect 214 806 216 808
rect 220 806 222 808
rect 286 806 288 808
rect 292 806 294 808
rect 316 806 318 808
rect 322 806 324 808
rect 378 806 380 808
rect 384 806 386 808
rect 408 806 410 808
rect 414 806 416 808
rect 438 806 440 808
rect 444 806 446 808
rect 468 806 470 808
rect 474 806 476 808
rect 498 806 500 808
rect 504 806 506 808
rect 528 806 530 808
rect 534 806 536 808
rect 558 806 560 808
rect 564 806 566 808
rect 42 804 44 806
rect 72 804 74 806
rect 102 804 104 806
rect 132 804 134 806
rect 162 804 164 806
rect 192 804 194 806
rect 222 804 224 806
rect 294 804 296 806
rect 324 804 326 806
rect 376 804 378 806
rect 406 804 408 806
rect 436 804 438 806
rect 466 804 468 806
rect 496 804 498 806
rect 526 804 528 806
rect 556 804 558 806
rect 42 798 44 800
rect 72 798 74 800
rect 102 798 104 800
rect 132 798 134 800
rect 162 798 164 800
rect 192 798 194 800
rect 222 798 224 800
rect 294 798 296 800
rect 324 798 326 800
rect 376 798 378 800
rect 406 798 408 800
rect 436 798 438 800
rect 466 798 468 800
rect 496 798 498 800
rect 526 798 528 800
rect 556 798 558 800
rect 34 796 36 798
rect 40 796 42 798
rect 64 796 66 798
rect 70 796 72 798
rect 94 796 96 798
rect 100 796 102 798
rect 124 796 126 798
rect 130 796 132 798
rect 154 796 156 798
rect 160 796 162 798
rect 184 796 186 798
rect 190 796 192 798
rect 214 796 216 798
rect 220 796 222 798
rect 286 796 288 798
rect 292 796 294 798
rect 316 796 318 798
rect 322 796 324 798
rect 378 796 380 798
rect 384 796 386 798
rect 408 796 410 798
rect 414 796 416 798
rect 438 796 440 798
rect 444 796 446 798
rect 468 796 470 798
rect 474 796 476 798
rect 498 796 500 798
rect 504 796 506 798
rect 528 796 530 798
rect 534 796 536 798
rect 558 796 560 798
rect 564 796 566 798
rect 32 794 34 796
rect 62 794 64 796
rect 92 794 94 796
rect 122 794 124 796
rect 152 794 154 796
rect 182 794 184 796
rect 212 794 214 796
rect 284 794 286 796
rect 314 794 316 796
rect 386 794 388 796
rect 416 794 418 796
rect 446 794 448 796
rect 476 794 478 796
rect 506 794 508 796
rect 536 794 538 796
rect 566 794 568 796
rect 32 788 34 790
rect 62 788 64 790
rect 92 788 94 790
rect 122 788 124 790
rect 152 788 154 790
rect 182 788 184 790
rect 212 788 214 790
rect 284 788 286 790
rect 314 788 316 790
rect 386 788 388 790
rect 416 788 418 790
rect 446 788 448 790
rect 476 788 478 790
rect 506 788 508 790
rect 536 788 538 790
rect 566 788 568 790
rect 34 786 36 788
rect 40 786 42 788
rect 64 786 66 788
rect 70 786 72 788
rect 94 786 96 788
rect 100 786 102 788
rect 124 786 126 788
rect 130 786 132 788
rect 154 786 156 788
rect 160 786 162 788
rect 184 786 186 788
rect 190 786 192 788
rect 214 786 216 788
rect 220 786 222 788
rect 286 786 288 788
rect 292 786 294 788
rect 316 786 318 788
rect 322 786 324 788
rect 378 786 380 788
rect 384 786 386 788
rect 408 786 410 788
rect 414 786 416 788
rect 438 786 440 788
rect 444 786 446 788
rect 468 786 470 788
rect 474 786 476 788
rect 498 786 500 788
rect 504 786 506 788
rect 528 786 530 788
rect 534 786 536 788
rect 558 786 560 788
rect 564 786 566 788
rect 42 784 44 786
rect 72 784 74 786
rect 102 784 104 786
rect 132 784 134 786
rect 162 784 164 786
rect 192 784 194 786
rect 222 784 224 786
rect 294 784 296 786
rect 324 784 326 786
rect 376 784 378 786
rect 406 784 408 786
rect 436 784 438 786
rect 466 784 468 786
rect 496 784 498 786
rect 526 784 528 786
rect 556 784 558 786
rect 42 778 44 780
rect 72 778 74 780
rect 526 778 528 780
rect 556 778 558 780
rect 34 776 36 778
rect 40 776 42 778
rect 64 776 66 778
rect 70 776 72 778
rect 94 776 96 778
rect 110 776 112 778
rect 124 776 126 778
rect 140 776 142 778
rect 154 776 156 778
rect 170 776 172 778
rect 184 776 186 778
rect 200 776 202 778
rect 214 776 216 778
rect 230 776 232 778
rect 244 776 246 778
rect 266 776 268 778
rect 272 776 274 778
rect 286 776 288 778
rect 302 776 304 778
rect 316 776 318 778
rect 332 776 334 778
rect 354 776 356 778
rect 368 776 370 778
rect 384 776 386 778
rect 398 776 400 778
rect 414 776 416 778
rect 428 776 430 778
rect 444 776 446 778
rect 458 776 460 778
rect 474 776 476 778
rect 488 776 490 778
rect 504 776 506 778
rect 528 776 530 778
rect 534 776 536 778
rect 558 776 560 778
rect 564 776 566 778
rect 32 774 34 776
rect 62 774 64 776
rect 92 774 94 776
rect 112 774 114 776
rect 122 774 124 776
rect 142 774 144 776
rect 152 774 154 776
rect 172 774 174 776
rect 182 774 184 776
rect 202 774 204 776
rect 212 774 214 776
rect 232 774 234 776
rect 242 774 244 776
rect 264 774 266 776
rect 274 774 276 776
rect 284 774 286 776
rect 304 774 306 776
rect 314 774 316 776
rect 334 774 336 776
rect 356 774 358 776
rect 366 774 368 776
rect 386 774 388 776
rect 396 774 398 776
rect 416 774 418 776
rect 426 774 428 776
rect 446 774 448 776
rect 456 774 458 776
rect 476 774 478 776
rect 486 774 488 776
rect 506 774 508 776
rect 536 774 538 776
rect 566 774 568 776
rect 32 768 34 770
rect 62 768 64 770
rect 92 768 94 770
rect 112 768 114 770
rect 122 768 124 770
rect 142 768 144 770
rect 152 768 154 770
rect 172 768 174 770
rect 182 768 184 770
rect 202 768 204 770
rect 212 768 214 770
rect 232 768 234 770
rect 242 768 244 770
rect 264 768 266 770
rect 274 768 276 770
rect 284 768 286 770
rect 304 768 306 770
rect 314 768 316 770
rect 334 768 336 770
rect 356 768 358 770
rect 366 768 368 770
rect 386 768 388 770
rect 396 768 398 770
rect 416 768 418 770
rect 426 768 428 770
rect 446 768 448 770
rect 456 768 458 770
rect 476 768 478 770
rect 486 768 488 770
rect 506 768 508 770
rect 536 768 538 770
rect 566 768 568 770
rect 34 766 36 768
rect 40 766 42 768
rect 64 766 66 768
rect 70 766 72 768
rect 94 766 96 768
rect 110 766 112 768
rect 124 766 126 768
rect 140 766 142 768
rect 154 766 156 768
rect 170 766 172 768
rect 184 766 186 768
rect 200 766 202 768
rect 214 766 216 768
rect 230 766 232 768
rect 244 766 246 768
rect 266 766 268 768
rect 272 766 274 768
rect 286 766 288 768
rect 302 766 304 768
rect 316 766 318 768
rect 332 766 334 768
rect 354 766 356 768
rect 368 766 370 768
rect 384 766 386 768
rect 398 766 400 768
rect 414 766 416 768
rect 428 766 430 768
rect 444 766 446 768
rect 458 766 460 768
rect 474 766 476 768
rect 488 766 490 768
rect 504 766 506 768
rect 528 766 530 768
rect 534 766 536 768
rect 558 766 560 768
rect 564 766 566 768
rect 42 764 44 766
rect 72 764 74 766
rect 526 764 528 766
rect 556 764 558 766
rect 42 758 44 760
rect 72 758 74 760
rect 102 758 104 760
rect 132 758 134 760
rect 162 758 164 760
rect 192 758 194 760
rect 222 758 224 760
rect 294 758 296 760
rect 324 758 326 760
rect 376 758 378 760
rect 406 758 408 760
rect 436 758 438 760
rect 466 758 468 760
rect 496 758 498 760
rect 526 758 528 760
rect 556 758 558 760
rect 34 756 36 758
rect 40 756 42 758
rect 64 756 66 758
rect 70 756 72 758
rect 94 756 96 758
rect 100 756 102 758
rect 124 756 126 758
rect 130 756 132 758
rect 154 756 156 758
rect 160 756 162 758
rect 184 756 186 758
rect 190 756 192 758
rect 214 756 216 758
rect 220 756 222 758
rect 286 756 288 758
rect 292 756 294 758
rect 316 756 318 758
rect 322 756 324 758
rect 378 756 380 758
rect 384 756 386 758
rect 408 756 410 758
rect 414 756 416 758
rect 438 756 440 758
rect 444 756 446 758
rect 468 756 470 758
rect 474 756 476 758
rect 498 756 500 758
rect 504 756 506 758
rect 528 756 530 758
rect 534 756 536 758
rect 558 756 560 758
rect 564 756 566 758
rect 32 754 34 756
rect 62 754 64 756
rect 92 754 94 756
rect 122 754 124 756
rect 152 754 154 756
rect 182 754 184 756
rect 212 754 214 756
rect 284 754 286 756
rect 314 754 316 756
rect 386 754 388 756
rect 416 754 418 756
rect 446 754 448 756
rect 476 754 478 756
rect 506 754 508 756
rect 536 754 538 756
rect 566 754 568 756
rect 32 748 34 750
rect 62 748 64 750
rect 92 748 94 750
rect 122 748 124 750
rect 152 748 154 750
rect 182 748 184 750
rect 212 748 214 750
rect 284 748 286 750
rect 314 748 316 750
rect 386 748 388 750
rect 416 748 418 750
rect 446 748 448 750
rect 476 748 478 750
rect 506 748 508 750
rect 536 748 538 750
rect 566 748 568 750
rect 34 746 36 748
rect 40 746 42 748
rect 64 746 66 748
rect 70 746 72 748
rect 94 746 96 748
rect 100 746 102 748
rect 124 746 126 748
rect 130 746 132 748
rect 154 746 156 748
rect 160 746 162 748
rect 184 746 186 748
rect 190 746 192 748
rect 214 746 216 748
rect 220 746 222 748
rect 286 746 288 748
rect 292 746 294 748
rect 316 746 318 748
rect 322 746 324 748
rect 378 746 380 748
rect 384 746 386 748
rect 408 746 410 748
rect 414 746 416 748
rect 438 746 440 748
rect 444 746 446 748
rect 468 746 470 748
rect 474 746 476 748
rect 498 746 500 748
rect 504 746 506 748
rect 528 746 530 748
rect 534 746 536 748
rect 558 746 560 748
rect 564 746 566 748
rect 42 744 44 746
rect 72 744 74 746
rect 102 744 104 746
rect 132 744 134 746
rect 162 744 164 746
rect 192 744 194 746
rect 222 744 224 746
rect 294 744 296 746
rect 324 744 326 746
rect 376 744 378 746
rect 406 744 408 746
rect 436 744 438 746
rect 466 744 468 746
rect 496 744 498 746
rect 526 744 528 746
rect 556 744 558 746
rect 222 738 224 740
rect 294 738 296 740
rect 324 738 326 740
rect 376 738 378 740
rect 220 736 222 738
rect 286 736 288 738
rect 292 736 294 738
rect 316 736 318 738
rect 322 736 324 738
rect 378 736 380 738
rect 284 734 286 736
rect 314 734 316 736
rect 284 728 286 730
rect 314 728 316 730
rect 220 726 222 728
rect 286 726 288 728
rect 292 726 294 728
rect 316 726 318 728
rect 322 726 324 728
rect 378 726 380 728
rect 222 724 224 726
rect 294 724 296 726
rect 324 724 326 726
rect 376 724 378 726
rect 42 718 44 720
rect 72 718 74 720
rect 102 718 104 720
rect 132 718 134 720
rect 162 718 164 720
rect 192 718 194 720
rect 222 718 224 720
rect 294 718 296 720
rect 324 718 326 720
rect 376 718 378 720
rect 406 718 408 720
rect 436 718 438 720
rect 466 718 468 720
rect 496 718 498 720
rect 526 718 528 720
rect 556 718 558 720
rect 34 716 36 718
rect 40 716 42 718
rect 64 716 66 718
rect 70 716 72 718
rect 94 716 96 718
rect 100 716 102 718
rect 124 716 126 718
rect 130 716 132 718
rect 154 716 156 718
rect 160 716 162 718
rect 184 716 186 718
rect 190 716 192 718
rect 214 716 216 718
rect 220 716 222 718
rect 286 716 288 718
rect 292 716 294 718
rect 316 716 318 718
rect 322 716 324 718
rect 378 716 380 718
rect 384 716 386 718
rect 408 716 410 718
rect 414 716 416 718
rect 438 716 440 718
rect 444 716 446 718
rect 468 716 470 718
rect 474 716 476 718
rect 498 716 500 718
rect 504 716 506 718
rect 528 716 530 718
rect 534 716 536 718
rect 558 716 560 718
rect 564 716 566 718
rect 32 714 34 716
rect 62 714 64 716
rect 92 714 94 716
rect 122 714 124 716
rect 152 714 154 716
rect 182 714 184 716
rect 212 714 214 716
rect 284 714 286 716
rect 314 714 316 716
rect 386 714 388 716
rect 416 714 418 716
rect 446 714 448 716
rect 476 714 478 716
rect 506 714 508 716
rect 536 714 538 716
rect 566 714 568 716
rect 32 708 34 710
rect 62 708 64 710
rect 92 708 94 710
rect 122 708 124 710
rect 152 708 154 710
rect 182 708 184 710
rect 212 708 214 710
rect 284 708 286 710
rect 314 708 316 710
rect 386 708 388 710
rect 416 708 418 710
rect 446 708 448 710
rect 476 708 478 710
rect 506 708 508 710
rect 536 708 538 710
rect 566 708 568 710
rect 34 706 36 708
rect 40 706 42 708
rect 64 706 66 708
rect 70 706 72 708
rect 94 706 96 708
rect 100 706 102 708
rect 124 706 126 708
rect 130 706 132 708
rect 154 706 156 708
rect 160 706 162 708
rect 184 706 186 708
rect 190 706 192 708
rect 214 706 216 708
rect 220 706 222 708
rect 286 706 288 708
rect 292 706 294 708
rect 316 706 318 708
rect 322 706 324 708
rect 378 706 380 708
rect 384 706 386 708
rect 408 706 410 708
rect 414 706 416 708
rect 438 706 440 708
rect 444 706 446 708
rect 468 706 470 708
rect 474 706 476 708
rect 498 706 500 708
rect 504 706 506 708
rect 528 706 530 708
rect 534 706 536 708
rect 558 706 560 708
rect 564 706 566 708
rect 42 704 44 706
rect 72 704 74 706
rect 102 704 104 706
rect 132 704 134 706
rect 162 704 164 706
rect 192 704 194 706
rect 222 704 224 706
rect 294 704 296 706
rect 324 704 326 706
rect 376 704 378 706
rect 406 704 408 706
rect 436 704 438 706
rect 466 704 468 706
rect 496 704 498 706
rect 526 704 528 706
rect 556 704 558 706
rect 42 698 44 700
rect 72 698 74 700
rect 102 698 104 700
rect 132 698 134 700
rect 162 698 164 700
rect 192 698 194 700
rect 222 698 224 700
rect 294 698 296 700
rect 324 698 326 700
rect 376 698 378 700
rect 406 698 408 700
rect 436 698 438 700
rect 466 698 468 700
rect 496 698 498 700
rect 526 698 528 700
rect 556 698 558 700
rect 34 696 36 698
rect 40 696 42 698
rect 64 696 66 698
rect 70 696 72 698
rect 94 696 96 698
rect 100 696 102 698
rect 124 696 126 698
rect 130 696 132 698
rect 154 696 156 698
rect 160 696 162 698
rect 184 696 186 698
rect 190 696 192 698
rect 214 696 216 698
rect 220 696 222 698
rect 286 696 288 698
rect 292 696 294 698
rect 316 696 318 698
rect 322 696 324 698
rect 378 696 380 698
rect 384 696 386 698
rect 408 696 410 698
rect 414 696 416 698
rect 438 696 440 698
rect 444 696 446 698
rect 468 696 470 698
rect 474 696 476 698
rect 498 696 500 698
rect 504 696 506 698
rect 528 696 530 698
rect 534 696 536 698
rect 558 696 560 698
rect 564 696 566 698
rect 32 694 34 696
rect 62 694 64 696
rect 92 694 94 696
rect 122 694 124 696
rect 152 694 154 696
rect 182 694 184 696
rect 212 694 214 696
rect 284 694 286 696
rect 314 694 316 696
rect 386 694 388 696
rect 416 694 418 696
rect 446 694 448 696
rect 476 694 478 696
rect 506 694 508 696
rect 536 694 538 696
rect 566 694 568 696
rect 32 644 34 646
rect 62 644 64 646
rect 92 644 94 646
rect 122 644 124 646
rect 152 644 154 646
rect 182 644 184 646
rect 212 644 214 646
rect 284 644 286 646
rect 314 644 316 646
rect 386 644 388 646
rect 416 644 418 646
rect 446 644 448 646
rect 476 644 478 646
rect 506 644 508 646
rect 536 644 538 646
rect 566 644 568 646
rect 34 642 36 644
rect 40 642 42 644
rect 64 642 66 644
rect 70 642 72 644
rect 94 642 96 644
rect 100 642 102 644
rect 124 642 126 644
rect 130 642 132 644
rect 154 642 156 644
rect 160 642 162 644
rect 184 642 186 644
rect 190 642 192 644
rect 214 642 216 644
rect 220 642 222 644
rect 286 642 288 644
rect 292 642 294 644
rect 316 642 318 644
rect 322 642 324 644
rect 378 642 380 644
rect 384 642 386 644
rect 408 642 410 644
rect 414 642 416 644
rect 438 642 440 644
rect 444 642 446 644
rect 468 642 470 644
rect 474 642 476 644
rect 498 642 500 644
rect 504 642 506 644
rect 528 642 530 644
rect 534 642 536 644
rect 558 642 560 644
rect 564 642 566 644
rect 42 640 44 642
rect 72 640 74 642
rect 102 640 104 642
rect 132 640 134 642
rect 162 640 164 642
rect 192 640 194 642
rect 222 640 224 642
rect 294 640 296 642
rect 324 640 326 642
rect 376 640 378 642
rect 406 640 408 642
rect 436 640 438 642
rect 466 640 468 642
rect 496 640 498 642
rect 526 640 528 642
rect 556 640 558 642
rect 42 634 44 636
rect 72 634 74 636
rect 102 634 104 636
rect 132 634 134 636
rect 162 634 164 636
rect 192 634 194 636
rect 222 634 224 636
rect 294 634 296 636
rect 324 634 326 636
rect 376 634 378 636
rect 406 634 408 636
rect 436 634 438 636
rect 466 634 468 636
rect 496 634 498 636
rect 526 634 528 636
rect 556 634 558 636
rect 34 632 36 634
rect 40 632 42 634
rect 64 632 66 634
rect 70 632 72 634
rect 94 632 96 634
rect 100 632 102 634
rect 124 632 126 634
rect 130 632 132 634
rect 154 632 156 634
rect 160 632 162 634
rect 184 632 186 634
rect 190 632 192 634
rect 214 632 216 634
rect 220 632 222 634
rect 286 632 288 634
rect 292 632 294 634
rect 316 632 318 634
rect 322 632 324 634
rect 378 632 380 634
rect 384 632 386 634
rect 408 632 410 634
rect 414 632 416 634
rect 438 632 440 634
rect 444 632 446 634
rect 468 632 470 634
rect 474 632 476 634
rect 498 632 500 634
rect 504 632 506 634
rect 528 632 530 634
rect 534 632 536 634
rect 558 632 560 634
rect 564 632 566 634
rect 32 630 34 632
rect 62 630 64 632
rect 92 630 94 632
rect 122 630 124 632
rect 152 630 154 632
rect 182 630 184 632
rect 212 630 214 632
rect 284 630 286 632
rect 314 630 316 632
rect 386 630 388 632
rect 416 630 418 632
rect 446 630 448 632
rect 476 630 478 632
rect 506 630 508 632
rect 536 630 538 632
rect 566 630 568 632
rect 32 624 34 626
rect 62 624 64 626
rect 92 624 94 626
rect 122 624 124 626
rect 152 624 154 626
rect 182 624 184 626
rect 212 624 214 626
rect 284 624 286 626
rect 314 624 316 626
rect 386 624 388 626
rect 416 624 418 626
rect 446 624 448 626
rect 476 624 478 626
rect 506 624 508 626
rect 536 624 538 626
rect 566 624 568 626
rect 34 622 36 624
rect 40 622 42 624
rect 64 622 66 624
rect 70 622 72 624
rect 94 622 96 624
rect 100 622 102 624
rect 124 622 126 624
rect 130 622 132 624
rect 154 622 156 624
rect 160 622 162 624
rect 184 622 186 624
rect 190 622 192 624
rect 214 622 216 624
rect 220 622 222 624
rect 286 622 288 624
rect 292 622 294 624
rect 316 622 318 624
rect 322 622 324 624
rect 378 622 380 624
rect 384 622 386 624
rect 408 622 410 624
rect 414 622 416 624
rect 438 622 440 624
rect 444 622 446 624
rect 468 622 470 624
rect 474 622 476 624
rect 498 622 500 624
rect 504 622 506 624
rect 528 622 530 624
rect 534 622 536 624
rect 558 622 560 624
rect 564 622 566 624
rect 42 620 44 622
rect 72 620 74 622
rect 102 620 104 622
rect 132 620 134 622
rect 162 620 164 622
rect 192 620 194 622
rect 222 620 224 622
rect 294 620 296 622
rect 324 620 326 622
rect 376 620 378 622
rect 406 620 408 622
rect 436 620 438 622
rect 466 620 468 622
rect 496 620 498 622
rect 526 620 528 622
rect 556 620 558 622
rect 222 614 224 616
rect 294 614 296 616
rect 324 614 326 616
rect 376 614 378 616
rect 220 612 222 614
rect 286 612 288 614
rect 292 612 294 614
rect 316 612 318 614
rect 322 612 324 614
rect 378 612 380 614
rect 284 610 286 612
rect 314 610 316 612
rect 284 604 286 606
rect 314 604 316 606
rect 220 602 222 604
rect 286 602 288 604
rect 292 602 294 604
rect 316 602 318 604
rect 322 602 324 604
rect 378 602 380 604
rect 222 600 224 602
rect 294 600 296 602
rect 324 600 326 602
rect 376 600 378 602
rect 42 594 44 596
rect 72 594 74 596
rect 102 594 104 596
rect 132 594 134 596
rect 162 594 164 596
rect 192 594 194 596
rect 222 594 224 596
rect 376 594 378 596
rect 406 594 408 596
rect 436 594 438 596
rect 466 594 468 596
rect 496 594 498 596
rect 526 594 528 596
rect 556 594 558 596
rect 34 592 36 594
rect 40 592 42 594
rect 64 592 66 594
rect 70 592 72 594
rect 94 592 96 594
rect 100 592 102 594
rect 124 592 126 594
rect 130 592 132 594
rect 154 592 156 594
rect 160 592 162 594
rect 184 592 186 594
rect 190 592 192 594
rect 214 592 216 594
rect 220 592 222 594
rect 266 592 268 594
rect 272 592 274 594
rect 286 592 288 594
rect 302 592 304 594
rect 316 592 318 594
rect 332 592 334 594
rect 378 592 380 594
rect 384 592 386 594
rect 408 592 410 594
rect 414 592 416 594
rect 438 592 440 594
rect 444 592 446 594
rect 468 592 470 594
rect 474 592 476 594
rect 498 592 500 594
rect 504 592 506 594
rect 528 592 530 594
rect 534 592 536 594
rect 558 592 560 594
rect 564 592 566 594
rect 32 590 34 592
rect 62 590 64 592
rect 92 590 94 592
rect 122 590 124 592
rect 152 590 154 592
rect 182 590 184 592
rect 212 590 214 592
rect 264 590 266 592
rect 274 590 276 592
rect 284 590 286 592
rect 304 590 306 592
rect 314 590 316 592
rect 334 590 336 592
rect 386 590 388 592
rect 416 590 418 592
rect 446 590 448 592
rect 476 590 478 592
rect 506 590 508 592
rect 536 590 538 592
rect 566 590 568 592
rect 32 584 34 586
rect 62 584 64 586
rect 92 584 94 586
rect 506 584 508 586
rect 536 584 538 586
rect 566 584 568 586
rect 34 582 36 584
rect 40 582 42 584
rect 64 582 66 584
rect 70 582 72 584
rect 94 582 96 584
rect 100 582 102 584
rect 114 582 116 584
rect 130 582 132 584
rect 144 582 146 584
rect 160 582 162 584
rect 174 582 176 584
rect 190 582 192 584
rect 204 582 206 584
rect 220 582 222 584
rect 234 582 236 584
rect 240 582 242 584
rect 358 582 360 584
rect 364 582 366 584
rect 378 582 380 584
rect 394 582 396 584
rect 408 582 410 584
rect 424 582 426 584
rect 438 582 440 584
rect 454 582 456 584
rect 468 582 470 584
rect 484 582 486 584
rect 498 582 500 584
rect 504 582 506 584
rect 528 582 530 584
rect 534 582 536 584
rect 558 582 560 584
rect 564 582 566 584
rect 42 580 44 582
rect 72 580 74 582
rect 102 580 104 582
rect 112 580 114 582
rect 132 580 134 582
rect 142 580 144 582
rect 162 580 164 582
rect 172 580 174 582
rect 192 580 194 582
rect 202 580 204 582
rect 222 580 224 582
rect 232 580 234 582
rect 242 580 244 582
rect 356 580 358 582
rect 366 580 368 582
rect 376 580 378 582
rect 396 580 398 582
rect 406 580 408 582
rect 426 580 428 582
rect 436 580 438 582
rect 456 580 458 582
rect 466 580 468 582
rect 486 580 488 582
rect 496 580 498 582
rect 526 580 528 582
rect 556 580 558 582
rect 42 574 44 576
rect 72 574 74 576
rect 102 574 104 576
rect 112 574 114 576
rect 132 574 134 576
rect 142 574 144 576
rect 162 574 164 576
rect 172 574 174 576
rect 192 574 194 576
rect 202 574 204 576
rect 222 574 224 576
rect 232 574 234 576
rect 242 574 244 576
rect 264 574 266 576
rect 274 574 276 576
rect 294 574 296 576
rect 304 574 306 576
rect 324 574 326 576
rect 334 574 336 576
rect 356 574 358 576
rect 366 574 368 576
rect 376 574 378 576
rect 396 574 398 576
rect 406 574 408 576
rect 426 574 428 576
rect 436 574 438 576
rect 456 574 458 576
rect 466 574 468 576
rect 486 574 488 576
rect 496 574 498 576
rect 526 574 528 576
rect 556 574 558 576
rect 34 572 36 574
rect 40 572 42 574
rect 64 572 66 574
rect 70 572 72 574
rect 94 572 96 574
rect 100 572 102 574
rect 114 572 116 574
rect 130 572 132 574
rect 144 572 146 574
rect 160 572 162 574
rect 174 572 176 574
rect 190 572 192 574
rect 204 572 206 574
rect 220 572 222 574
rect 234 572 236 574
rect 240 572 242 574
rect 262 572 264 574
rect 276 572 278 574
rect 292 572 294 574
rect 306 572 308 574
rect 322 572 324 574
rect 336 572 338 574
rect 358 572 360 574
rect 364 572 366 574
rect 378 572 380 574
rect 394 572 396 574
rect 408 572 410 574
rect 424 572 426 574
rect 438 572 440 574
rect 454 572 456 574
rect 468 572 470 574
rect 484 572 486 574
rect 498 572 500 574
rect 504 572 506 574
rect 528 572 530 574
rect 534 572 536 574
rect 558 572 560 574
rect 564 572 566 574
rect 32 570 34 572
rect 62 570 64 572
rect 92 570 94 572
rect 506 570 508 572
rect 536 570 538 572
rect 566 570 568 572
rect 32 564 34 566
rect 62 564 64 566
rect 92 564 94 566
rect 122 564 124 566
rect 152 564 154 566
rect 182 564 184 566
rect 212 564 214 566
rect 284 564 286 566
rect 314 564 316 566
rect 386 564 388 566
rect 416 564 418 566
rect 446 564 448 566
rect 476 564 478 566
rect 506 564 508 566
rect 536 564 538 566
rect 566 564 568 566
rect 34 562 36 564
rect 40 562 42 564
rect 64 562 66 564
rect 70 562 72 564
rect 94 562 96 564
rect 100 562 102 564
rect 124 562 126 564
rect 130 562 132 564
rect 154 562 156 564
rect 160 562 162 564
rect 184 562 186 564
rect 190 562 192 564
rect 214 562 216 564
rect 220 562 222 564
rect 286 562 288 564
rect 292 562 294 564
rect 316 562 318 564
rect 322 562 324 564
rect 378 562 380 564
rect 384 562 386 564
rect 408 562 410 564
rect 414 562 416 564
rect 438 562 440 564
rect 444 562 446 564
rect 468 562 470 564
rect 474 562 476 564
rect 498 562 500 564
rect 504 562 506 564
rect 528 562 530 564
rect 534 562 536 564
rect 558 562 560 564
rect 564 562 566 564
rect 42 560 44 562
rect 72 560 74 562
rect 102 560 104 562
rect 132 560 134 562
rect 162 560 164 562
rect 192 560 194 562
rect 222 560 224 562
rect 294 560 296 562
rect 324 560 326 562
rect 376 560 378 562
rect 406 560 408 562
rect 436 560 438 562
rect 466 560 468 562
rect 496 560 498 562
rect 526 560 528 562
rect 556 560 558 562
rect 42 554 44 556
rect 72 554 74 556
rect 102 554 104 556
rect 132 554 134 556
rect 162 554 164 556
rect 192 554 194 556
rect 222 554 224 556
rect 294 554 296 556
rect 324 554 326 556
rect 376 554 378 556
rect 406 554 408 556
rect 436 554 438 556
rect 466 554 468 556
rect 496 554 498 556
rect 526 554 528 556
rect 556 554 558 556
rect 34 552 36 554
rect 40 552 42 554
rect 64 552 66 554
rect 70 552 72 554
rect 94 552 96 554
rect 100 552 102 554
rect 124 552 126 554
rect 130 552 132 554
rect 154 552 156 554
rect 160 552 162 554
rect 184 552 186 554
rect 190 552 192 554
rect 214 552 216 554
rect 220 552 222 554
rect 286 552 288 554
rect 292 552 294 554
rect 316 552 318 554
rect 322 552 324 554
rect 378 552 380 554
rect 384 552 386 554
rect 408 552 410 554
rect 414 552 416 554
rect 438 552 440 554
rect 444 552 446 554
rect 468 552 470 554
rect 474 552 476 554
rect 498 552 500 554
rect 504 552 506 554
rect 528 552 530 554
rect 534 552 536 554
rect 558 552 560 554
rect 564 552 566 554
rect 32 550 34 552
rect 62 550 64 552
rect 92 550 94 552
rect 122 550 124 552
rect 152 550 154 552
rect 182 550 184 552
rect 212 550 214 552
rect 284 550 286 552
rect 314 550 316 552
rect 386 550 388 552
rect 416 550 418 552
rect 446 550 448 552
rect 476 550 478 552
rect 506 550 508 552
rect 536 550 538 552
rect 566 550 568 552
rect 32 544 34 546
rect 62 544 64 546
rect 92 544 94 546
rect 122 544 124 546
rect 152 544 154 546
rect 182 544 184 546
rect 212 544 214 546
rect 284 544 286 546
rect 314 544 316 546
rect 386 544 388 546
rect 416 544 418 546
rect 446 544 448 546
rect 476 544 478 546
rect 506 544 508 546
rect 536 544 538 546
rect 566 544 568 546
rect 34 542 36 544
rect 40 542 42 544
rect 64 542 66 544
rect 70 542 72 544
rect 94 542 96 544
rect 100 542 102 544
rect 124 542 126 544
rect 130 542 132 544
rect 154 542 156 544
rect 160 542 162 544
rect 184 542 186 544
rect 190 542 192 544
rect 214 542 216 544
rect 220 542 222 544
rect 286 542 288 544
rect 292 542 294 544
rect 316 542 318 544
rect 322 542 324 544
rect 378 542 380 544
rect 384 542 386 544
rect 408 542 410 544
rect 414 542 416 544
rect 438 542 440 544
rect 444 542 446 544
rect 468 542 470 544
rect 474 542 476 544
rect 498 542 500 544
rect 504 542 506 544
rect 528 542 530 544
rect 534 542 536 544
rect 558 542 560 544
rect 564 542 566 544
rect 42 540 44 542
rect 72 540 74 542
rect 102 540 104 542
rect 132 540 134 542
rect 162 540 164 542
rect 192 540 194 542
rect 222 540 224 542
rect 294 540 296 542
rect 324 540 326 542
rect 376 540 378 542
rect 406 540 408 542
rect 436 540 438 542
rect 466 540 468 542
rect 496 540 498 542
rect 526 540 528 542
rect 556 540 558 542
rect 42 534 44 536
rect 72 534 74 536
rect 102 534 104 536
rect 132 534 134 536
rect 162 534 164 536
rect 192 534 194 536
rect 222 534 224 536
rect 294 534 296 536
rect 324 534 326 536
rect 376 534 378 536
rect 406 534 408 536
rect 436 534 438 536
rect 466 534 468 536
rect 496 534 498 536
rect 526 534 528 536
rect 556 534 558 536
rect 34 532 36 534
rect 40 532 42 534
rect 64 532 66 534
rect 70 532 72 534
rect 94 532 96 534
rect 100 532 102 534
rect 124 532 126 534
rect 130 532 132 534
rect 154 532 156 534
rect 160 532 162 534
rect 184 532 186 534
rect 190 532 192 534
rect 214 532 216 534
rect 220 532 222 534
rect 286 532 288 534
rect 292 532 294 534
rect 316 532 318 534
rect 322 532 324 534
rect 378 532 380 534
rect 384 532 386 534
rect 408 532 410 534
rect 414 532 416 534
rect 438 532 440 534
rect 444 532 446 534
rect 468 532 470 534
rect 474 532 476 534
rect 498 532 500 534
rect 504 532 506 534
rect 528 532 530 534
rect 534 532 536 534
rect 558 532 560 534
rect 564 532 566 534
rect 32 530 34 532
rect 62 530 64 532
rect 92 530 94 532
rect 122 530 124 532
rect 152 530 154 532
rect 182 530 184 532
rect 212 530 214 532
rect 284 530 286 532
rect 314 530 316 532
rect 386 530 388 532
rect 416 530 418 532
rect 446 530 448 532
rect 476 530 478 532
rect 506 530 508 532
rect 536 530 538 532
rect 566 530 568 532
rect 586 514 596 516
rect 584 512 596 514
rect 586 508 588 512
rect 588 506 590 508
rect 40 460 42 462
rect 50 460 52 462
rect 60 460 62 462
rect 80 460 82 462
rect 90 460 92 462
rect 110 460 112 462
rect 120 460 122 462
rect 140 460 142 462
rect 150 460 152 462
rect 170 460 172 462
rect 180 460 182 462
rect 200 460 202 462
rect 210 460 212 462
rect 230 460 232 462
rect 240 460 242 462
rect 260 460 262 462
rect 270 460 272 462
rect 290 460 292 462
rect 300 460 302 462
rect 320 460 322 462
rect 330 460 332 462
rect 350 460 352 462
rect 360 460 362 462
rect 380 460 382 462
rect 390 460 392 462
rect 410 460 412 462
rect 420 460 422 462
rect 440 460 442 462
rect 450 460 452 462
rect 470 460 472 462
rect 480 460 482 462
rect 500 460 502 462
rect 510 460 512 462
rect 530 460 532 462
rect 540 460 542 462
rect 560 460 562 462
rect 42 458 44 460
rect 48 458 50 460
rect 62 458 64 460
rect 78 458 80 460
rect 92 458 94 460
rect 108 458 110 460
rect 122 458 124 460
rect 138 458 140 460
rect 152 458 154 460
rect 168 458 170 460
rect 182 458 184 460
rect 198 458 200 460
rect 212 458 214 460
rect 228 458 230 460
rect 242 458 244 460
rect 258 458 260 460
rect 272 458 274 460
rect 288 458 290 460
rect 302 458 304 460
rect 318 458 320 460
rect 332 458 334 460
rect 348 458 350 460
rect 362 458 364 460
rect 378 458 380 460
rect 392 458 394 460
rect 408 458 410 460
rect 422 458 424 460
rect 438 458 440 460
rect 452 458 454 460
rect 468 458 470 460
rect 482 458 484 460
rect 498 458 500 460
rect 512 458 514 460
rect 528 458 530 460
rect 542 458 544 460
rect 558 458 560 460
rect 70 450 72 452
rect 100 450 102 452
rect 130 450 132 452
rect 160 450 162 452
rect 190 450 192 452
rect 220 450 222 452
rect 250 450 252 452
rect 280 450 282 452
rect 310 450 312 452
rect 340 450 342 452
rect 370 450 372 452
rect 400 450 402 452
rect 430 450 432 452
rect 460 450 462 452
rect 490 450 492 452
rect 520 450 522 452
rect 550 450 552 452
rect 62 448 64 450
rect 68 448 70 450
rect 92 448 94 450
rect 98 448 100 450
rect 122 448 124 450
rect 128 448 130 450
rect 152 448 154 450
rect 158 448 160 450
rect 182 448 184 450
rect 188 448 190 450
rect 212 448 214 450
rect 218 448 220 450
rect 242 448 244 450
rect 248 448 250 450
rect 272 448 274 450
rect 278 448 280 450
rect 302 448 304 450
rect 308 448 310 450
rect 332 448 334 450
rect 338 448 340 450
rect 362 448 364 450
rect 368 448 370 450
rect 392 448 394 450
rect 398 448 400 450
rect 422 448 424 450
rect 428 448 430 450
rect 452 448 454 450
rect 458 448 460 450
rect 482 448 484 450
rect 488 448 490 450
rect 512 448 514 450
rect 518 448 520 450
rect 542 448 544 450
rect 548 448 550 450
rect 60 446 62 448
rect 90 446 92 448
rect 120 446 122 448
rect 150 446 152 448
rect 180 446 182 448
rect 210 446 212 448
rect 240 446 242 448
rect 270 446 272 448
rect 300 446 302 448
rect 330 446 332 448
rect 360 446 362 448
rect 390 446 392 448
rect 420 446 422 448
rect 450 446 452 448
rect 480 446 482 448
rect 510 446 512 448
rect 540 446 542 448
rect 60 440 62 442
rect 90 440 92 442
rect 120 440 122 442
rect 150 440 152 442
rect 180 440 182 442
rect 210 440 212 442
rect 240 440 242 442
rect 270 440 272 442
rect 300 440 302 442
rect 330 440 332 442
rect 360 440 362 442
rect 390 440 392 442
rect 420 440 422 442
rect 450 440 452 442
rect 480 440 482 442
rect 510 440 512 442
rect 540 440 542 442
rect 62 438 64 440
rect 68 438 70 440
rect 92 438 94 440
rect 98 438 100 440
rect 122 438 124 440
rect 128 438 130 440
rect 152 438 154 440
rect 158 438 160 440
rect 182 438 184 440
rect 188 438 190 440
rect 212 438 214 440
rect 218 438 220 440
rect 242 438 244 440
rect 248 438 250 440
rect 272 438 274 440
rect 278 438 280 440
rect 302 438 304 440
rect 308 438 310 440
rect 332 438 334 440
rect 338 438 340 440
rect 362 438 364 440
rect 368 438 370 440
rect 392 438 394 440
rect 398 438 400 440
rect 422 438 424 440
rect 428 438 430 440
rect 452 438 454 440
rect 458 438 460 440
rect 482 438 484 440
rect 488 438 490 440
rect 512 438 514 440
rect 518 438 520 440
rect 542 438 544 440
rect 548 438 550 440
rect 70 436 72 438
rect 100 436 102 438
rect 130 436 132 438
rect 160 436 162 438
rect 190 436 192 438
rect 220 436 222 438
rect 250 436 252 438
rect 280 436 282 438
rect 310 436 312 438
rect 340 436 342 438
rect 370 436 372 438
rect 400 436 402 438
rect 430 436 432 438
rect 460 436 462 438
rect 490 436 492 438
rect 520 436 522 438
rect 550 436 552 438
rect 70 430 72 432
rect 100 430 102 432
rect 130 430 132 432
rect 160 430 162 432
rect 190 430 192 432
rect 220 430 222 432
rect 250 430 252 432
rect 280 430 282 432
rect 310 430 312 432
rect 340 430 342 432
rect 370 430 372 432
rect 400 430 402 432
rect 430 430 432 432
rect 460 430 462 432
rect 490 430 492 432
rect 520 430 522 432
rect 550 430 552 432
rect 62 428 64 430
rect 68 428 70 430
rect 92 428 94 430
rect 98 428 100 430
rect 122 428 124 430
rect 128 428 130 430
rect 152 428 154 430
rect 158 428 160 430
rect 182 428 184 430
rect 188 428 190 430
rect 212 428 214 430
rect 218 428 220 430
rect 242 428 244 430
rect 248 428 250 430
rect 272 428 274 430
rect 278 428 280 430
rect 302 428 304 430
rect 308 428 310 430
rect 332 428 334 430
rect 338 428 340 430
rect 362 428 364 430
rect 368 428 370 430
rect 392 428 394 430
rect 398 428 400 430
rect 422 428 424 430
rect 428 428 430 430
rect 452 428 454 430
rect 458 428 460 430
rect 482 428 484 430
rect 488 428 490 430
rect 512 428 514 430
rect 518 428 520 430
rect 542 428 544 430
rect 548 428 550 430
rect 60 426 62 428
rect 90 426 92 428
rect 120 426 122 428
rect 150 426 152 428
rect 180 426 182 428
rect 210 426 212 428
rect 240 426 242 428
rect 270 426 272 428
rect 300 426 302 428
rect 330 426 332 428
rect 360 426 362 428
rect 390 426 392 428
rect 420 426 422 428
rect 450 426 452 428
rect 480 426 482 428
rect 510 426 512 428
rect 540 426 542 428
rect 60 420 62 422
rect 90 420 92 422
rect 120 420 122 422
rect 150 420 152 422
rect 180 420 182 422
rect 210 420 212 422
rect 240 420 242 422
rect 270 420 272 422
rect 300 420 302 422
rect 330 420 332 422
rect 360 420 362 422
rect 390 420 392 422
rect 420 420 422 422
rect 450 420 452 422
rect 480 420 482 422
rect 510 420 512 422
rect 540 420 542 422
rect 62 418 64 420
rect 68 418 70 420
rect 92 418 94 420
rect 98 418 100 420
rect 122 418 124 420
rect 128 418 130 420
rect 152 418 154 420
rect 158 418 160 420
rect 182 418 184 420
rect 188 418 190 420
rect 212 418 214 420
rect 218 418 220 420
rect 242 418 244 420
rect 248 418 250 420
rect 272 418 274 420
rect 278 418 280 420
rect 302 418 304 420
rect 308 418 310 420
rect 332 418 334 420
rect 338 418 340 420
rect 362 418 364 420
rect 368 418 370 420
rect 392 418 394 420
rect 398 418 400 420
rect 422 418 424 420
rect 428 418 430 420
rect 452 418 454 420
rect 458 418 460 420
rect 482 418 484 420
rect 488 418 490 420
rect 512 418 514 420
rect 518 418 520 420
rect 542 418 544 420
rect 548 418 550 420
rect 70 416 72 418
rect 100 416 102 418
rect 130 416 132 418
rect 160 416 162 418
rect 190 416 192 418
rect 220 416 222 418
rect 250 416 252 418
rect 280 416 282 418
rect 310 416 312 418
rect 340 416 342 418
rect 370 416 372 418
rect 400 416 402 418
rect 430 416 432 418
rect 460 416 462 418
rect 490 416 492 418
rect 520 416 522 418
rect 550 416 552 418
rect 70 410 72 412
rect 100 410 102 412
rect 130 410 132 412
rect 160 410 162 412
rect 190 410 192 412
rect 220 410 222 412
rect 250 410 252 412
rect 280 410 282 412
rect 310 410 312 412
rect 340 410 342 412
rect 370 410 372 412
rect 400 410 402 412
rect 430 410 432 412
rect 460 410 462 412
rect 490 410 492 412
rect 520 410 522 412
rect 550 410 552 412
rect 62 408 64 410
rect 68 408 70 410
rect 92 408 94 410
rect 98 408 100 410
rect 122 408 124 410
rect 128 408 130 410
rect 152 408 154 410
rect 158 408 160 410
rect 182 408 184 410
rect 188 408 190 410
rect 212 408 214 410
rect 218 408 220 410
rect 242 408 244 410
rect 248 408 250 410
rect 272 408 274 410
rect 278 408 280 410
rect 302 408 304 410
rect 308 408 310 410
rect 332 408 334 410
rect 338 408 340 410
rect 362 408 364 410
rect 368 408 370 410
rect 392 408 394 410
rect 398 408 400 410
rect 422 408 424 410
rect 428 408 430 410
rect 452 408 454 410
rect 458 408 460 410
rect 482 408 484 410
rect 488 408 490 410
rect 512 408 514 410
rect 518 408 520 410
rect 542 408 544 410
rect 548 408 550 410
rect 60 406 62 408
rect 90 406 92 408
rect 120 406 122 408
rect 150 406 152 408
rect 180 406 182 408
rect 210 406 212 408
rect 240 406 242 408
rect 270 406 272 408
rect 300 406 302 408
rect 330 406 332 408
rect 360 406 362 408
rect 390 406 392 408
rect 420 406 422 408
rect 450 406 452 408
rect 480 406 482 408
rect 510 406 512 408
rect 540 406 542 408
rect 60 400 62 402
rect 90 400 92 402
rect 120 400 122 402
rect 150 400 152 402
rect 180 400 182 402
rect 210 400 212 402
rect 240 400 242 402
rect 270 400 272 402
rect 300 400 302 402
rect 330 400 332 402
rect 360 400 362 402
rect 390 400 392 402
rect 420 400 422 402
rect 450 400 452 402
rect 480 400 482 402
rect 510 400 512 402
rect 540 400 542 402
rect 62 398 64 400
rect 68 398 70 400
rect 92 398 94 400
rect 98 398 100 400
rect 122 398 124 400
rect 128 398 130 400
rect 152 398 154 400
rect 158 398 160 400
rect 182 398 184 400
rect 188 398 190 400
rect 212 398 214 400
rect 218 398 220 400
rect 242 398 244 400
rect 248 398 250 400
rect 272 398 274 400
rect 278 398 280 400
rect 302 398 304 400
rect 308 398 310 400
rect 332 398 334 400
rect 338 398 340 400
rect 362 398 364 400
rect 368 398 370 400
rect 392 398 394 400
rect 398 398 400 400
rect 422 398 424 400
rect 428 398 430 400
rect 452 398 454 400
rect 458 398 460 400
rect 482 398 484 400
rect 488 398 490 400
rect 512 398 514 400
rect 518 398 520 400
rect 542 398 544 400
rect 548 398 550 400
rect 70 396 72 398
rect 100 396 102 398
rect 130 396 132 398
rect 160 396 162 398
rect 190 396 192 398
rect 220 396 222 398
rect 250 396 252 398
rect 280 396 282 398
rect 310 396 312 398
rect 340 396 342 398
rect 370 396 372 398
rect 400 396 402 398
rect 430 396 432 398
rect 460 396 462 398
rect 490 396 492 398
rect 520 396 522 398
rect 550 396 552 398
rect 100 390 102 392
rect 520 390 522 392
rect 550 390 552 392
rect 98 388 100 390
rect 518 388 520 390
rect 542 388 544 390
rect 548 388 550 390
rect 540 386 542 388
rect 540 380 542 382
rect 98 378 100 380
rect 518 378 520 380
rect 542 378 544 380
rect 548 378 550 380
rect 100 376 102 378
rect 520 376 522 378
rect 550 376 552 378
rect 70 370 72 372
rect 100 370 102 372
rect 130 370 132 372
rect 160 370 162 372
rect 190 370 192 372
rect 220 370 222 372
rect 250 370 252 372
rect 280 370 282 372
rect 310 370 312 372
rect 340 370 342 372
rect 370 370 372 372
rect 400 370 402 372
rect 430 370 432 372
rect 460 370 462 372
rect 490 370 492 372
rect 520 370 522 372
rect 550 370 552 372
rect 62 368 64 370
rect 68 368 70 370
rect 92 368 94 370
rect 98 368 100 370
rect 122 368 124 370
rect 128 368 130 370
rect 152 368 154 370
rect 158 368 160 370
rect 182 368 184 370
rect 188 368 190 370
rect 212 368 214 370
rect 218 368 220 370
rect 242 368 244 370
rect 248 368 250 370
rect 272 368 274 370
rect 278 368 280 370
rect 302 368 304 370
rect 308 368 310 370
rect 332 368 334 370
rect 338 368 340 370
rect 362 368 364 370
rect 368 368 370 370
rect 392 368 394 370
rect 398 368 400 370
rect 422 368 424 370
rect 428 368 430 370
rect 452 368 454 370
rect 458 368 460 370
rect 482 368 484 370
rect 488 368 490 370
rect 512 368 514 370
rect 518 368 520 370
rect 542 368 544 370
rect 548 368 550 370
rect 60 366 62 368
rect 90 366 92 368
rect 120 366 122 368
rect 150 366 152 368
rect 180 366 182 368
rect 210 366 212 368
rect 240 366 242 368
rect 270 366 272 368
rect 300 366 302 368
rect 330 366 332 368
rect 360 366 362 368
rect 390 366 392 368
rect 420 366 422 368
rect 450 366 452 368
rect 480 366 482 368
rect 510 366 512 368
rect 540 366 542 368
rect 60 360 62 362
rect 90 360 92 362
rect 120 360 122 362
rect 150 360 152 362
rect 180 360 182 362
rect 210 360 212 362
rect 240 360 242 362
rect 270 360 272 362
rect 300 360 302 362
rect 330 360 332 362
rect 360 360 362 362
rect 390 360 392 362
rect 420 360 422 362
rect 450 360 452 362
rect 480 360 482 362
rect 510 360 512 362
rect 540 360 542 362
rect 62 358 64 360
rect 68 358 70 360
rect 92 358 94 360
rect 98 358 100 360
rect 122 358 124 360
rect 128 358 130 360
rect 152 358 154 360
rect 158 358 160 360
rect 182 358 184 360
rect 188 358 190 360
rect 212 358 214 360
rect 218 358 220 360
rect 242 358 244 360
rect 248 358 250 360
rect 272 358 274 360
rect 278 358 280 360
rect 302 358 304 360
rect 308 358 310 360
rect 332 358 334 360
rect 338 358 340 360
rect 362 358 364 360
rect 368 358 370 360
rect 392 358 394 360
rect 398 358 400 360
rect 422 358 424 360
rect 428 358 430 360
rect 452 358 454 360
rect 458 358 460 360
rect 482 358 484 360
rect 488 358 490 360
rect 512 358 514 360
rect 518 358 520 360
rect 542 358 544 360
rect 548 358 550 360
rect 70 356 72 358
rect 100 356 102 358
rect 130 356 132 358
rect 160 356 162 358
rect 190 356 192 358
rect 220 356 222 358
rect 250 356 252 358
rect 280 356 282 358
rect 310 356 312 358
rect 340 356 342 358
rect 370 356 372 358
rect 400 356 402 358
rect 430 356 432 358
rect 460 356 462 358
rect 490 356 492 358
rect 520 356 522 358
rect 550 356 552 358
rect 70 350 72 352
rect 100 350 102 352
rect 130 350 132 352
rect 160 350 162 352
rect 190 350 192 352
rect 220 350 222 352
rect 250 350 252 352
rect 280 350 282 352
rect 310 350 312 352
rect 340 350 342 352
rect 370 350 372 352
rect 400 350 402 352
rect 430 350 432 352
rect 460 350 462 352
rect 490 350 492 352
rect 520 350 522 352
rect 550 350 552 352
rect 62 348 64 350
rect 68 348 70 350
rect 92 348 94 350
rect 98 348 100 350
rect 122 348 124 350
rect 128 348 130 350
rect 152 348 154 350
rect 158 348 160 350
rect 182 348 184 350
rect 188 348 190 350
rect 212 348 214 350
rect 218 348 220 350
rect 242 348 244 350
rect 248 348 250 350
rect 272 348 274 350
rect 278 348 280 350
rect 302 348 304 350
rect 308 348 310 350
rect 332 348 334 350
rect 338 348 340 350
rect 362 348 364 350
rect 368 348 370 350
rect 392 348 394 350
rect 398 348 400 350
rect 422 348 424 350
rect 428 348 430 350
rect 452 348 454 350
rect 458 348 460 350
rect 482 348 484 350
rect 488 348 490 350
rect 512 348 514 350
rect 518 348 520 350
rect 542 348 544 350
rect 548 348 550 350
rect 60 346 62 348
rect 90 346 92 348
rect 120 346 122 348
rect 150 346 152 348
rect 180 346 182 348
rect 210 346 212 348
rect 240 346 242 348
rect 270 346 272 348
rect 300 346 302 348
rect 330 346 332 348
rect 360 346 362 348
rect 390 346 392 348
rect 420 346 422 348
rect 450 346 452 348
rect 480 346 482 348
rect 510 346 512 348
rect 540 346 542 348
rect 60 340 62 342
rect 90 340 92 342
rect 120 340 122 342
rect 150 340 152 342
rect 180 340 182 342
rect 210 340 212 342
rect 240 340 242 342
rect 270 340 272 342
rect 300 340 302 342
rect 330 340 332 342
rect 360 340 362 342
rect 390 340 392 342
rect 420 340 422 342
rect 450 340 452 342
rect 480 340 482 342
rect 510 340 512 342
rect 540 340 542 342
rect 62 338 64 340
rect 68 338 70 340
rect 92 338 94 340
rect 98 338 100 340
rect 122 338 124 340
rect 128 338 130 340
rect 152 338 154 340
rect 158 338 160 340
rect 182 338 184 340
rect 188 338 190 340
rect 212 338 214 340
rect 218 338 220 340
rect 242 338 244 340
rect 248 338 250 340
rect 272 338 274 340
rect 278 338 280 340
rect 302 338 304 340
rect 308 338 310 340
rect 332 338 334 340
rect 338 338 340 340
rect 362 338 364 340
rect 368 338 370 340
rect 392 338 394 340
rect 398 338 400 340
rect 422 338 424 340
rect 428 338 430 340
rect 452 338 454 340
rect 458 338 460 340
rect 482 338 484 340
rect 488 338 490 340
rect 512 338 514 340
rect 518 338 520 340
rect 542 338 544 340
rect 548 338 550 340
rect 70 336 72 338
rect 100 336 102 338
rect 130 336 132 338
rect 160 336 162 338
rect 190 336 192 338
rect 220 336 222 338
rect 250 336 252 338
rect 280 336 282 338
rect 310 336 312 338
rect 340 336 342 338
rect 370 336 372 338
rect 400 336 402 338
rect 430 336 432 338
rect 460 336 462 338
rect 490 336 492 338
rect 520 336 522 338
rect 550 336 552 338
rect 70 330 72 332
rect 100 330 102 332
rect 130 330 132 332
rect 160 330 162 332
rect 190 330 192 332
rect 220 330 222 332
rect 250 330 252 332
rect 280 330 282 332
rect 310 330 312 332
rect 340 330 342 332
rect 370 330 372 332
rect 400 330 402 332
rect 430 330 432 332
rect 460 330 462 332
rect 490 330 492 332
rect 520 330 522 332
rect 550 330 552 332
rect 62 328 64 330
rect 68 328 70 330
rect 92 328 94 330
rect 98 328 100 330
rect 122 328 124 330
rect 128 328 130 330
rect 152 328 154 330
rect 158 328 160 330
rect 182 328 184 330
rect 188 328 190 330
rect 212 328 214 330
rect 218 328 220 330
rect 242 328 244 330
rect 248 328 250 330
rect 272 328 274 330
rect 278 328 280 330
rect 302 328 304 330
rect 308 328 310 330
rect 332 328 334 330
rect 338 328 340 330
rect 362 328 364 330
rect 368 328 370 330
rect 392 328 394 330
rect 398 328 400 330
rect 422 328 424 330
rect 428 328 430 330
rect 452 328 454 330
rect 458 328 460 330
rect 482 328 484 330
rect 488 328 490 330
rect 512 328 514 330
rect 518 328 520 330
rect 542 328 544 330
rect 548 328 550 330
rect 60 326 62 328
rect 90 326 92 328
rect 120 326 122 328
rect 150 326 152 328
rect 180 326 182 328
rect 210 326 212 328
rect 240 326 242 328
rect 270 326 272 328
rect 300 326 302 328
rect 330 326 332 328
rect 360 326 362 328
rect 390 326 392 328
rect 420 326 422 328
rect 450 326 452 328
rect 480 326 482 328
rect 510 326 512 328
rect 540 326 542 328
rect 60 320 62 322
rect 90 320 92 322
rect 120 320 122 322
rect 150 320 152 322
rect 180 320 182 322
rect 210 320 212 322
rect 240 320 242 322
rect 270 320 272 322
rect 300 320 302 322
rect 330 320 332 322
rect 360 320 362 322
rect 390 320 392 322
rect 420 320 422 322
rect 450 320 452 322
rect 480 320 482 322
rect 510 320 512 322
rect 540 320 542 322
rect 62 318 64 320
rect 68 318 70 320
rect 92 318 94 320
rect 98 318 100 320
rect 122 318 124 320
rect 128 318 130 320
rect 152 318 154 320
rect 158 318 160 320
rect 182 318 184 320
rect 188 318 190 320
rect 212 318 214 320
rect 218 318 220 320
rect 242 318 244 320
rect 248 318 250 320
rect 272 318 274 320
rect 278 318 280 320
rect 302 318 304 320
rect 308 318 310 320
rect 332 318 334 320
rect 338 318 340 320
rect 362 318 364 320
rect 368 318 370 320
rect 392 318 394 320
rect 398 318 400 320
rect 422 318 424 320
rect 428 318 430 320
rect 452 318 454 320
rect 458 318 460 320
rect 482 318 484 320
rect 488 318 490 320
rect 512 318 514 320
rect 518 318 520 320
rect 542 318 544 320
rect 548 318 550 320
rect 70 316 72 318
rect 100 316 102 318
rect 130 316 132 318
rect 160 316 162 318
rect 190 316 192 318
rect 220 316 222 318
rect 250 316 252 318
rect 280 316 282 318
rect 310 316 312 318
rect 340 316 342 318
rect 370 316 372 318
rect 400 316 402 318
rect 430 316 432 318
rect 460 316 462 318
rect 490 316 492 318
rect 520 316 522 318
rect 550 316 552 318
rect 70 310 72 312
rect 520 310 522 312
rect 550 310 552 312
rect 62 308 64 310
rect 68 308 70 310
rect 512 308 514 310
rect 518 308 520 310
rect 542 308 544 310
rect 548 308 550 310
rect 60 306 62 308
rect 510 306 512 308
rect 540 306 542 308
rect 60 300 62 302
rect 510 300 512 302
rect 540 300 542 302
rect 62 298 64 300
rect 68 298 70 300
rect 512 298 514 300
rect 518 298 520 300
rect 542 298 544 300
rect 548 298 550 300
rect 70 296 72 298
rect 520 296 522 298
rect 550 296 552 298
rect 70 290 72 292
rect 100 290 102 292
rect 130 290 132 292
rect 160 290 162 292
rect 190 290 192 292
rect 220 290 222 292
rect 250 290 252 292
rect 280 290 282 292
rect 310 290 312 292
rect 340 290 342 292
rect 370 290 372 292
rect 400 290 402 292
rect 430 290 432 292
rect 460 290 462 292
rect 490 290 492 292
rect 520 290 522 292
rect 550 290 552 292
rect 62 288 64 290
rect 68 288 70 290
rect 92 288 94 290
rect 98 288 100 290
rect 122 288 124 290
rect 128 288 130 290
rect 152 288 154 290
rect 158 288 160 290
rect 182 288 184 290
rect 188 288 190 290
rect 212 288 214 290
rect 218 288 220 290
rect 242 288 244 290
rect 248 288 250 290
rect 272 288 274 290
rect 278 288 280 290
rect 302 288 304 290
rect 308 288 310 290
rect 332 288 334 290
rect 338 288 340 290
rect 362 288 364 290
rect 368 288 370 290
rect 392 288 394 290
rect 398 288 400 290
rect 422 288 424 290
rect 428 288 430 290
rect 452 288 454 290
rect 458 288 460 290
rect 482 288 484 290
rect 488 288 490 290
rect 512 288 514 290
rect 518 288 520 290
rect 542 288 544 290
rect 548 288 550 290
rect 60 286 62 288
rect 90 286 92 288
rect 120 286 122 288
rect 150 286 152 288
rect 180 286 182 288
rect 210 286 212 288
rect 240 286 242 288
rect 270 286 272 288
rect 300 286 302 288
rect 330 286 332 288
rect 360 286 362 288
rect 390 286 392 288
rect 420 286 422 288
rect 450 286 452 288
rect 480 286 482 288
rect 510 286 512 288
rect 540 286 542 288
rect 60 280 62 282
rect 90 280 92 282
rect 120 280 122 282
rect 150 280 152 282
rect 180 280 182 282
rect 210 280 212 282
rect 240 280 242 282
rect 270 280 272 282
rect 300 280 302 282
rect 330 280 332 282
rect 360 280 362 282
rect 390 280 392 282
rect 420 280 422 282
rect 450 280 452 282
rect 480 280 482 282
rect 510 280 512 282
rect 540 280 542 282
rect 62 278 64 280
rect 68 278 70 280
rect 92 278 94 280
rect 98 278 100 280
rect 122 278 124 280
rect 128 278 130 280
rect 152 278 154 280
rect 158 278 160 280
rect 182 278 184 280
rect 188 278 190 280
rect 212 278 214 280
rect 218 278 220 280
rect 242 278 244 280
rect 248 278 250 280
rect 272 278 274 280
rect 278 278 280 280
rect 302 278 304 280
rect 308 278 310 280
rect 332 278 334 280
rect 338 278 340 280
rect 362 278 364 280
rect 368 278 370 280
rect 392 278 394 280
rect 398 278 400 280
rect 422 278 424 280
rect 428 278 430 280
rect 452 278 454 280
rect 458 278 460 280
rect 482 278 484 280
rect 488 278 490 280
rect 512 278 514 280
rect 518 278 520 280
rect 542 278 544 280
rect 548 278 550 280
rect 70 276 72 278
rect 100 276 102 278
rect 130 276 132 278
rect 160 276 162 278
rect 190 276 192 278
rect 220 276 222 278
rect 250 276 252 278
rect 280 276 282 278
rect 310 276 312 278
rect 340 276 342 278
rect 370 276 372 278
rect 400 276 402 278
rect 430 276 432 278
rect 460 276 462 278
rect 490 276 492 278
rect 520 276 522 278
rect 550 276 552 278
rect 70 270 72 272
rect 100 270 102 272
rect 130 270 132 272
rect 160 270 162 272
rect 190 270 192 272
rect 220 270 222 272
rect 250 270 252 272
rect 280 270 282 272
rect 310 270 312 272
rect 340 270 342 272
rect 370 270 372 272
rect 400 270 402 272
rect 430 270 432 272
rect 460 270 462 272
rect 490 270 492 272
rect 520 270 522 272
rect 550 270 552 272
rect 62 268 64 270
rect 68 268 70 270
rect 92 268 94 270
rect 98 268 100 270
rect 122 268 124 270
rect 128 268 130 270
rect 152 268 154 270
rect 158 268 160 270
rect 182 268 184 270
rect 188 268 190 270
rect 212 268 214 270
rect 218 268 220 270
rect 242 268 244 270
rect 248 268 250 270
rect 272 268 274 270
rect 278 268 280 270
rect 302 268 304 270
rect 308 268 310 270
rect 332 268 334 270
rect 338 268 340 270
rect 362 268 364 270
rect 368 268 370 270
rect 392 268 394 270
rect 398 268 400 270
rect 422 268 424 270
rect 428 268 430 270
rect 452 268 454 270
rect 458 268 460 270
rect 482 268 484 270
rect 488 268 490 270
rect 512 268 514 270
rect 518 268 520 270
rect 542 268 544 270
rect 548 268 550 270
rect 60 266 62 268
rect 90 266 92 268
rect 120 266 122 268
rect 150 266 152 268
rect 180 266 182 268
rect 210 266 212 268
rect 240 266 242 268
rect 270 266 272 268
rect 300 266 302 268
rect 330 266 332 268
rect 360 266 362 268
rect 390 266 392 268
rect 420 266 422 268
rect 450 266 452 268
rect 480 266 482 268
rect 510 266 512 268
rect 540 266 542 268
rect 60 260 62 262
rect 90 260 92 262
rect 120 260 122 262
rect 150 260 152 262
rect 180 260 182 262
rect 210 260 212 262
rect 240 260 242 262
rect 270 260 272 262
rect 300 260 302 262
rect 330 260 332 262
rect 360 260 362 262
rect 390 260 392 262
rect 420 260 422 262
rect 450 260 452 262
rect 480 260 482 262
rect 510 260 512 262
rect 540 260 542 262
rect 62 258 64 260
rect 68 258 70 260
rect 92 258 94 260
rect 98 258 100 260
rect 122 258 124 260
rect 128 258 130 260
rect 152 258 154 260
rect 158 258 160 260
rect 182 258 184 260
rect 188 258 190 260
rect 212 258 214 260
rect 218 258 220 260
rect 242 258 244 260
rect 248 258 250 260
rect 272 258 274 260
rect 278 258 280 260
rect 302 258 304 260
rect 308 258 310 260
rect 332 258 334 260
rect 338 258 340 260
rect 362 258 364 260
rect 368 258 370 260
rect 392 258 394 260
rect 398 258 400 260
rect 422 258 424 260
rect 428 258 430 260
rect 452 258 454 260
rect 458 258 460 260
rect 482 258 484 260
rect 488 258 490 260
rect 512 258 514 260
rect 518 258 520 260
rect 542 258 544 260
rect 548 258 550 260
rect 70 256 72 258
rect 100 256 102 258
rect 130 256 132 258
rect 160 256 162 258
rect 190 256 192 258
rect 220 256 222 258
rect 250 256 252 258
rect 280 256 282 258
rect 310 256 312 258
rect 340 256 342 258
rect 370 256 372 258
rect 400 256 402 258
rect 430 256 432 258
rect 460 256 462 258
rect 490 256 492 258
rect 520 256 522 258
rect 550 256 552 258
rect 70 250 72 252
rect 100 250 102 252
rect 130 250 132 252
rect 160 250 162 252
rect 190 250 192 252
rect 220 250 222 252
rect 250 250 252 252
rect 280 250 282 252
rect 310 250 312 252
rect 340 250 342 252
rect 370 250 372 252
rect 400 250 402 252
rect 430 250 432 252
rect 460 250 462 252
rect 490 250 492 252
rect 520 250 522 252
rect 550 250 552 252
rect 62 248 64 250
rect 68 248 70 250
rect 92 248 94 250
rect 98 248 100 250
rect 122 248 124 250
rect 128 248 130 250
rect 152 248 154 250
rect 158 248 160 250
rect 182 248 184 250
rect 188 248 190 250
rect 212 248 214 250
rect 218 248 220 250
rect 242 248 244 250
rect 248 248 250 250
rect 272 248 274 250
rect 278 248 280 250
rect 302 248 304 250
rect 308 248 310 250
rect 332 248 334 250
rect 338 248 340 250
rect 362 248 364 250
rect 368 248 370 250
rect 392 248 394 250
rect 398 248 400 250
rect 422 248 424 250
rect 428 248 430 250
rect 452 248 454 250
rect 458 248 460 250
rect 482 248 484 250
rect 488 248 490 250
rect 512 248 514 250
rect 518 248 520 250
rect 542 248 544 250
rect 548 248 550 250
rect 60 246 62 248
rect 90 246 92 248
rect 120 246 122 248
rect 150 246 152 248
rect 180 246 182 248
rect 210 246 212 248
rect 240 246 242 248
rect 270 246 272 248
rect 300 246 302 248
rect 330 246 332 248
rect 360 246 362 248
rect 390 246 392 248
rect 420 246 422 248
rect 450 246 452 248
rect 480 246 482 248
rect 510 246 512 248
rect 540 246 542 248
rect 60 240 62 242
rect 90 240 92 242
rect 510 240 512 242
rect 540 240 542 242
rect 62 238 64 240
rect 88 238 90 240
rect 508 238 510 240
rect 542 238 544 240
rect 548 238 550 240
rect 550 236 552 238
rect 550 230 552 232
rect 62 228 64 230
rect 88 228 90 230
rect 508 228 510 230
rect 542 228 544 230
rect 548 228 550 230
rect 60 226 62 228
rect 90 226 92 228
rect 510 226 512 228
rect 540 226 542 228
rect 60 220 62 222
rect 90 220 92 222
rect 120 220 122 222
rect 150 220 152 222
rect 180 220 182 222
rect 210 220 212 222
rect 240 220 242 222
rect 270 220 272 222
rect 300 220 302 222
rect 330 220 332 222
rect 360 220 362 222
rect 390 220 392 222
rect 420 220 422 222
rect 450 220 452 222
rect 480 220 482 222
rect 510 220 512 222
rect 540 220 542 222
rect 62 218 64 220
rect 68 218 70 220
rect 92 218 94 220
rect 98 218 100 220
rect 122 218 124 220
rect 128 218 130 220
rect 152 218 154 220
rect 158 218 160 220
rect 182 218 184 220
rect 188 218 190 220
rect 212 218 214 220
rect 218 218 220 220
rect 242 218 244 220
rect 248 218 250 220
rect 272 218 274 220
rect 278 218 280 220
rect 302 218 304 220
rect 308 218 310 220
rect 332 218 334 220
rect 338 218 340 220
rect 362 218 364 220
rect 368 218 370 220
rect 392 218 394 220
rect 398 218 400 220
rect 422 218 424 220
rect 428 218 430 220
rect 452 218 454 220
rect 458 218 460 220
rect 482 218 484 220
rect 488 218 490 220
rect 512 218 514 220
rect 518 218 520 220
rect 542 218 544 220
rect 548 218 550 220
rect 70 216 72 218
rect 100 216 102 218
rect 130 216 132 218
rect 160 216 162 218
rect 190 216 192 218
rect 220 216 222 218
rect 250 216 252 218
rect 280 216 282 218
rect 310 216 312 218
rect 340 216 342 218
rect 370 216 372 218
rect 400 216 402 218
rect 430 216 432 218
rect 460 216 462 218
rect 490 216 492 218
rect 520 216 522 218
rect 550 216 552 218
rect 70 210 72 212
rect 100 210 102 212
rect 130 210 132 212
rect 160 210 162 212
rect 190 210 192 212
rect 220 210 222 212
rect 250 210 252 212
rect 280 210 282 212
rect 310 210 312 212
rect 340 210 342 212
rect 370 210 372 212
rect 400 210 402 212
rect 430 210 432 212
rect 460 210 462 212
rect 490 210 492 212
rect 520 210 522 212
rect 550 210 552 212
rect 62 208 64 210
rect 68 208 70 210
rect 92 208 94 210
rect 98 208 100 210
rect 122 208 124 210
rect 128 208 130 210
rect 152 208 154 210
rect 158 208 160 210
rect 182 208 184 210
rect 188 208 190 210
rect 212 208 214 210
rect 218 208 220 210
rect 242 208 244 210
rect 248 208 250 210
rect 272 208 274 210
rect 278 208 280 210
rect 302 208 304 210
rect 308 208 310 210
rect 332 208 334 210
rect 338 208 340 210
rect 362 208 364 210
rect 368 208 370 210
rect 392 208 394 210
rect 398 208 400 210
rect 422 208 424 210
rect 428 208 430 210
rect 452 208 454 210
rect 458 208 460 210
rect 482 208 484 210
rect 488 208 490 210
rect 512 208 514 210
rect 518 208 520 210
rect 542 208 544 210
rect 548 208 550 210
rect 60 206 62 208
rect 90 206 92 208
rect 120 206 122 208
rect 150 206 152 208
rect 180 206 182 208
rect 210 206 212 208
rect 240 206 242 208
rect 270 206 272 208
rect 300 206 302 208
rect 330 206 332 208
rect 360 206 362 208
rect 390 206 392 208
rect 420 206 422 208
rect 450 206 452 208
rect 480 206 482 208
rect 510 206 512 208
rect 540 206 542 208
rect 60 200 62 202
rect 90 200 92 202
rect 120 200 122 202
rect 150 200 152 202
rect 180 200 182 202
rect 210 200 212 202
rect 240 200 242 202
rect 270 200 272 202
rect 300 200 302 202
rect 330 200 332 202
rect 360 200 362 202
rect 390 200 392 202
rect 420 200 422 202
rect 450 200 452 202
rect 480 200 482 202
rect 510 200 512 202
rect 540 200 542 202
rect 62 198 64 200
rect 68 198 70 200
rect 92 198 94 200
rect 98 198 100 200
rect 122 198 124 200
rect 128 198 130 200
rect 152 198 154 200
rect 158 198 160 200
rect 182 198 184 200
rect 188 198 190 200
rect 212 198 214 200
rect 218 198 220 200
rect 242 198 244 200
rect 248 198 250 200
rect 272 198 274 200
rect 278 198 280 200
rect 302 198 304 200
rect 308 198 310 200
rect 332 198 334 200
rect 338 198 340 200
rect 362 198 364 200
rect 368 198 370 200
rect 392 198 394 200
rect 398 198 400 200
rect 422 198 424 200
rect 428 198 430 200
rect 452 198 454 200
rect 458 198 460 200
rect 482 198 484 200
rect 488 198 490 200
rect 512 198 514 200
rect 518 198 520 200
rect 542 198 544 200
rect 548 198 550 200
rect 70 196 72 198
rect 100 196 102 198
rect 130 196 132 198
rect 160 196 162 198
rect 190 196 192 198
rect 220 196 222 198
rect 250 196 252 198
rect 280 196 282 198
rect 310 196 312 198
rect 340 196 342 198
rect 370 196 372 198
rect 400 196 402 198
rect 430 196 432 198
rect 460 196 462 198
rect 490 196 492 198
rect 520 196 522 198
rect 550 196 552 198
rect 70 190 72 192
rect 100 190 102 192
rect 130 190 132 192
rect 160 190 162 192
rect 190 190 192 192
rect 220 190 222 192
rect 250 190 252 192
rect 280 190 282 192
rect 310 190 312 192
rect 340 190 342 192
rect 370 190 372 192
rect 400 190 402 192
rect 430 190 432 192
rect 460 190 462 192
rect 490 190 492 192
rect 520 190 522 192
rect 550 190 552 192
rect 62 188 64 190
rect 68 188 70 190
rect 92 188 94 190
rect 98 188 100 190
rect 122 188 124 190
rect 128 188 130 190
rect 152 188 154 190
rect 158 188 160 190
rect 182 188 184 190
rect 188 188 190 190
rect 212 188 214 190
rect 218 188 220 190
rect 242 188 244 190
rect 248 188 250 190
rect 272 188 274 190
rect 278 188 280 190
rect 302 188 304 190
rect 308 188 310 190
rect 332 188 334 190
rect 338 188 340 190
rect 362 188 364 190
rect 368 188 370 190
rect 392 188 394 190
rect 398 188 400 190
rect 422 188 424 190
rect 428 188 430 190
rect 452 188 454 190
rect 458 188 460 190
rect 482 188 484 190
rect 488 188 490 190
rect 512 188 514 190
rect 518 188 520 190
rect 542 188 544 190
rect 548 188 550 190
rect 60 186 62 188
rect 90 186 92 188
rect 120 186 122 188
rect 150 186 152 188
rect 180 186 182 188
rect 210 186 212 188
rect 240 186 242 188
rect 270 186 272 188
rect 300 186 302 188
rect 330 186 332 188
rect 360 186 362 188
rect 390 186 392 188
rect 420 186 422 188
rect 450 186 452 188
rect 480 186 482 188
rect 510 186 512 188
rect 540 186 542 188
rect 60 180 62 182
rect 90 180 92 182
rect 120 180 122 182
rect 150 180 152 182
rect 180 180 182 182
rect 210 180 212 182
rect 240 180 242 182
rect 270 180 272 182
rect 300 180 302 182
rect 330 180 332 182
rect 360 180 362 182
rect 390 180 392 182
rect 420 180 422 182
rect 450 180 452 182
rect 480 180 482 182
rect 510 180 512 182
rect 540 180 542 182
rect 62 178 64 180
rect 68 178 70 180
rect 92 178 94 180
rect 98 178 100 180
rect 122 178 124 180
rect 128 178 130 180
rect 152 178 154 180
rect 158 178 160 180
rect 182 178 184 180
rect 188 178 190 180
rect 212 178 214 180
rect 218 178 220 180
rect 242 178 244 180
rect 248 178 250 180
rect 272 178 274 180
rect 278 178 280 180
rect 302 178 304 180
rect 308 178 310 180
rect 332 178 334 180
rect 338 178 340 180
rect 362 178 364 180
rect 368 178 370 180
rect 392 178 394 180
rect 398 178 400 180
rect 422 178 424 180
rect 428 178 430 180
rect 452 178 454 180
rect 458 178 460 180
rect 482 178 484 180
rect 488 178 490 180
rect 512 178 514 180
rect 518 178 520 180
rect 542 178 544 180
rect 548 178 550 180
rect 70 176 72 178
rect 100 176 102 178
rect 130 176 132 178
rect 160 176 162 178
rect 190 176 192 178
rect 220 176 222 178
rect 250 176 252 178
rect 280 176 282 178
rect 310 176 312 178
rect 340 176 342 178
rect 370 176 372 178
rect 400 176 402 178
rect 430 176 432 178
rect 460 176 462 178
rect 490 176 492 178
rect 520 176 522 178
rect 550 176 552 178
rect 70 170 72 172
rect 100 170 102 172
rect 130 170 132 172
rect 160 170 162 172
rect 190 170 192 172
rect 220 170 222 172
rect 250 170 252 172
rect 280 170 282 172
rect 310 170 312 172
rect 340 170 342 172
rect 370 170 372 172
rect 400 170 402 172
rect 430 170 432 172
rect 460 170 462 172
rect 490 170 492 172
rect 520 170 522 172
rect 550 170 552 172
rect 62 168 64 170
rect 68 168 70 170
rect 92 168 94 170
rect 98 168 100 170
rect 122 168 124 170
rect 128 168 130 170
rect 152 168 154 170
rect 158 168 160 170
rect 182 168 184 170
rect 188 168 190 170
rect 212 168 214 170
rect 218 168 220 170
rect 242 168 244 170
rect 248 168 250 170
rect 272 168 274 170
rect 278 168 280 170
rect 302 168 304 170
rect 308 168 310 170
rect 332 168 334 170
rect 338 168 340 170
rect 362 168 364 170
rect 368 168 370 170
rect 392 168 394 170
rect 398 168 400 170
rect 422 168 424 170
rect 428 168 430 170
rect 452 168 454 170
rect 458 168 460 170
rect 482 168 484 170
rect 488 168 490 170
rect 512 168 514 170
rect 518 168 520 170
rect 542 168 544 170
rect 548 168 550 170
rect 60 166 62 168
rect 90 166 92 168
rect 120 166 122 168
rect 150 166 152 168
rect 180 166 182 168
rect 210 166 212 168
rect 240 166 242 168
rect 270 166 272 168
rect 300 166 302 168
rect 330 166 332 168
rect 360 166 362 168
rect 390 166 392 168
rect 420 166 422 168
rect 450 166 452 168
rect 480 166 482 168
rect 510 166 512 168
rect 540 166 542 168
rect 60 160 62 162
rect 90 160 92 162
rect 510 160 512 162
rect 540 160 542 162
rect 62 158 64 160
rect 68 158 70 160
rect 92 158 94 160
rect 508 158 510 160
rect 542 158 544 160
rect 548 158 550 160
rect 70 156 72 158
rect 550 156 552 158
rect 70 150 72 152
rect 550 150 552 152
rect 62 148 64 150
rect 68 148 70 150
rect 92 148 94 150
rect 508 148 510 150
rect 542 148 544 150
rect 548 148 550 150
rect 60 146 62 148
rect 90 146 92 148
rect 510 146 512 148
rect 540 146 542 148
rect 60 140 62 142
rect 90 140 92 142
rect 120 140 122 142
rect 150 140 152 142
rect 180 140 182 142
rect 210 140 212 142
rect 240 140 242 142
rect 270 140 272 142
rect 300 140 302 142
rect 330 140 332 142
rect 360 140 362 142
rect 390 140 392 142
rect 420 140 422 142
rect 450 140 452 142
rect 480 140 482 142
rect 510 140 512 142
rect 540 140 542 142
rect 62 138 64 140
rect 68 138 70 140
rect 92 138 94 140
rect 98 138 100 140
rect 122 138 124 140
rect 128 138 130 140
rect 152 138 154 140
rect 158 138 160 140
rect 182 138 184 140
rect 188 138 190 140
rect 212 138 214 140
rect 218 138 220 140
rect 242 138 244 140
rect 248 138 250 140
rect 272 138 274 140
rect 278 138 280 140
rect 302 138 304 140
rect 308 138 310 140
rect 332 138 334 140
rect 338 138 340 140
rect 362 138 364 140
rect 368 138 370 140
rect 392 138 394 140
rect 398 138 400 140
rect 422 138 424 140
rect 428 138 430 140
rect 452 138 454 140
rect 458 138 460 140
rect 482 138 484 140
rect 488 138 490 140
rect 512 138 514 140
rect 518 138 520 140
rect 542 138 544 140
rect 548 138 550 140
rect 70 136 72 138
rect 100 136 102 138
rect 130 136 132 138
rect 160 136 162 138
rect 190 136 192 138
rect 220 136 222 138
rect 250 136 252 138
rect 280 136 282 138
rect 310 136 312 138
rect 340 136 342 138
rect 370 136 372 138
rect 400 136 402 138
rect 430 136 432 138
rect 460 136 462 138
rect 490 136 492 138
rect 520 136 522 138
rect 550 136 552 138
rect 70 130 72 132
rect 100 130 102 132
rect 130 130 132 132
rect 160 130 162 132
rect 190 130 192 132
rect 220 130 222 132
rect 250 130 252 132
rect 280 130 282 132
rect 310 130 312 132
rect 340 130 342 132
rect 370 130 372 132
rect 400 130 402 132
rect 430 130 432 132
rect 460 130 462 132
rect 490 130 492 132
rect 520 130 522 132
rect 550 130 552 132
rect 62 128 64 130
rect 68 128 70 130
rect 92 128 94 130
rect 98 128 100 130
rect 122 128 124 130
rect 128 128 130 130
rect 152 128 154 130
rect 158 128 160 130
rect 182 128 184 130
rect 188 128 190 130
rect 212 128 214 130
rect 218 128 220 130
rect 242 128 244 130
rect 248 128 250 130
rect 272 128 274 130
rect 278 128 280 130
rect 302 128 304 130
rect 308 128 310 130
rect 332 128 334 130
rect 338 128 340 130
rect 362 128 364 130
rect 368 128 370 130
rect 392 128 394 130
rect 398 128 400 130
rect 422 128 424 130
rect 428 128 430 130
rect 452 128 454 130
rect 458 128 460 130
rect 482 128 484 130
rect 488 128 490 130
rect 512 128 514 130
rect 518 128 520 130
rect 542 128 544 130
rect 548 128 550 130
rect 60 126 62 128
rect 90 126 92 128
rect 120 126 122 128
rect 150 126 152 128
rect 180 126 182 128
rect 210 126 212 128
rect 240 126 242 128
rect 270 126 272 128
rect 300 126 302 128
rect 330 126 332 128
rect 360 126 362 128
rect 390 126 392 128
rect 420 126 422 128
rect 450 126 452 128
rect 480 126 482 128
rect 510 126 512 128
rect 540 126 542 128
rect 60 120 62 122
rect 90 120 92 122
rect 120 120 122 122
rect 150 120 152 122
rect 180 120 182 122
rect 210 120 212 122
rect 240 120 242 122
rect 270 120 272 122
rect 300 120 302 122
rect 330 120 332 122
rect 360 120 362 122
rect 390 120 392 122
rect 420 120 422 122
rect 450 120 452 122
rect 480 120 482 122
rect 510 120 512 122
rect 540 120 542 122
rect 62 118 64 120
rect 68 118 70 120
rect 92 118 94 120
rect 98 118 100 120
rect 122 118 124 120
rect 128 118 130 120
rect 152 118 154 120
rect 158 118 160 120
rect 182 118 184 120
rect 188 118 190 120
rect 212 118 214 120
rect 218 118 220 120
rect 242 118 244 120
rect 248 118 250 120
rect 272 118 274 120
rect 278 118 280 120
rect 302 118 304 120
rect 308 118 310 120
rect 332 118 334 120
rect 338 118 340 120
rect 362 118 364 120
rect 368 118 370 120
rect 392 118 394 120
rect 398 118 400 120
rect 422 118 424 120
rect 428 118 430 120
rect 452 118 454 120
rect 458 118 460 120
rect 482 118 484 120
rect 488 118 490 120
rect 512 118 514 120
rect 518 118 520 120
rect 542 118 544 120
rect 548 118 550 120
rect 70 116 72 118
rect 100 116 102 118
rect 130 116 132 118
rect 160 116 162 118
rect 190 116 192 118
rect 220 116 222 118
rect 250 116 252 118
rect 280 116 282 118
rect 310 116 312 118
rect 340 116 342 118
rect 370 116 372 118
rect 400 116 402 118
rect 430 116 432 118
rect 460 116 462 118
rect 490 116 492 118
rect 520 116 522 118
rect 550 116 552 118
rect 70 110 72 112
rect 100 110 102 112
rect 130 110 132 112
rect 160 110 162 112
rect 190 110 192 112
rect 220 110 222 112
rect 250 110 252 112
rect 280 110 282 112
rect 310 110 312 112
rect 340 110 342 112
rect 370 110 372 112
rect 400 110 402 112
rect 430 110 432 112
rect 460 110 462 112
rect 490 110 492 112
rect 520 110 522 112
rect 550 110 552 112
rect 62 108 64 110
rect 68 108 70 110
rect 92 108 94 110
rect 98 108 100 110
rect 122 108 124 110
rect 128 108 130 110
rect 152 108 154 110
rect 158 108 160 110
rect 182 108 184 110
rect 188 108 190 110
rect 212 108 214 110
rect 218 108 220 110
rect 242 108 244 110
rect 248 108 250 110
rect 272 108 274 110
rect 278 108 280 110
rect 302 108 304 110
rect 308 108 310 110
rect 332 108 334 110
rect 338 108 340 110
rect 362 108 364 110
rect 368 108 370 110
rect 392 108 394 110
rect 398 108 400 110
rect 422 108 424 110
rect 428 108 430 110
rect 452 108 454 110
rect 458 108 460 110
rect 482 108 484 110
rect 488 108 490 110
rect 512 108 514 110
rect 518 108 520 110
rect 542 108 544 110
rect 548 108 550 110
rect 60 106 62 108
rect 90 106 92 108
rect 120 106 122 108
rect 150 106 152 108
rect 180 106 182 108
rect 210 106 212 108
rect 240 106 242 108
rect 270 106 272 108
rect 300 106 302 108
rect 330 106 332 108
rect 360 106 362 108
rect 390 106 392 108
rect 420 106 422 108
rect 450 106 452 108
rect 480 106 482 108
rect 510 106 512 108
rect 540 106 542 108
rect 60 100 62 102
rect 90 100 92 102
rect 120 100 122 102
rect 150 100 152 102
rect 180 100 182 102
rect 210 100 212 102
rect 240 100 242 102
rect 270 100 272 102
rect 300 100 302 102
rect 330 100 332 102
rect 360 100 362 102
rect 390 100 392 102
rect 420 100 422 102
rect 450 100 452 102
rect 480 100 482 102
rect 510 100 512 102
rect 540 100 542 102
rect 62 98 64 100
rect 68 98 70 100
rect 92 98 94 100
rect 98 98 100 100
rect 122 98 124 100
rect 128 98 130 100
rect 152 98 154 100
rect 158 98 160 100
rect 182 98 184 100
rect 188 98 190 100
rect 212 98 214 100
rect 218 98 220 100
rect 242 98 244 100
rect 248 98 250 100
rect 272 98 274 100
rect 278 98 280 100
rect 302 98 304 100
rect 308 98 310 100
rect 332 98 334 100
rect 338 98 340 100
rect 362 98 364 100
rect 368 98 370 100
rect 392 98 394 100
rect 398 98 400 100
rect 422 98 424 100
rect 428 98 430 100
rect 452 98 454 100
rect 458 98 460 100
rect 482 98 484 100
rect 488 98 490 100
rect 512 98 514 100
rect 518 98 520 100
rect 542 98 544 100
rect 548 98 550 100
rect 70 96 72 98
rect 100 96 102 98
rect 130 96 132 98
rect 160 96 162 98
rect 190 96 192 98
rect 220 96 222 98
rect 250 96 252 98
rect 280 96 282 98
rect 310 96 312 98
rect 340 96 342 98
rect 370 96 372 98
rect 400 96 402 98
rect 430 96 432 98
rect 460 96 462 98
rect 490 96 492 98
rect 520 96 522 98
rect 550 96 552 98
rect 70 90 72 92
rect 100 90 102 92
rect 130 90 132 92
rect 160 90 162 92
rect 190 90 192 92
rect 220 90 222 92
rect 250 90 252 92
rect 280 90 282 92
rect 310 90 312 92
rect 340 90 342 92
rect 370 90 372 92
rect 400 90 402 92
rect 430 90 432 92
rect 460 90 462 92
rect 490 90 492 92
rect 520 90 522 92
rect 550 90 552 92
rect 62 88 64 90
rect 68 88 70 90
rect 92 88 94 90
rect 98 88 100 90
rect 122 88 124 90
rect 128 88 130 90
rect 152 88 154 90
rect 158 88 160 90
rect 182 88 184 90
rect 188 88 190 90
rect 212 88 214 90
rect 218 88 220 90
rect 242 88 244 90
rect 248 88 250 90
rect 272 88 274 90
rect 278 88 280 90
rect 302 88 304 90
rect 308 88 310 90
rect 332 88 334 90
rect 338 88 340 90
rect 362 88 364 90
rect 368 88 370 90
rect 392 88 394 90
rect 398 88 400 90
rect 422 88 424 90
rect 428 88 430 90
rect 452 88 454 90
rect 458 88 460 90
rect 482 88 484 90
rect 488 88 490 90
rect 512 88 514 90
rect 518 88 520 90
rect 542 88 544 90
rect 548 88 550 90
rect 60 86 62 88
rect 90 86 92 88
rect 120 86 122 88
rect 150 86 152 88
rect 180 86 182 88
rect 210 86 212 88
rect 240 86 242 88
rect 270 86 272 88
rect 300 86 302 88
rect 330 86 332 88
rect 360 86 362 88
rect 390 86 392 88
rect 420 86 422 88
rect 450 86 452 88
rect 480 86 482 88
rect 510 86 512 88
rect 540 86 542 88
rect 60 80 62 82
rect 90 80 92 82
rect 120 80 122 82
rect 150 80 152 82
rect 180 80 182 82
rect 210 80 212 82
rect 240 80 242 82
rect 270 80 272 82
rect 300 80 302 82
rect 330 80 332 82
rect 360 80 362 82
rect 390 80 392 82
rect 420 80 422 82
rect 450 80 452 82
rect 480 80 482 82
rect 510 80 512 82
rect 540 80 542 82
rect 62 78 64 80
rect 68 78 70 80
rect 92 78 94 80
rect 98 78 100 80
rect 122 78 124 80
rect 128 78 130 80
rect 152 78 154 80
rect 158 78 160 80
rect 182 78 184 80
rect 188 78 190 80
rect 212 78 214 80
rect 218 78 220 80
rect 242 78 244 80
rect 248 78 250 80
rect 272 78 274 80
rect 278 78 280 80
rect 302 78 304 80
rect 308 78 310 80
rect 332 78 334 80
rect 338 78 340 80
rect 362 78 364 80
rect 368 78 370 80
rect 392 78 394 80
rect 398 78 400 80
rect 422 78 424 80
rect 428 78 430 80
rect 452 78 454 80
rect 458 78 460 80
rect 482 78 484 80
rect 488 78 490 80
rect 512 78 514 80
rect 518 78 520 80
rect 542 78 544 80
rect 548 78 550 80
rect 70 76 72 78
rect 100 76 102 78
rect 130 76 132 78
rect 160 76 162 78
rect 190 76 192 78
rect 220 76 222 78
rect 250 76 252 78
rect 280 76 282 78
rect 310 76 312 78
rect 340 76 342 78
rect 370 76 372 78
rect 400 76 402 78
rect 430 76 432 78
rect 460 76 462 78
rect 490 76 492 78
rect 520 76 522 78
rect 550 76 552 78
rect 70 70 72 72
rect 100 70 102 72
rect 130 70 132 72
rect 160 70 162 72
rect 190 70 192 72
rect 220 70 222 72
rect 250 70 252 72
rect 280 70 282 72
rect 310 70 312 72
rect 340 70 342 72
rect 370 70 372 72
rect 400 70 402 72
rect 430 70 432 72
rect 460 70 462 72
rect 490 70 492 72
rect 520 70 522 72
rect 550 70 552 72
rect 62 68 64 70
rect 68 68 70 70
rect 92 68 94 70
rect 98 68 100 70
rect 122 68 124 70
rect 128 68 130 70
rect 152 68 154 70
rect 158 68 160 70
rect 182 68 184 70
rect 188 68 190 70
rect 212 68 214 70
rect 218 68 220 70
rect 242 68 244 70
rect 248 68 250 70
rect 272 68 274 70
rect 278 68 280 70
rect 302 68 304 70
rect 308 68 310 70
rect 332 68 334 70
rect 338 68 340 70
rect 362 68 364 70
rect 368 68 370 70
rect 392 68 394 70
rect 398 68 400 70
rect 422 68 424 70
rect 428 68 430 70
rect 452 68 454 70
rect 458 68 460 70
rect 482 68 484 70
rect 488 68 490 70
rect 512 68 514 70
rect 518 68 520 70
rect 542 68 544 70
rect 548 68 550 70
rect 60 66 62 68
rect 90 66 92 68
rect 120 66 122 68
rect 150 66 152 68
rect 180 66 182 68
rect 210 66 212 68
rect 240 66 242 68
rect 270 66 272 68
rect 300 66 302 68
rect 330 66 332 68
rect 360 66 362 68
rect 390 66 392 68
rect 420 66 422 68
rect 450 66 452 68
rect 480 66 482 68
rect 510 66 512 68
rect 540 66 542 68
rect 60 60 62 62
rect 90 60 92 62
rect 120 60 122 62
rect 150 60 152 62
rect 180 60 182 62
rect 210 60 212 62
rect 240 60 242 62
rect 270 60 272 62
rect 300 60 302 62
rect 330 60 332 62
rect 360 60 362 62
rect 390 60 392 62
rect 420 60 422 62
rect 450 60 452 62
rect 480 60 482 62
rect 510 60 512 62
rect 540 60 542 62
rect 62 58 64 60
rect 68 58 70 60
rect 92 58 94 60
rect 98 58 100 60
rect 122 58 124 60
rect 128 58 130 60
rect 152 58 154 60
rect 158 58 160 60
rect 182 58 184 60
rect 188 58 190 60
rect 212 58 214 60
rect 218 58 220 60
rect 242 58 244 60
rect 248 58 250 60
rect 272 58 274 60
rect 278 58 280 60
rect 302 58 304 60
rect 308 58 310 60
rect 332 58 334 60
rect 338 58 340 60
rect 362 58 364 60
rect 368 58 370 60
rect 392 58 394 60
rect 398 58 400 60
rect 422 58 424 60
rect 428 58 430 60
rect 452 58 454 60
rect 458 58 460 60
rect 482 58 484 60
rect 488 58 490 60
rect 512 58 514 60
rect 518 58 520 60
rect 542 58 544 60
rect 548 58 550 60
rect 70 56 72 58
rect 100 56 102 58
rect 130 56 132 58
rect 160 56 162 58
rect 190 56 192 58
rect 220 56 222 58
rect 250 56 252 58
rect 280 56 282 58
rect 310 56 312 58
rect 340 56 342 58
rect 370 56 372 58
rect 400 56 402 58
rect 430 56 432 58
rect 460 56 462 58
rect 490 56 492 58
rect 520 56 522 58
rect 550 56 552 58
rect 70 50 72 52
rect 100 50 102 52
rect 130 50 132 52
rect 160 50 162 52
rect 190 50 192 52
rect 220 50 222 52
rect 250 50 252 52
rect 280 50 282 52
rect 310 50 312 52
rect 340 50 342 52
rect 370 50 372 52
rect 400 50 402 52
rect 430 50 432 52
rect 460 50 462 52
rect 490 50 492 52
rect 520 50 522 52
rect 550 50 552 52
rect 62 48 64 50
rect 68 48 70 50
rect 92 48 94 50
rect 98 48 100 50
rect 122 48 124 50
rect 128 48 130 50
rect 152 48 154 50
rect 158 48 160 50
rect 182 48 184 50
rect 188 48 190 50
rect 212 48 214 50
rect 218 48 220 50
rect 242 48 244 50
rect 248 48 250 50
rect 272 48 274 50
rect 278 48 280 50
rect 302 48 304 50
rect 308 48 310 50
rect 332 48 334 50
rect 338 48 340 50
rect 362 48 364 50
rect 368 48 370 50
rect 392 48 394 50
rect 398 48 400 50
rect 422 48 424 50
rect 428 48 430 50
rect 452 48 454 50
rect 458 48 460 50
rect 482 48 484 50
rect 488 48 490 50
rect 512 48 514 50
rect 518 48 520 50
rect 542 48 544 50
rect 548 48 550 50
rect 60 46 62 48
rect 90 46 92 48
rect 120 46 122 48
rect 150 46 152 48
rect 180 46 182 48
rect 210 46 212 48
rect 240 46 242 48
rect 270 46 272 48
rect 300 46 302 48
rect 330 46 332 48
rect 360 46 362 48
rect 390 46 392 48
rect 420 46 422 48
rect 450 46 452 48
rect 480 46 482 48
rect 510 46 512 48
rect 540 46 542 48
rect 60 40 62 42
rect 90 40 92 42
rect 120 40 122 42
rect 150 40 152 42
rect 180 40 182 42
rect 210 40 212 42
rect 240 40 242 42
rect 270 40 272 42
rect 300 40 302 42
rect 330 40 332 42
rect 360 40 362 42
rect 390 40 392 42
rect 420 40 422 42
rect 450 40 452 42
rect 480 40 482 42
rect 510 40 512 42
rect 540 40 542 42
rect 62 38 64 40
rect 68 38 70 40
rect 92 38 94 40
rect 98 38 100 40
rect 122 38 124 40
rect 128 38 130 40
rect 152 38 154 40
rect 158 38 160 40
rect 182 38 184 40
rect 188 38 190 40
rect 212 38 214 40
rect 218 38 220 40
rect 242 38 244 40
rect 248 38 250 40
rect 272 38 274 40
rect 278 38 280 40
rect 302 38 304 40
rect 308 38 310 40
rect 332 38 334 40
rect 338 38 340 40
rect 362 38 364 40
rect 368 38 370 40
rect 392 38 394 40
rect 398 38 400 40
rect 422 38 424 40
rect 428 38 430 40
rect 452 38 454 40
rect 458 38 460 40
rect 482 38 484 40
rect 488 38 490 40
rect 512 38 514 40
rect 518 38 520 40
rect 542 38 544 40
rect 548 38 550 40
rect 70 36 72 38
rect 100 36 102 38
rect 130 36 132 38
rect 160 36 162 38
rect 190 36 192 38
rect 220 36 222 38
rect 250 36 252 38
rect 280 36 282 38
rect 310 36 312 38
rect 340 36 342 38
rect 370 36 372 38
rect 400 36 402 38
rect 430 36 432 38
rect 460 36 462 38
rect 490 36 492 38
rect 520 36 522 38
rect 550 36 552 38
<< nwell >>
rect 34 858 566 1306
rect -6 498 606 660
rect -6 22 22 498
rect 578 22 606 498
rect -6 -6 606 22
<< psubstratepdiff >>
rect 0 1336 600 1340
rect 0 828 4 1336
rect 332 1328 338 1336
rect 12 1318 588 1328
rect 12 846 22 1318
rect 578 846 588 1318
rect 12 836 588 846
rect 12 828 24 836
rect 42 828 54 836
rect 72 828 84 836
rect 102 828 114 836
rect 132 828 144 836
rect 162 828 174 836
rect 192 828 204 836
rect 222 828 234 836
rect 242 828 256 836
rect 264 828 276 836
rect 294 828 306 836
rect 324 828 336 836
rect 344 828 358 836
rect 366 828 378 836
rect 396 828 408 836
rect 426 828 438 836
rect 456 828 468 836
rect 486 828 498 836
rect 516 828 528 836
rect 546 828 558 836
rect 576 828 588 836
rect 596 828 600 1336
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 184 828
rect 192 826 214 828
rect 222 826 286 828
rect 294 826 316 828
rect 324 826 378 828
rect 386 826 408 828
rect 416 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 0 818 14 826
rect 22 818 34 826
rect 52 818 64 826
rect 82 818 94 826
rect 112 818 124 826
rect 142 818 154 826
rect 172 818 184 826
rect 202 818 214 826
rect 232 818 244 826
rect 252 818 266 826
rect 274 818 286 826
rect 304 818 316 826
rect 334 818 348 826
rect 356 818 368 826
rect 386 818 398 826
rect 416 818 428 826
rect 446 818 458 826
rect 476 818 488 826
rect 506 818 518 826
rect 536 818 548 826
rect 566 818 578 826
rect 586 818 600 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 184 818
rect 192 816 214 818
rect 222 816 286 818
rect 294 816 316 818
rect 324 816 378 818
rect 386 816 408 818
rect 416 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 0 808 4 816
rect 12 808 24 816
rect 42 808 54 816
rect 72 808 84 816
rect 102 808 114 816
rect 132 808 144 816
rect 162 808 174 816
rect 192 808 204 816
rect 222 808 234 816
rect 242 808 256 816
rect 264 808 276 816
rect 294 808 306 816
rect 324 808 336 816
rect 344 808 358 816
rect 366 808 378 816
rect 396 808 408 816
rect 426 808 438 816
rect 456 808 468 816
rect 486 808 498 816
rect 516 808 528 816
rect 546 808 558 816
rect 576 808 588 816
rect 596 808 600 816
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 184 808
rect 192 806 214 808
rect 222 806 286 808
rect 294 806 316 808
rect 324 806 378 808
rect 386 806 408 808
rect 416 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 0 798 14 806
rect 22 798 34 806
rect 52 798 64 806
rect 82 798 94 806
rect 112 798 124 806
rect 142 798 154 806
rect 172 798 184 806
rect 202 798 214 806
rect 232 798 244 806
rect 252 798 266 806
rect 274 798 286 806
rect 304 798 316 806
rect 334 798 348 806
rect 356 798 368 806
rect 386 798 398 806
rect 416 798 428 806
rect 446 798 458 806
rect 476 798 488 806
rect 506 798 518 806
rect 536 798 548 806
rect 566 798 578 806
rect 586 798 600 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 184 798
rect 192 796 214 798
rect 222 796 286 798
rect 294 796 316 798
rect 324 796 378 798
rect 386 796 408 798
rect 416 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 0 788 4 796
rect 12 788 24 796
rect 42 788 54 796
rect 72 788 84 796
rect 102 788 114 796
rect 132 788 144 796
rect 162 788 174 796
rect 192 788 204 796
rect 222 788 234 796
rect 242 788 256 796
rect 264 788 276 796
rect 294 788 306 796
rect 324 788 336 796
rect 344 788 358 796
rect 366 788 378 796
rect 396 788 408 796
rect 426 788 438 796
rect 456 788 468 796
rect 486 788 498 796
rect 516 788 528 796
rect 546 788 558 796
rect 576 788 588 796
rect 596 788 600 796
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 184 788
rect 192 786 214 788
rect 222 786 286 788
rect 294 786 316 788
rect 324 786 378 788
rect 386 786 408 788
rect 416 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 0 778 14 786
rect 22 778 34 786
rect 52 778 64 786
rect 82 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 776 124 786
rect 142 776 154 786
rect 172 776 184 786
rect 202 776 214 786
rect 232 776 244 786
rect 252 776 266 786
rect 274 776 286 786
rect 304 776 316 786
rect 334 776 348 786
rect 356 776 368 786
rect 386 776 398 786
rect 416 776 428 786
rect 446 776 458 786
rect 476 776 488 786
rect 506 778 518 786
rect 536 778 548 786
rect 566 778 578 786
rect 586 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 0 768 4 776
rect 12 768 24 776
rect 42 768 54 776
rect 72 768 84 776
rect 252 768 256 776
rect 344 768 348 776
rect 516 768 528 776
rect 546 768 558 776
rect 576 768 588 776
rect 596 768 600 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 14 766
rect 22 758 34 766
rect 52 758 64 766
rect 82 758 94 766
rect 112 758 124 768
rect 142 758 154 768
rect 172 758 184 768
rect 202 758 214 768
rect 232 758 244 768
rect 252 758 266 768
rect 274 758 286 768
rect 304 758 316 768
rect 334 758 348 768
rect 356 758 368 768
rect 386 758 398 768
rect 416 758 428 768
rect 446 758 458 768
rect 476 758 488 768
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 518 766
rect 536 758 548 766
rect 566 758 578 766
rect 586 758 600 766
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 184 758
rect 192 756 214 758
rect 222 756 286 758
rect 294 756 316 758
rect 324 756 378 758
rect 386 756 408 758
rect 416 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 0 748 4 756
rect 12 748 24 756
rect 42 748 54 756
rect 72 748 84 756
rect 102 748 114 756
rect 132 748 144 756
rect 162 748 174 756
rect 192 748 204 756
rect 222 748 234 756
rect 242 748 256 756
rect 264 748 276 756
rect 294 748 306 756
rect 324 748 336 756
rect 344 748 358 756
rect 366 748 378 756
rect 396 748 408 756
rect 426 748 438 756
rect 456 748 468 756
rect 486 748 498 756
rect 516 748 528 756
rect 546 748 558 756
rect 576 748 588 756
rect 596 748 600 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 184 748
rect 192 746 214 748
rect 222 746 286 748
rect 294 746 316 748
rect 324 746 378 748
rect 386 746 408 748
rect 416 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 0 738 14 746
rect 22 738 34 746
rect 52 738 64 746
rect 82 738 94 746
rect 112 738 124 746
rect 142 738 154 746
rect 172 738 184 746
rect 202 738 214 746
rect 232 738 244 746
rect 252 738 266 746
rect 274 738 286 746
rect 304 738 316 746
rect 334 738 348 746
rect 356 738 368 746
rect 386 738 398 746
rect 416 738 428 746
rect 446 738 458 746
rect 476 738 488 746
rect 506 738 518 746
rect 536 738 548 746
rect 566 738 578 746
rect 586 738 600 746
rect 0 736 214 738
rect 0 728 4 736
rect 12 728 24 736
rect 32 728 214 736
rect 0 726 214 728
rect 222 736 286 738
rect 294 736 316 738
rect 324 736 378 738
rect 222 728 234 736
rect 242 728 256 736
rect 264 728 276 736
rect 294 728 306 736
rect 324 728 336 736
rect 344 728 358 736
rect 366 728 378 736
rect 222 726 286 728
rect 294 726 316 728
rect 324 726 378 728
rect 386 736 600 738
rect 386 728 568 736
rect 576 728 588 736
rect 596 728 600 736
rect 386 726 600 728
rect 0 718 14 726
rect 22 718 34 726
rect 52 718 64 726
rect 82 718 94 726
rect 112 718 124 726
rect 142 718 154 726
rect 172 718 184 726
rect 202 718 214 726
rect 232 718 244 726
rect 252 718 266 726
rect 274 718 286 726
rect 304 718 316 726
rect 334 718 348 726
rect 356 718 368 726
rect 386 718 398 726
rect 416 718 428 726
rect 446 718 458 726
rect 476 718 488 726
rect 506 718 518 726
rect 536 718 548 726
rect 566 718 578 726
rect 586 718 600 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 184 718
rect 192 716 214 718
rect 222 716 286 718
rect 294 716 316 718
rect 324 716 378 718
rect 386 716 408 718
rect 416 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 0 708 4 716
rect 12 708 24 716
rect 42 708 54 716
rect 72 708 84 716
rect 102 708 114 716
rect 132 708 144 716
rect 162 708 174 716
rect 192 708 204 716
rect 222 708 234 716
rect 242 708 256 716
rect 264 708 276 716
rect 294 708 306 716
rect 324 708 336 716
rect 344 708 358 716
rect 366 708 378 716
rect 396 708 408 716
rect 426 708 438 716
rect 456 708 468 716
rect 486 708 498 716
rect 516 708 528 716
rect 546 708 558 716
rect 576 708 588 716
rect 596 708 600 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 184 708
rect 192 706 214 708
rect 222 706 286 708
rect 294 706 316 708
rect 324 706 378 708
rect 386 706 408 708
rect 416 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 0 698 14 706
rect 22 698 34 706
rect 52 698 64 706
rect 82 698 94 706
rect 112 698 124 706
rect 142 698 154 706
rect 172 698 184 706
rect 202 698 214 706
rect 232 698 244 706
rect 252 698 266 706
rect 274 698 286 706
rect 304 698 316 706
rect 334 698 348 706
rect 356 698 368 706
rect 386 698 398 706
rect 416 698 428 706
rect 446 698 458 706
rect 476 698 488 706
rect 506 698 518 706
rect 536 698 548 706
rect 566 698 578 706
rect 586 698 600 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 184 698
rect 192 696 214 698
rect 222 696 286 698
rect 294 696 316 698
rect 324 696 378 698
rect 386 696 408 698
rect 416 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 0 688 4 696
rect 12 688 24 696
rect 42 688 54 696
rect 72 688 84 696
rect 102 688 114 696
rect 132 688 144 696
rect 162 688 174 696
rect 192 688 204 696
rect 222 688 234 696
rect 242 688 256 696
rect 264 688 276 696
rect 294 688 306 696
rect 324 688 336 696
rect 344 688 358 696
rect 366 688 378 696
rect 396 688 408 696
rect 426 688 438 696
rect 456 688 468 696
rect 486 688 498 696
rect 516 688 528 696
rect 546 688 558 696
rect 576 688 588 696
rect 596 688 600 696
rect 0 686 600 688
rect 28 488 572 492
rect 28 460 32 488
rect 570 460 572 488
rect 28 450 42 460
rect 50 450 62 460
rect 80 450 92 460
rect 110 450 122 460
rect 140 450 152 460
rect 170 450 182 460
rect 200 450 212 460
rect 230 450 242 460
rect 260 450 272 460
rect 290 450 302 460
rect 320 450 332 460
rect 350 450 362 460
rect 380 450 392 460
rect 410 450 422 460
rect 440 450 452 460
rect 470 450 482 460
rect 500 450 512 460
rect 530 450 542 460
rect 560 450 572 460
rect 28 448 62 450
rect 70 448 92 450
rect 100 448 122 450
rect 130 448 152 450
rect 160 448 182 450
rect 190 448 212 450
rect 220 448 242 450
rect 250 448 272 450
rect 280 448 302 450
rect 310 448 332 450
rect 340 448 362 450
rect 370 448 392 450
rect 400 448 422 450
rect 430 448 452 450
rect 460 448 482 450
rect 490 448 512 450
rect 520 448 542 450
rect 550 448 572 450
rect 28 440 32 448
rect 40 440 52 448
rect 70 440 82 448
rect 100 440 112 448
rect 130 440 142 448
rect 160 440 172 448
rect 190 440 202 448
rect 220 440 232 448
rect 250 440 262 448
rect 280 440 292 448
rect 310 440 322 448
rect 340 440 352 448
rect 370 440 382 448
rect 400 440 412 448
rect 430 440 442 448
rect 460 440 472 448
rect 490 440 502 448
rect 520 440 532 448
rect 550 440 562 448
rect 570 440 572 448
rect 28 438 62 440
rect 70 438 92 440
rect 100 438 122 440
rect 130 438 152 440
rect 160 438 182 440
rect 190 438 212 440
rect 220 438 242 440
rect 250 438 272 440
rect 280 438 302 440
rect 310 438 332 440
rect 340 438 362 440
rect 370 438 392 440
rect 400 438 422 440
rect 430 438 452 440
rect 460 438 482 440
rect 490 438 512 440
rect 520 438 542 440
rect 550 438 572 440
rect 28 430 42 438
rect 50 430 62 438
rect 80 430 92 438
rect 110 430 122 438
rect 140 430 152 438
rect 170 430 182 438
rect 200 430 212 438
rect 230 430 242 438
rect 260 430 272 438
rect 290 430 302 438
rect 320 430 332 438
rect 350 430 362 438
rect 380 430 392 438
rect 410 430 422 438
rect 440 430 452 438
rect 470 430 482 438
rect 500 430 512 438
rect 530 430 542 438
rect 560 430 572 438
rect 28 428 62 430
rect 70 428 92 430
rect 100 428 122 430
rect 130 428 152 430
rect 160 428 182 430
rect 190 428 212 430
rect 220 428 242 430
rect 250 428 272 430
rect 280 428 302 430
rect 310 428 332 430
rect 340 428 362 430
rect 370 428 392 430
rect 400 428 422 430
rect 430 428 452 430
rect 460 428 482 430
rect 490 428 512 430
rect 520 428 542 430
rect 550 428 572 430
rect 28 420 32 428
rect 40 420 52 428
rect 70 420 82 428
rect 100 420 112 428
rect 130 420 142 428
rect 160 420 172 428
rect 190 420 202 428
rect 220 420 232 428
rect 250 420 262 428
rect 280 420 292 428
rect 310 420 322 428
rect 340 420 352 428
rect 370 420 382 428
rect 400 420 412 428
rect 430 420 442 428
rect 460 420 472 428
rect 490 420 502 428
rect 520 420 532 428
rect 550 420 562 428
rect 570 420 572 428
rect 28 418 62 420
rect 70 418 92 420
rect 100 418 122 420
rect 130 418 152 420
rect 160 418 182 420
rect 190 418 212 420
rect 220 418 242 420
rect 250 418 272 420
rect 280 418 302 420
rect 310 418 332 420
rect 340 418 362 420
rect 370 418 392 420
rect 400 418 422 420
rect 430 418 452 420
rect 460 418 482 420
rect 490 418 512 420
rect 520 418 542 420
rect 550 418 572 420
rect 28 410 42 418
rect 50 410 62 418
rect 80 410 92 418
rect 110 410 122 418
rect 140 410 152 418
rect 170 410 182 418
rect 200 410 212 418
rect 230 410 242 418
rect 260 410 272 418
rect 290 410 302 418
rect 320 410 332 418
rect 350 410 362 418
rect 380 410 392 418
rect 410 410 422 418
rect 440 410 452 418
rect 470 410 482 418
rect 500 410 512 418
rect 530 410 542 418
rect 560 410 572 418
rect 28 408 62 410
rect 70 408 92 410
rect 100 408 122 410
rect 130 408 152 410
rect 160 408 182 410
rect 190 408 212 410
rect 220 408 242 410
rect 250 408 272 410
rect 280 408 302 410
rect 310 408 332 410
rect 340 408 362 410
rect 370 408 392 410
rect 400 408 422 410
rect 430 408 452 410
rect 460 408 482 410
rect 490 408 512 410
rect 520 408 542 410
rect 550 408 572 410
rect 28 400 32 408
rect 40 400 52 408
rect 70 400 82 408
rect 100 400 112 408
rect 130 400 142 408
rect 160 400 172 408
rect 190 400 202 408
rect 220 400 232 408
rect 250 400 262 408
rect 280 400 292 408
rect 310 400 322 408
rect 340 400 352 408
rect 370 400 382 408
rect 400 400 412 408
rect 430 400 442 408
rect 460 400 472 408
rect 490 400 502 408
rect 520 400 532 408
rect 550 400 562 408
rect 570 400 572 408
rect 28 398 62 400
rect 70 398 92 400
rect 100 398 122 400
rect 130 398 152 400
rect 160 398 182 400
rect 190 398 212 400
rect 220 398 242 400
rect 250 398 272 400
rect 280 398 302 400
rect 310 398 332 400
rect 340 398 362 400
rect 370 398 392 400
rect 400 398 422 400
rect 430 398 452 400
rect 460 398 482 400
rect 490 398 512 400
rect 520 398 542 400
rect 550 398 572 400
rect 28 370 42 398
rect 50 370 62 398
rect 80 370 92 398
rect 110 390 122 398
rect 140 390 152 398
rect 170 390 182 398
rect 200 390 212 398
rect 230 390 242 398
rect 260 390 272 398
rect 290 390 302 398
rect 320 390 332 398
rect 350 390 362 398
rect 380 390 392 398
rect 410 390 422 398
rect 440 390 452 398
rect 470 390 482 398
rect 500 390 512 398
rect 530 390 542 398
rect 560 390 572 398
rect 100 378 512 390
rect 520 388 542 390
rect 550 388 572 390
rect 520 380 532 388
rect 550 380 562 388
rect 570 380 572 388
rect 520 378 542 380
rect 550 378 572 380
rect 110 370 122 378
rect 140 370 152 378
rect 170 370 182 378
rect 200 370 212 378
rect 230 370 242 378
rect 260 370 272 378
rect 290 370 302 378
rect 320 370 332 378
rect 350 370 362 378
rect 380 370 392 378
rect 410 370 422 378
rect 440 370 452 378
rect 470 370 482 378
rect 500 370 512 378
rect 530 370 542 378
rect 560 370 572 378
rect 28 368 62 370
rect 70 368 92 370
rect 100 368 122 370
rect 130 368 152 370
rect 160 368 182 370
rect 190 368 212 370
rect 220 368 242 370
rect 250 368 272 370
rect 280 368 302 370
rect 310 368 332 370
rect 340 368 362 370
rect 370 368 392 370
rect 400 368 422 370
rect 430 368 452 370
rect 460 368 482 370
rect 490 368 512 370
rect 520 368 542 370
rect 550 368 572 370
rect 28 360 32 368
rect 40 360 52 368
rect 70 360 82 368
rect 100 360 112 368
rect 130 360 142 368
rect 160 360 172 368
rect 190 360 202 368
rect 220 360 232 368
rect 250 360 262 368
rect 280 360 292 368
rect 310 360 322 368
rect 340 360 352 368
rect 370 360 382 368
rect 400 360 412 368
rect 430 360 442 368
rect 460 360 472 368
rect 490 360 502 368
rect 520 360 532 368
rect 550 360 562 368
rect 570 360 572 368
rect 28 358 62 360
rect 70 358 92 360
rect 100 358 122 360
rect 130 358 152 360
rect 160 358 182 360
rect 190 358 212 360
rect 220 358 242 360
rect 250 358 272 360
rect 280 358 302 360
rect 310 358 332 360
rect 340 358 362 360
rect 370 358 392 360
rect 400 358 422 360
rect 430 358 452 360
rect 460 358 482 360
rect 490 358 512 360
rect 520 358 542 360
rect 550 358 572 360
rect 28 350 42 358
rect 50 350 62 358
rect 80 350 92 358
rect 110 350 122 358
rect 140 350 152 358
rect 170 350 182 358
rect 200 350 212 358
rect 230 350 242 358
rect 260 350 272 358
rect 290 350 302 358
rect 320 350 332 358
rect 350 350 362 358
rect 380 350 392 358
rect 410 350 422 358
rect 440 350 452 358
rect 470 350 482 358
rect 500 350 512 358
rect 530 350 542 358
rect 560 350 572 358
rect 28 348 62 350
rect 70 348 92 350
rect 100 348 122 350
rect 130 348 152 350
rect 160 348 182 350
rect 190 348 212 350
rect 220 348 242 350
rect 250 348 272 350
rect 280 348 302 350
rect 310 348 332 350
rect 340 348 362 350
rect 370 348 392 350
rect 400 348 422 350
rect 430 348 452 350
rect 460 348 482 350
rect 490 348 512 350
rect 520 348 542 350
rect 550 348 572 350
rect 28 340 32 348
rect 40 340 52 348
rect 70 340 82 348
rect 100 340 112 348
rect 130 340 142 348
rect 160 340 172 348
rect 190 340 202 348
rect 220 340 232 348
rect 250 340 262 348
rect 280 340 292 348
rect 310 340 322 348
rect 340 340 352 348
rect 370 340 382 348
rect 400 340 412 348
rect 430 340 442 348
rect 460 340 472 348
rect 490 340 502 348
rect 520 340 532 348
rect 550 340 562 348
rect 570 340 572 348
rect 28 338 62 340
rect 70 338 92 340
rect 100 338 122 340
rect 130 338 152 340
rect 160 338 182 340
rect 190 338 212 340
rect 220 338 242 340
rect 250 338 272 340
rect 280 338 302 340
rect 310 338 332 340
rect 340 338 362 340
rect 370 338 392 340
rect 400 338 422 340
rect 430 338 452 340
rect 460 338 482 340
rect 490 338 512 340
rect 520 338 542 340
rect 550 338 572 340
rect 28 330 42 338
rect 50 330 62 338
rect 80 330 92 338
rect 110 330 122 338
rect 140 330 152 338
rect 170 330 182 338
rect 200 330 212 338
rect 230 330 242 338
rect 260 330 272 338
rect 290 330 302 338
rect 320 330 332 338
rect 350 330 362 338
rect 380 330 392 338
rect 410 330 422 338
rect 440 330 452 338
rect 470 330 482 338
rect 500 330 512 338
rect 530 330 542 338
rect 560 330 572 338
rect 28 328 62 330
rect 70 328 92 330
rect 100 328 122 330
rect 130 328 152 330
rect 160 328 182 330
rect 190 328 212 330
rect 220 328 242 330
rect 250 328 272 330
rect 280 328 302 330
rect 310 328 332 330
rect 340 328 362 330
rect 370 328 392 330
rect 400 328 422 330
rect 430 328 452 330
rect 460 328 482 330
rect 490 328 512 330
rect 520 328 542 330
rect 550 328 572 330
rect 28 320 32 328
rect 40 320 52 328
rect 70 320 82 328
rect 100 320 112 328
rect 130 320 142 328
rect 160 320 172 328
rect 190 320 202 328
rect 220 320 232 328
rect 250 320 262 328
rect 280 320 292 328
rect 310 320 322 328
rect 340 320 352 328
rect 370 320 382 328
rect 400 320 412 328
rect 430 320 442 328
rect 460 320 472 328
rect 490 320 502 328
rect 520 320 532 328
rect 550 320 562 328
rect 570 320 572 328
rect 28 318 62 320
rect 70 318 92 320
rect 100 318 122 320
rect 130 318 152 320
rect 160 318 182 320
rect 190 318 212 320
rect 220 318 242 320
rect 250 318 272 320
rect 280 318 302 320
rect 310 318 332 320
rect 340 318 362 320
rect 370 318 392 320
rect 400 318 422 320
rect 430 318 452 320
rect 460 318 482 320
rect 490 318 512 320
rect 520 318 542 320
rect 550 318 572 320
rect 28 310 42 318
rect 50 310 62 318
rect 80 310 92 318
rect 110 310 122 318
rect 140 310 152 318
rect 170 310 182 318
rect 200 310 212 318
rect 230 310 242 318
rect 260 310 272 318
rect 290 310 302 318
rect 320 310 332 318
rect 350 310 362 318
rect 380 310 392 318
rect 410 310 422 318
rect 440 310 452 318
rect 470 310 482 318
rect 500 310 512 318
rect 530 310 542 318
rect 560 310 572 318
rect 28 308 62 310
rect 70 308 512 310
rect 520 308 542 310
rect 550 308 572 310
rect 28 300 32 308
rect 40 300 52 308
rect 70 300 82 308
rect 90 300 502 308
rect 520 300 532 308
rect 550 300 562 308
rect 570 300 572 308
rect 28 298 62 300
rect 70 298 512 300
rect 520 298 542 300
rect 550 298 572 300
rect 28 290 42 298
rect 50 290 62 298
rect 80 290 92 298
rect 110 290 122 298
rect 140 290 152 298
rect 170 290 182 298
rect 200 290 212 298
rect 230 290 242 298
rect 260 290 272 298
rect 290 290 302 298
rect 320 290 332 298
rect 350 290 362 298
rect 380 290 392 298
rect 410 290 422 298
rect 440 290 452 298
rect 470 290 482 298
rect 500 290 512 298
rect 530 290 542 298
rect 560 290 572 298
rect 28 288 62 290
rect 70 288 92 290
rect 100 288 122 290
rect 130 288 152 290
rect 160 288 182 290
rect 190 288 212 290
rect 220 288 242 290
rect 250 288 272 290
rect 280 288 302 290
rect 310 288 332 290
rect 340 288 362 290
rect 370 288 392 290
rect 400 288 422 290
rect 430 288 452 290
rect 460 288 482 290
rect 490 288 512 290
rect 520 288 542 290
rect 550 288 572 290
rect 28 280 32 288
rect 40 280 52 288
rect 70 280 82 288
rect 100 280 112 288
rect 130 280 142 288
rect 160 280 172 288
rect 190 280 202 288
rect 220 280 232 288
rect 250 280 262 288
rect 280 280 292 288
rect 310 280 322 288
rect 340 280 352 288
rect 370 280 382 288
rect 400 280 412 288
rect 430 280 442 288
rect 460 280 472 288
rect 490 280 502 288
rect 520 280 532 288
rect 550 280 562 288
rect 570 280 572 288
rect 28 278 62 280
rect 70 278 92 280
rect 100 278 122 280
rect 130 278 152 280
rect 160 278 182 280
rect 190 278 212 280
rect 220 278 242 280
rect 250 278 272 280
rect 280 278 302 280
rect 310 278 332 280
rect 340 278 362 280
rect 370 278 392 280
rect 400 278 422 280
rect 430 278 452 280
rect 460 278 482 280
rect 490 278 512 280
rect 520 278 542 280
rect 550 278 572 280
rect 28 270 42 278
rect 50 270 62 278
rect 80 270 92 278
rect 110 270 122 278
rect 140 270 152 278
rect 170 270 182 278
rect 200 270 212 278
rect 230 270 242 278
rect 260 270 272 278
rect 290 270 302 278
rect 320 270 332 278
rect 350 270 362 278
rect 380 270 392 278
rect 410 270 422 278
rect 440 270 452 278
rect 470 270 482 278
rect 500 270 512 278
rect 530 270 542 278
rect 560 270 572 278
rect 28 268 62 270
rect 70 268 92 270
rect 100 268 122 270
rect 130 268 152 270
rect 160 268 182 270
rect 190 268 212 270
rect 220 268 242 270
rect 250 268 272 270
rect 280 268 302 270
rect 310 268 332 270
rect 340 268 362 270
rect 370 268 392 270
rect 400 268 422 270
rect 430 268 452 270
rect 460 268 482 270
rect 490 268 512 270
rect 520 268 542 270
rect 550 268 572 270
rect 28 260 32 268
rect 40 260 52 268
rect 70 260 82 268
rect 100 260 112 268
rect 130 260 142 268
rect 160 260 172 268
rect 190 260 202 268
rect 220 260 232 268
rect 250 260 262 268
rect 280 260 292 268
rect 310 260 322 268
rect 340 260 352 268
rect 370 260 382 268
rect 400 260 412 268
rect 430 260 442 268
rect 460 260 472 268
rect 490 260 502 268
rect 520 260 532 268
rect 550 260 562 268
rect 570 260 572 268
rect 28 258 62 260
rect 70 258 92 260
rect 100 258 122 260
rect 130 258 152 260
rect 160 258 182 260
rect 190 258 212 260
rect 220 258 242 260
rect 250 258 272 260
rect 280 258 302 260
rect 310 258 332 260
rect 340 258 362 260
rect 370 258 392 260
rect 400 258 422 260
rect 430 258 452 260
rect 460 258 482 260
rect 490 258 512 260
rect 520 258 542 260
rect 550 258 572 260
rect 28 250 42 258
rect 50 250 62 258
rect 80 250 92 258
rect 110 250 122 258
rect 140 250 152 258
rect 170 250 182 258
rect 200 250 212 258
rect 230 250 242 258
rect 260 250 272 258
rect 290 250 302 258
rect 320 250 332 258
rect 350 250 362 258
rect 380 250 392 258
rect 410 250 422 258
rect 440 250 452 258
rect 470 250 482 258
rect 500 250 512 258
rect 530 250 542 258
rect 560 250 572 258
rect 28 248 62 250
rect 70 248 92 250
rect 100 248 122 250
rect 130 248 152 250
rect 160 248 182 250
rect 190 248 212 250
rect 220 248 242 250
rect 250 248 272 250
rect 280 248 302 250
rect 310 248 332 250
rect 340 248 362 250
rect 370 248 392 250
rect 400 248 422 250
rect 430 248 452 250
rect 460 248 482 250
rect 490 248 512 250
rect 520 248 542 250
rect 550 248 572 250
rect 28 240 32 248
rect 40 240 52 248
rect 28 238 62 240
rect 28 230 42 238
rect 50 230 62 238
rect 28 228 62 230
rect 28 220 32 228
rect 40 220 52 228
rect 70 220 82 248
rect 100 240 112 248
rect 130 240 142 248
rect 160 240 172 248
rect 190 240 202 248
rect 220 240 232 248
rect 250 240 262 248
rect 280 240 292 248
rect 310 240 322 248
rect 340 240 352 248
rect 370 240 382 248
rect 400 240 412 248
rect 430 240 442 248
rect 460 240 472 248
rect 490 240 502 248
rect 520 240 532 248
rect 550 240 562 248
rect 570 240 572 248
rect 90 228 502 240
rect 510 238 542 240
rect 550 238 572 240
rect 510 230 522 238
rect 530 230 542 238
rect 560 230 572 238
rect 510 228 542 230
rect 550 228 572 230
rect 100 220 112 228
rect 130 220 142 228
rect 160 220 172 228
rect 190 220 202 228
rect 220 220 232 228
rect 250 220 262 228
rect 280 220 292 228
rect 310 220 322 228
rect 340 220 352 228
rect 370 220 382 228
rect 400 220 412 228
rect 430 220 442 228
rect 460 220 472 228
rect 490 220 502 228
rect 520 220 532 228
rect 550 220 562 228
rect 570 220 572 228
rect 28 218 62 220
rect 70 218 92 220
rect 100 218 122 220
rect 130 218 152 220
rect 160 218 182 220
rect 190 218 212 220
rect 220 218 242 220
rect 250 218 272 220
rect 280 218 302 220
rect 310 218 332 220
rect 340 218 362 220
rect 370 218 392 220
rect 400 218 422 220
rect 430 218 452 220
rect 460 218 482 220
rect 490 218 512 220
rect 520 218 542 220
rect 550 218 572 220
rect 28 210 42 218
rect 50 210 62 218
rect 80 210 92 218
rect 110 210 122 218
rect 140 210 152 218
rect 170 210 182 218
rect 200 210 212 218
rect 230 210 242 218
rect 260 210 272 218
rect 290 210 302 218
rect 320 210 332 218
rect 350 210 362 218
rect 380 210 392 218
rect 410 210 422 218
rect 440 210 452 218
rect 470 210 482 218
rect 500 210 512 218
rect 530 210 542 218
rect 560 210 572 218
rect 28 208 62 210
rect 70 208 92 210
rect 100 208 122 210
rect 130 208 152 210
rect 160 208 182 210
rect 190 208 212 210
rect 220 208 242 210
rect 250 208 272 210
rect 280 208 302 210
rect 310 208 332 210
rect 340 208 362 210
rect 370 208 392 210
rect 400 208 422 210
rect 430 208 452 210
rect 460 208 482 210
rect 490 208 512 210
rect 520 208 542 210
rect 550 208 572 210
rect 28 200 32 208
rect 40 200 52 208
rect 70 200 82 208
rect 100 200 112 208
rect 130 200 142 208
rect 160 200 172 208
rect 190 200 202 208
rect 220 200 232 208
rect 250 200 262 208
rect 280 200 292 208
rect 310 200 322 208
rect 340 200 352 208
rect 370 200 382 208
rect 400 200 412 208
rect 430 200 442 208
rect 460 200 472 208
rect 490 200 502 208
rect 520 200 532 208
rect 550 200 562 208
rect 570 200 572 208
rect 28 198 62 200
rect 70 198 92 200
rect 100 198 122 200
rect 130 198 152 200
rect 160 198 182 200
rect 190 198 212 200
rect 220 198 242 200
rect 250 198 272 200
rect 280 198 302 200
rect 310 198 332 200
rect 340 198 362 200
rect 370 198 392 200
rect 400 198 422 200
rect 430 198 452 200
rect 460 198 482 200
rect 490 198 512 200
rect 520 198 542 200
rect 550 198 572 200
rect 28 190 42 198
rect 50 190 62 198
rect 80 190 92 198
rect 110 190 122 198
rect 140 190 152 198
rect 170 190 182 198
rect 200 190 212 198
rect 230 190 242 198
rect 260 190 272 198
rect 290 190 302 198
rect 320 190 332 198
rect 350 190 362 198
rect 380 190 392 198
rect 410 190 422 198
rect 440 190 452 198
rect 470 190 482 198
rect 500 190 512 198
rect 530 190 542 198
rect 560 190 572 198
rect 28 188 62 190
rect 70 188 92 190
rect 100 188 122 190
rect 130 188 152 190
rect 160 188 182 190
rect 190 188 212 190
rect 220 188 242 190
rect 250 188 272 190
rect 280 188 302 190
rect 310 188 332 190
rect 340 188 362 190
rect 370 188 392 190
rect 400 188 422 190
rect 430 188 452 190
rect 460 188 482 190
rect 490 188 512 190
rect 520 188 542 190
rect 550 188 572 190
rect 28 180 32 188
rect 40 180 52 188
rect 70 180 82 188
rect 100 180 112 188
rect 130 180 142 188
rect 160 180 172 188
rect 190 180 202 188
rect 220 180 232 188
rect 250 180 262 188
rect 280 180 292 188
rect 310 180 322 188
rect 340 180 352 188
rect 370 180 382 188
rect 400 180 412 188
rect 430 180 442 188
rect 460 180 472 188
rect 490 180 502 188
rect 520 180 532 188
rect 550 180 562 188
rect 570 180 572 188
rect 28 178 62 180
rect 70 178 92 180
rect 100 178 122 180
rect 130 178 152 180
rect 160 178 182 180
rect 190 178 212 180
rect 220 178 242 180
rect 250 178 272 180
rect 280 178 302 180
rect 310 178 332 180
rect 340 178 362 180
rect 370 178 392 180
rect 400 178 422 180
rect 430 178 452 180
rect 460 178 482 180
rect 490 178 512 180
rect 520 178 542 180
rect 550 178 572 180
rect 28 170 42 178
rect 50 170 62 178
rect 80 170 92 178
rect 110 170 122 178
rect 140 170 152 178
rect 170 170 182 178
rect 200 170 212 178
rect 230 170 242 178
rect 260 170 272 178
rect 290 170 302 178
rect 320 170 332 178
rect 350 170 362 178
rect 380 170 392 178
rect 410 170 422 178
rect 440 170 452 178
rect 470 170 482 178
rect 500 170 512 178
rect 530 170 542 178
rect 560 170 572 178
rect 28 168 62 170
rect 70 168 92 170
rect 100 168 122 170
rect 130 168 152 170
rect 160 168 182 170
rect 190 168 212 170
rect 220 168 242 170
rect 250 168 272 170
rect 280 168 302 170
rect 310 168 332 170
rect 340 168 362 170
rect 370 168 392 170
rect 400 168 422 170
rect 430 168 452 170
rect 460 168 482 170
rect 490 168 512 170
rect 520 168 542 170
rect 550 168 572 170
rect 28 160 32 168
rect 40 160 52 168
rect 70 160 82 168
rect 100 160 112 168
rect 130 160 142 168
rect 160 160 172 168
rect 190 160 202 168
rect 220 160 232 168
rect 250 160 262 168
rect 280 160 292 168
rect 310 160 322 168
rect 340 160 352 168
rect 370 160 382 168
rect 400 160 412 168
rect 430 160 442 168
rect 460 160 472 168
rect 490 160 502 168
rect 520 160 532 168
rect 550 160 562 168
rect 570 160 572 168
rect 28 158 62 160
rect 70 158 92 160
rect 28 150 42 158
rect 50 150 62 158
rect 80 150 92 158
rect 28 148 62 150
rect 70 148 92 150
rect 100 148 502 160
rect 510 158 542 160
rect 550 158 572 160
rect 510 150 522 158
rect 530 150 542 158
rect 560 150 572 158
rect 510 148 542 150
rect 550 148 572 150
rect 28 140 32 148
rect 40 140 52 148
rect 70 140 82 148
rect 100 140 112 148
rect 130 140 142 148
rect 160 140 172 148
rect 190 140 202 148
rect 220 140 232 148
rect 250 140 262 148
rect 280 140 292 148
rect 310 140 322 148
rect 340 140 352 148
rect 370 140 382 148
rect 400 140 412 148
rect 430 140 442 148
rect 460 140 472 148
rect 490 140 502 148
rect 520 140 532 148
rect 550 140 562 148
rect 570 140 572 148
rect 28 138 62 140
rect 70 138 92 140
rect 100 138 122 140
rect 130 138 152 140
rect 160 138 182 140
rect 190 138 212 140
rect 220 138 242 140
rect 250 138 272 140
rect 280 138 302 140
rect 310 138 332 140
rect 340 138 362 140
rect 370 138 392 140
rect 400 138 422 140
rect 430 138 452 140
rect 460 138 482 140
rect 490 138 512 140
rect 520 138 542 140
rect 550 138 572 140
rect 28 130 42 138
rect 50 130 62 138
rect 80 130 92 138
rect 110 130 122 138
rect 140 130 152 138
rect 170 130 182 138
rect 200 130 212 138
rect 230 130 242 138
rect 260 130 272 138
rect 290 130 302 138
rect 320 130 332 138
rect 350 130 362 138
rect 380 130 392 138
rect 410 130 422 138
rect 440 130 452 138
rect 470 130 482 138
rect 500 130 512 138
rect 530 130 542 138
rect 560 130 572 138
rect 28 128 62 130
rect 70 128 92 130
rect 100 128 122 130
rect 130 128 152 130
rect 160 128 182 130
rect 190 128 212 130
rect 220 128 242 130
rect 250 128 272 130
rect 280 128 302 130
rect 310 128 332 130
rect 340 128 362 130
rect 370 128 392 130
rect 400 128 422 130
rect 430 128 452 130
rect 460 128 482 130
rect 490 128 512 130
rect 520 128 542 130
rect 550 128 572 130
rect 28 120 32 128
rect 40 120 52 128
rect 70 120 82 128
rect 100 120 112 128
rect 130 120 142 128
rect 160 120 172 128
rect 190 120 202 128
rect 220 120 232 128
rect 250 120 262 128
rect 280 120 292 128
rect 310 120 322 128
rect 340 120 352 128
rect 370 120 382 128
rect 400 120 412 128
rect 430 120 442 128
rect 460 120 472 128
rect 490 120 502 128
rect 520 120 532 128
rect 550 120 562 128
rect 570 120 572 128
rect 28 118 62 120
rect 70 118 92 120
rect 100 118 122 120
rect 130 118 152 120
rect 160 118 182 120
rect 190 118 212 120
rect 220 118 242 120
rect 250 118 272 120
rect 280 118 302 120
rect 310 118 332 120
rect 340 118 362 120
rect 370 118 392 120
rect 400 118 422 120
rect 430 118 452 120
rect 460 118 482 120
rect 490 118 512 120
rect 520 118 542 120
rect 550 118 572 120
rect 28 110 42 118
rect 50 110 62 118
rect 80 110 92 118
rect 110 110 122 118
rect 140 110 152 118
rect 170 110 182 118
rect 200 110 212 118
rect 230 110 242 118
rect 260 110 272 118
rect 290 110 302 118
rect 320 110 332 118
rect 350 110 362 118
rect 380 110 392 118
rect 410 110 422 118
rect 440 110 452 118
rect 470 110 482 118
rect 500 110 512 118
rect 530 110 542 118
rect 560 110 572 118
rect 28 108 62 110
rect 70 108 92 110
rect 100 108 122 110
rect 130 108 152 110
rect 160 108 182 110
rect 190 108 212 110
rect 220 108 242 110
rect 250 108 272 110
rect 280 108 302 110
rect 310 108 332 110
rect 340 108 362 110
rect 370 108 392 110
rect 400 108 422 110
rect 430 108 452 110
rect 460 108 482 110
rect 490 108 512 110
rect 520 108 542 110
rect 550 108 572 110
rect 28 100 32 108
rect 40 100 52 108
rect 70 100 82 108
rect 100 100 112 108
rect 130 100 142 108
rect 160 100 172 108
rect 190 100 202 108
rect 220 100 232 108
rect 250 100 262 108
rect 280 100 292 108
rect 310 100 322 108
rect 340 100 352 108
rect 370 100 382 108
rect 400 100 412 108
rect 430 100 442 108
rect 460 100 472 108
rect 490 100 502 108
rect 520 100 532 108
rect 550 100 562 108
rect 570 100 572 108
rect 28 98 62 100
rect 70 98 92 100
rect 100 98 122 100
rect 130 98 152 100
rect 160 98 182 100
rect 190 98 212 100
rect 220 98 242 100
rect 250 98 272 100
rect 280 98 302 100
rect 310 98 332 100
rect 340 98 362 100
rect 370 98 392 100
rect 400 98 422 100
rect 430 98 452 100
rect 460 98 482 100
rect 490 98 512 100
rect 520 98 542 100
rect 550 98 572 100
rect 28 90 42 98
rect 50 90 62 98
rect 80 90 92 98
rect 110 90 122 98
rect 140 90 152 98
rect 170 90 182 98
rect 200 90 212 98
rect 230 90 242 98
rect 260 90 272 98
rect 290 90 302 98
rect 320 90 332 98
rect 350 90 362 98
rect 380 90 392 98
rect 410 90 422 98
rect 440 90 452 98
rect 470 90 482 98
rect 500 90 512 98
rect 530 90 542 98
rect 560 90 572 98
rect 28 88 62 90
rect 70 88 92 90
rect 100 88 122 90
rect 130 88 152 90
rect 160 88 182 90
rect 190 88 212 90
rect 220 88 242 90
rect 250 88 272 90
rect 280 88 302 90
rect 310 88 332 90
rect 340 88 362 90
rect 370 88 392 90
rect 400 88 422 90
rect 430 88 452 90
rect 460 88 482 90
rect 490 88 512 90
rect 520 88 542 90
rect 550 88 572 90
rect 28 80 32 88
rect 40 80 52 88
rect 70 80 82 88
rect 100 80 112 88
rect 130 80 142 88
rect 160 80 172 88
rect 190 80 202 88
rect 220 80 232 88
rect 250 80 262 88
rect 280 80 292 88
rect 310 80 322 88
rect 340 80 352 88
rect 370 80 382 88
rect 400 80 412 88
rect 430 80 442 88
rect 460 80 472 88
rect 490 80 502 88
rect 520 80 532 88
rect 550 80 562 88
rect 570 80 572 88
rect 28 78 62 80
rect 70 78 92 80
rect 100 78 122 80
rect 130 78 152 80
rect 160 78 182 80
rect 190 78 212 80
rect 220 78 242 80
rect 250 78 272 80
rect 280 78 302 80
rect 310 78 332 80
rect 340 78 362 80
rect 370 78 392 80
rect 400 78 422 80
rect 430 78 452 80
rect 460 78 482 80
rect 490 78 512 80
rect 520 78 542 80
rect 550 78 572 80
rect 28 70 42 78
rect 50 70 62 78
rect 80 70 92 78
rect 110 70 122 78
rect 140 70 152 78
rect 170 70 182 78
rect 200 70 212 78
rect 230 70 242 78
rect 260 70 272 78
rect 290 70 302 78
rect 320 70 332 78
rect 350 70 362 78
rect 380 70 392 78
rect 410 70 422 78
rect 440 70 452 78
rect 470 70 482 78
rect 500 70 512 78
rect 530 70 542 78
rect 560 70 572 78
rect 28 68 62 70
rect 70 68 92 70
rect 100 68 122 70
rect 130 68 152 70
rect 160 68 182 70
rect 190 68 212 70
rect 220 68 242 70
rect 250 68 272 70
rect 280 68 302 70
rect 310 68 332 70
rect 340 68 362 70
rect 370 68 392 70
rect 400 68 422 70
rect 430 68 452 70
rect 460 68 482 70
rect 490 68 512 70
rect 520 68 542 70
rect 550 68 572 70
rect 28 60 32 68
rect 40 60 52 68
rect 70 60 82 68
rect 100 60 112 68
rect 130 60 142 68
rect 160 60 172 68
rect 190 60 202 68
rect 220 60 232 68
rect 250 60 262 68
rect 280 60 292 68
rect 310 60 322 68
rect 340 60 352 68
rect 370 60 382 68
rect 400 60 412 68
rect 430 60 442 68
rect 460 60 472 68
rect 490 60 502 68
rect 520 60 532 68
rect 550 60 562 68
rect 570 60 572 68
rect 28 58 62 60
rect 70 58 92 60
rect 100 58 122 60
rect 130 58 152 60
rect 160 58 182 60
rect 190 58 212 60
rect 220 58 242 60
rect 250 58 272 60
rect 280 58 302 60
rect 310 58 332 60
rect 340 58 362 60
rect 370 58 392 60
rect 400 58 422 60
rect 430 58 452 60
rect 460 58 482 60
rect 490 58 512 60
rect 520 58 542 60
rect 550 58 572 60
rect 28 50 42 58
rect 50 50 62 58
rect 80 50 92 58
rect 110 50 122 58
rect 140 50 152 58
rect 170 50 182 58
rect 200 50 212 58
rect 230 50 242 58
rect 260 50 272 58
rect 290 50 302 58
rect 320 50 332 58
rect 350 50 362 58
rect 380 50 392 58
rect 410 50 422 58
rect 440 50 452 58
rect 470 50 482 58
rect 500 50 512 58
rect 530 50 542 58
rect 560 50 572 58
rect 28 48 62 50
rect 70 48 92 50
rect 100 48 122 50
rect 130 48 152 50
rect 160 48 182 50
rect 190 48 212 50
rect 220 48 242 50
rect 250 48 272 50
rect 280 48 302 50
rect 310 48 332 50
rect 340 48 362 50
rect 370 48 392 50
rect 400 48 422 50
rect 430 48 452 50
rect 460 48 482 50
rect 490 48 512 50
rect 520 48 542 50
rect 550 48 572 50
rect 28 40 32 48
rect 40 40 52 48
rect 70 40 82 48
rect 100 40 112 48
rect 130 40 142 48
rect 160 40 172 48
rect 190 40 202 48
rect 220 40 232 48
rect 250 40 262 48
rect 280 40 292 48
rect 310 40 322 48
rect 340 40 352 48
rect 370 40 382 48
rect 400 40 412 48
rect 430 40 442 48
rect 460 40 472 48
rect 490 40 502 48
rect 520 40 532 48
rect 550 40 562 48
rect 570 40 572 48
rect 28 38 62 40
rect 70 38 92 40
rect 100 38 122 40
rect 130 38 152 40
rect 160 38 182 40
rect 190 38 212 40
rect 220 38 242 40
rect 250 38 272 40
rect 280 38 302 40
rect 310 38 332 40
rect 340 38 362 40
rect 370 38 392 40
rect 400 38 422 40
rect 430 38 452 40
rect 460 38 482 40
rect 490 38 512 40
rect 520 38 542 40
rect 550 38 572 40
rect 28 30 42 38
rect 50 30 62 38
rect 80 30 92 38
rect 110 30 122 38
rect 140 30 152 38
rect 170 30 182 38
rect 200 30 212 38
rect 230 30 242 38
rect 260 30 272 38
rect 290 30 302 38
rect 320 30 332 38
rect 350 30 362 38
rect 380 30 392 38
rect 410 30 422 38
rect 440 30 452 38
rect 470 30 482 38
rect 500 30 512 38
rect 530 30 542 38
rect 560 30 572 38
rect 28 28 572 30
<< nsubstratendiff >>
rect 40 1298 560 1300
rect 40 1290 46 1298
rect 54 1290 66 1298
rect 84 1290 96 1298
rect 114 1290 126 1298
rect 144 1290 156 1298
rect 174 1290 186 1298
rect 204 1290 216 1298
rect 234 1290 246 1298
rect 264 1290 276 1298
rect 294 1290 306 1298
rect 324 1290 336 1298
rect 354 1290 366 1298
rect 384 1290 396 1298
rect 414 1290 426 1298
rect 444 1290 456 1298
rect 474 1290 486 1298
rect 504 1290 516 1298
rect 534 1290 546 1298
rect 554 1290 560 1298
rect 40 1288 76 1290
rect 84 1288 106 1290
rect 114 1288 136 1290
rect 144 1288 166 1290
rect 174 1288 196 1290
rect 204 1288 226 1290
rect 234 1288 256 1290
rect 264 1288 286 1290
rect 294 1288 316 1290
rect 324 1288 346 1290
rect 354 1288 376 1290
rect 384 1288 406 1290
rect 414 1288 436 1290
rect 444 1288 466 1290
rect 474 1288 496 1290
rect 504 1288 526 1290
rect 534 1288 560 1290
rect 40 1280 56 1288
rect 64 1280 76 1288
rect 94 1280 106 1288
rect 124 1280 136 1288
rect 154 1280 166 1288
rect 184 1280 196 1288
rect 214 1280 226 1288
rect 244 1280 256 1288
rect 274 1280 286 1288
rect 304 1280 316 1288
rect 334 1280 346 1288
rect 364 1280 376 1288
rect 394 1280 406 1288
rect 424 1280 436 1288
rect 454 1280 466 1288
rect 484 1280 496 1288
rect 514 1280 526 1288
rect 544 1280 560 1288
rect 40 1278 76 1280
rect 84 1278 106 1280
rect 114 1278 136 1280
rect 144 1278 166 1280
rect 174 1278 196 1280
rect 204 1278 226 1280
rect 234 1278 256 1280
rect 264 1278 286 1280
rect 294 1278 316 1280
rect 324 1278 346 1280
rect 354 1278 376 1280
rect 384 1278 406 1280
rect 414 1278 436 1280
rect 444 1278 466 1280
rect 474 1278 496 1280
rect 504 1278 526 1280
rect 534 1278 560 1280
rect 40 1270 46 1278
rect 54 1270 66 1278
rect 84 1270 96 1278
rect 114 1270 126 1278
rect 144 1270 156 1278
rect 174 1270 186 1278
rect 204 1270 216 1278
rect 234 1270 246 1278
rect 264 1270 276 1278
rect 294 1270 306 1278
rect 324 1270 336 1278
rect 354 1270 366 1278
rect 384 1270 396 1278
rect 414 1270 426 1278
rect 444 1270 456 1278
rect 474 1270 486 1278
rect 504 1270 516 1278
rect 534 1270 546 1278
rect 554 1270 560 1278
rect 40 1268 76 1270
rect 84 1268 106 1270
rect 114 1268 136 1270
rect 144 1268 166 1270
rect 174 1268 196 1270
rect 204 1268 226 1270
rect 234 1268 256 1270
rect 264 1268 286 1270
rect 294 1268 316 1270
rect 324 1268 346 1270
rect 354 1268 376 1270
rect 384 1268 406 1270
rect 414 1268 436 1270
rect 444 1268 466 1270
rect 474 1268 496 1270
rect 504 1268 526 1270
rect 534 1268 560 1270
rect 40 1260 56 1268
rect 64 1260 76 1268
rect 94 1260 106 1268
rect 124 1260 136 1268
rect 154 1260 166 1268
rect 184 1260 196 1268
rect 214 1260 226 1268
rect 244 1260 256 1268
rect 274 1260 286 1268
rect 304 1260 316 1268
rect 334 1260 346 1268
rect 364 1260 376 1268
rect 394 1260 406 1268
rect 424 1260 436 1268
rect 454 1260 466 1268
rect 484 1260 496 1268
rect 514 1260 526 1268
rect 544 1260 560 1268
rect 40 1258 76 1260
rect 84 1258 106 1260
rect 114 1258 136 1260
rect 144 1258 166 1260
rect 174 1258 196 1260
rect 204 1258 226 1260
rect 234 1258 256 1260
rect 264 1258 286 1260
rect 294 1258 316 1260
rect 324 1258 346 1260
rect 354 1258 376 1260
rect 384 1258 406 1260
rect 414 1258 436 1260
rect 444 1258 466 1260
rect 474 1258 496 1260
rect 504 1258 526 1260
rect 534 1258 560 1260
rect 40 1250 46 1258
rect 54 1250 66 1258
rect 84 1250 96 1258
rect 114 1250 126 1258
rect 144 1250 156 1258
rect 174 1250 186 1258
rect 204 1250 216 1258
rect 234 1250 246 1258
rect 264 1250 276 1258
rect 294 1250 306 1258
rect 324 1250 336 1258
rect 354 1250 366 1258
rect 384 1250 396 1258
rect 414 1250 426 1258
rect 444 1250 456 1258
rect 474 1250 486 1258
rect 504 1250 516 1258
rect 534 1250 546 1258
rect 554 1250 560 1258
rect 40 1248 76 1250
rect 84 1248 106 1250
rect 114 1248 136 1250
rect 144 1248 166 1250
rect 174 1248 196 1250
rect 204 1248 226 1250
rect 234 1248 256 1250
rect 264 1248 286 1250
rect 294 1248 316 1250
rect 324 1248 346 1250
rect 354 1248 376 1250
rect 384 1248 406 1250
rect 414 1248 436 1250
rect 444 1248 466 1250
rect 474 1248 496 1250
rect 504 1248 526 1250
rect 534 1248 560 1250
rect 40 1240 56 1248
rect 64 1240 76 1248
rect 94 1240 106 1248
rect 124 1240 136 1248
rect 154 1240 166 1248
rect 184 1240 196 1248
rect 214 1240 226 1248
rect 244 1240 256 1248
rect 274 1240 286 1248
rect 304 1240 316 1248
rect 334 1240 346 1248
rect 364 1240 376 1248
rect 394 1240 406 1248
rect 424 1240 436 1248
rect 454 1240 466 1248
rect 484 1240 496 1248
rect 514 1240 526 1248
rect 544 1240 560 1248
rect 40 1238 76 1240
rect 84 1238 106 1240
rect 114 1238 136 1240
rect 144 1238 166 1240
rect 174 1238 196 1240
rect 204 1238 226 1240
rect 234 1238 256 1240
rect 264 1238 286 1240
rect 294 1238 316 1240
rect 324 1238 346 1240
rect 354 1238 376 1240
rect 384 1238 406 1240
rect 414 1238 436 1240
rect 444 1238 466 1240
rect 474 1238 496 1240
rect 504 1238 526 1240
rect 534 1238 560 1240
rect 40 1230 46 1238
rect 54 1230 66 1238
rect 84 1230 96 1238
rect 114 1230 126 1238
rect 144 1230 156 1238
rect 174 1230 186 1238
rect 204 1230 216 1238
rect 234 1230 246 1238
rect 264 1230 276 1238
rect 294 1230 306 1238
rect 324 1230 336 1238
rect 354 1230 366 1238
rect 384 1230 396 1238
rect 414 1230 426 1238
rect 444 1230 456 1238
rect 474 1230 486 1238
rect 504 1230 516 1238
rect 534 1230 546 1238
rect 554 1230 560 1238
rect 40 1228 76 1230
rect 84 1228 106 1230
rect 114 1228 136 1230
rect 144 1228 166 1230
rect 174 1228 196 1230
rect 204 1228 226 1230
rect 234 1228 256 1230
rect 264 1228 286 1230
rect 294 1228 316 1230
rect 324 1228 346 1230
rect 354 1228 376 1230
rect 384 1228 406 1230
rect 414 1228 436 1230
rect 444 1228 466 1230
rect 474 1228 496 1230
rect 504 1228 526 1230
rect 534 1228 560 1230
rect 40 1220 56 1228
rect 64 1220 76 1228
rect 94 1220 106 1228
rect 124 1220 136 1228
rect 154 1220 166 1228
rect 184 1220 196 1228
rect 214 1220 226 1228
rect 244 1220 256 1228
rect 274 1220 286 1228
rect 304 1220 316 1228
rect 334 1220 346 1228
rect 364 1220 376 1228
rect 394 1220 406 1228
rect 424 1220 436 1228
rect 454 1220 466 1228
rect 484 1220 496 1228
rect 514 1220 526 1228
rect 544 1220 560 1228
rect 40 1218 76 1220
rect 84 1218 106 1220
rect 114 1218 136 1220
rect 144 1218 166 1220
rect 174 1218 196 1220
rect 204 1218 226 1220
rect 234 1218 256 1220
rect 264 1218 286 1220
rect 294 1218 316 1220
rect 324 1218 346 1220
rect 354 1218 376 1220
rect 384 1218 406 1220
rect 414 1218 436 1220
rect 444 1218 466 1220
rect 474 1218 496 1220
rect 504 1218 526 1220
rect 534 1218 560 1220
rect 40 1210 46 1218
rect 54 1210 66 1218
rect 84 1210 96 1218
rect 114 1210 126 1218
rect 144 1210 156 1218
rect 174 1210 186 1218
rect 204 1210 216 1218
rect 234 1210 246 1218
rect 264 1210 276 1218
rect 294 1210 306 1218
rect 324 1210 336 1218
rect 354 1210 366 1218
rect 384 1210 396 1218
rect 414 1210 426 1218
rect 444 1210 456 1218
rect 474 1210 486 1218
rect 504 1210 516 1218
rect 534 1210 546 1218
rect 554 1210 560 1218
rect 40 1208 76 1210
rect 84 1208 106 1210
rect 114 1208 136 1210
rect 144 1208 166 1210
rect 174 1208 196 1210
rect 204 1208 226 1210
rect 234 1208 256 1210
rect 264 1208 286 1210
rect 294 1208 316 1210
rect 324 1208 346 1210
rect 354 1208 376 1210
rect 384 1208 406 1210
rect 414 1208 436 1210
rect 444 1208 466 1210
rect 474 1208 496 1210
rect 504 1208 526 1210
rect 534 1208 560 1210
rect 40 1200 56 1208
rect 64 1200 76 1208
rect 94 1200 106 1208
rect 124 1200 136 1208
rect 154 1200 166 1208
rect 184 1200 196 1208
rect 214 1200 226 1208
rect 244 1200 256 1208
rect 274 1200 286 1208
rect 304 1200 316 1208
rect 334 1200 346 1208
rect 364 1200 376 1208
rect 394 1200 406 1208
rect 424 1200 436 1208
rect 454 1200 466 1208
rect 484 1200 496 1208
rect 514 1200 526 1208
rect 544 1200 560 1208
rect 40 1198 76 1200
rect 84 1198 106 1200
rect 114 1198 136 1200
rect 144 1198 166 1200
rect 174 1198 196 1200
rect 204 1198 226 1200
rect 234 1198 256 1200
rect 264 1198 286 1200
rect 294 1198 316 1200
rect 324 1198 346 1200
rect 354 1198 376 1200
rect 384 1198 406 1200
rect 414 1198 436 1200
rect 444 1198 466 1200
rect 474 1198 496 1200
rect 504 1198 526 1200
rect 534 1198 560 1200
rect 40 1190 46 1198
rect 54 1190 66 1198
rect 84 1190 96 1198
rect 114 1190 126 1198
rect 144 1190 156 1198
rect 174 1190 186 1198
rect 204 1190 216 1198
rect 234 1190 246 1198
rect 264 1190 276 1198
rect 294 1190 306 1198
rect 324 1190 336 1198
rect 354 1190 366 1198
rect 384 1190 396 1198
rect 414 1190 426 1198
rect 444 1190 456 1198
rect 474 1190 486 1198
rect 504 1190 516 1198
rect 534 1190 546 1198
rect 554 1190 560 1198
rect 40 1188 76 1190
rect 84 1188 526 1190
rect 534 1188 560 1190
rect 40 1180 56 1188
rect 64 1180 76 1188
rect 94 1180 506 1188
rect 514 1180 526 1188
rect 544 1180 560 1188
rect 40 1178 76 1180
rect 84 1178 526 1180
rect 534 1178 560 1180
rect 40 1170 46 1178
rect 54 1170 66 1178
rect 84 1170 96 1178
rect 114 1170 126 1178
rect 144 1170 156 1178
rect 174 1170 186 1178
rect 204 1170 216 1178
rect 234 1170 246 1178
rect 264 1170 276 1178
rect 294 1170 306 1178
rect 324 1170 336 1178
rect 354 1170 366 1178
rect 384 1170 396 1178
rect 414 1170 426 1178
rect 444 1170 456 1178
rect 474 1170 486 1178
rect 504 1170 516 1178
rect 534 1170 546 1178
rect 554 1170 560 1178
rect 40 1168 76 1170
rect 84 1168 106 1170
rect 114 1168 136 1170
rect 144 1168 166 1170
rect 174 1168 196 1170
rect 204 1168 226 1170
rect 234 1168 256 1170
rect 264 1168 286 1170
rect 294 1168 316 1170
rect 324 1168 346 1170
rect 354 1168 376 1170
rect 384 1168 406 1170
rect 414 1168 436 1170
rect 444 1168 466 1170
rect 474 1168 496 1170
rect 504 1168 526 1170
rect 534 1168 560 1170
rect 40 1160 56 1168
rect 64 1160 76 1168
rect 94 1160 106 1168
rect 124 1160 136 1168
rect 154 1160 166 1168
rect 184 1160 196 1168
rect 214 1160 226 1168
rect 244 1160 256 1168
rect 274 1160 286 1168
rect 304 1160 316 1168
rect 334 1160 346 1168
rect 364 1160 376 1168
rect 394 1160 406 1168
rect 424 1160 436 1168
rect 454 1160 466 1168
rect 484 1160 496 1168
rect 514 1160 526 1168
rect 544 1160 560 1168
rect 40 1158 76 1160
rect 84 1158 106 1160
rect 114 1158 136 1160
rect 144 1158 166 1160
rect 174 1158 196 1160
rect 204 1158 226 1160
rect 234 1158 256 1160
rect 264 1158 286 1160
rect 294 1158 316 1160
rect 324 1158 346 1160
rect 354 1158 376 1160
rect 384 1158 406 1160
rect 414 1158 436 1160
rect 444 1158 466 1160
rect 474 1158 496 1160
rect 504 1158 526 1160
rect 534 1158 560 1160
rect 40 1150 46 1158
rect 54 1150 66 1158
rect 84 1150 96 1158
rect 114 1150 126 1158
rect 144 1150 156 1158
rect 174 1150 186 1158
rect 204 1150 216 1158
rect 234 1150 246 1158
rect 264 1150 276 1158
rect 294 1150 306 1158
rect 324 1150 336 1158
rect 354 1150 366 1158
rect 384 1150 396 1158
rect 414 1150 426 1158
rect 444 1150 456 1158
rect 474 1150 486 1158
rect 504 1150 516 1158
rect 534 1150 546 1158
rect 554 1150 560 1158
rect 40 1148 76 1150
rect 84 1148 106 1150
rect 114 1148 136 1150
rect 144 1148 166 1150
rect 174 1148 196 1150
rect 204 1148 226 1150
rect 234 1148 256 1150
rect 264 1148 286 1150
rect 294 1148 316 1150
rect 324 1148 346 1150
rect 354 1148 376 1150
rect 384 1148 406 1150
rect 414 1148 436 1150
rect 444 1148 466 1150
rect 474 1148 496 1150
rect 504 1148 526 1150
rect 534 1148 560 1150
rect 40 1140 56 1148
rect 64 1140 76 1148
rect 94 1140 106 1148
rect 124 1140 136 1148
rect 154 1140 166 1148
rect 184 1140 196 1148
rect 214 1140 226 1148
rect 244 1140 256 1148
rect 274 1140 286 1148
rect 304 1140 316 1148
rect 334 1140 346 1148
rect 364 1140 376 1148
rect 394 1140 406 1148
rect 424 1140 436 1148
rect 454 1140 466 1148
rect 484 1140 496 1148
rect 514 1140 526 1148
rect 544 1140 560 1148
rect 40 1138 76 1140
rect 84 1138 106 1140
rect 114 1138 136 1140
rect 144 1138 166 1140
rect 174 1138 196 1140
rect 204 1138 226 1140
rect 234 1138 256 1140
rect 264 1138 286 1140
rect 294 1138 316 1140
rect 324 1138 346 1140
rect 354 1138 376 1140
rect 384 1138 406 1140
rect 414 1138 436 1140
rect 444 1138 466 1140
rect 474 1138 496 1140
rect 504 1138 526 1140
rect 534 1138 560 1140
rect 40 1130 46 1138
rect 54 1130 66 1138
rect 84 1130 96 1138
rect 114 1130 126 1138
rect 144 1130 156 1138
rect 174 1130 186 1138
rect 204 1130 216 1138
rect 234 1130 246 1138
rect 264 1130 276 1138
rect 294 1130 306 1138
rect 324 1130 336 1138
rect 354 1130 366 1138
rect 384 1130 396 1138
rect 414 1130 426 1138
rect 444 1130 456 1138
rect 474 1130 486 1138
rect 504 1130 516 1138
rect 534 1130 546 1138
rect 554 1130 560 1138
rect 40 1128 76 1130
rect 84 1128 106 1130
rect 114 1128 136 1130
rect 144 1128 166 1130
rect 174 1128 196 1130
rect 204 1128 226 1130
rect 234 1128 256 1130
rect 264 1128 286 1130
rect 294 1128 316 1130
rect 324 1128 346 1130
rect 354 1128 376 1130
rect 384 1128 406 1130
rect 414 1128 436 1130
rect 444 1128 466 1130
rect 474 1128 496 1130
rect 504 1128 526 1130
rect 534 1128 560 1130
rect 40 1120 56 1128
rect 64 1120 76 1128
rect 94 1120 106 1128
rect 124 1120 136 1128
rect 154 1120 166 1128
rect 184 1120 196 1128
rect 214 1120 226 1128
rect 244 1120 256 1128
rect 274 1120 286 1128
rect 304 1120 316 1128
rect 334 1120 346 1128
rect 364 1120 376 1128
rect 394 1120 406 1128
rect 424 1120 436 1128
rect 454 1120 466 1128
rect 484 1120 496 1128
rect 40 1118 86 1120
rect 40 1110 46 1118
rect 54 1110 66 1118
rect 74 1110 86 1118
rect 40 1108 86 1110
rect 94 1108 506 1120
rect 40 1100 56 1108
rect 64 1100 76 1108
rect 94 1100 106 1108
rect 124 1100 136 1108
rect 154 1100 166 1108
rect 184 1100 196 1108
rect 214 1100 226 1108
rect 244 1100 256 1108
rect 274 1100 286 1108
rect 304 1100 316 1108
rect 334 1100 346 1108
rect 364 1100 376 1108
rect 394 1100 406 1108
rect 424 1100 436 1108
rect 454 1100 466 1108
rect 484 1100 496 1108
rect 514 1100 526 1128
rect 544 1120 560 1128
rect 534 1118 560 1120
rect 534 1110 546 1118
rect 554 1110 560 1118
rect 534 1108 560 1110
rect 544 1100 560 1108
rect 40 1098 76 1100
rect 84 1098 106 1100
rect 114 1098 136 1100
rect 144 1098 166 1100
rect 174 1098 196 1100
rect 204 1098 226 1100
rect 234 1098 256 1100
rect 264 1098 286 1100
rect 294 1098 316 1100
rect 324 1098 346 1100
rect 354 1098 376 1100
rect 384 1098 406 1100
rect 414 1098 436 1100
rect 444 1098 466 1100
rect 474 1098 496 1100
rect 504 1098 526 1100
rect 534 1098 560 1100
rect 40 1090 46 1098
rect 54 1090 66 1098
rect 84 1090 96 1098
rect 114 1090 126 1098
rect 144 1090 156 1098
rect 174 1090 186 1098
rect 204 1090 216 1098
rect 234 1090 246 1098
rect 264 1090 276 1098
rect 294 1090 306 1098
rect 324 1090 336 1098
rect 354 1090 366 1098
rect 384 1090 396 1098
rect 414 1090 426 1098
rect 444 1090 456 1098
rect 474 1090 486 1098
rect 504 1090 516 1098
rect 534 1090 546 1098
rect 554 1090 560 1098
rect 40 1088 76 1090
rect 84 1088 106 1090
rect 114 1088 136 1090
rect 144 1088 166 1090
rect 174 1088 196 1090
rect 204 1088 226 1090
rect 234 1088 256 1090
rect 264 1088 286 1090
rect 294 1088 316 1090
rect 324 1088 346 1090
rect 354 1088 376 1090
rect 384 1088 406 1090
rect 414 1088 436 1090
rect 444 1088 466 1090
rect 474 1088 496 1090
rect 504 1088 526 1090
rect 534 1088 560 1090
rect 40 1080 56 1088
rect 64 1080 76 1088
rect 94 1080 106 1088
rect 124 1080 136 1088
rect 154 1080 166 1088
rect 184 1080 196 1088
rect 214 1080 226 1088
rect 244 1080 256 1088
rect 274 1080 286 1088
rect 304 1080 316 1088
rect 334 1080 346 1088
rect 364 1080 376 1088
rect 394 1080 406 1088
rect 424 1080 436 1088
rect 454 1080 466 1088
rect 484 1080 496 1088
rect 514 1080 526 1088
rect 544 1080 560 1088
rect 40 1078 76 1080
rect 84 1078 106 1080
rect 114 1078 136 1080
rect 144 1078 166 1080
rect 174 1078 196 1080
rect 204 1078 226 1080
rect 234 1078 256 1080
rect 264 1078 286 1080
rect 294 1078 316 1080
rect 324 1078 346 1080
rect 354 1078 376 1080
rect 384 1078 406 1080
rect 414 1078 436 1080
rect 444 1078 466 1080
rect 474 1078 496 1080
rect 504 1078 526 1080
rect 534 1078 560 1080
rect 40 1070 46 1078
rect 54 1070 66 1078
rect 84 1070 96 1078
rect 114 1070 126 1078
rect 144 1070 156 1078
rect 174 1070 186 1078
rect 204 1070 216 1078
rect 234 1070 246 1078
rect 264 1070 276 1078
rect 294 1070 306 1078
rect 324 1070 336 1078
rect 354 1070 366 1078
rect 384 1070 396 1078
rect 414 1070 426 1078
rect 444 1070 456 1078
rect 474 1070 486 1078
rect 504 1070 516 1078
rect 534 1070 546 1078
rect 554 1070 560 1078
rect 40 1068 76 1070
rect 84 1068 106 1070
rect 114 1068 136 1070
rect 144 1068 166 1070
rect 174 1068 196 1070
rect 204 1068 226 1070
rect 234 1068 256 1070
rect 264 1068 286 1070
rect 294 1068 316 1070
rect 324 1068 346 1070
rect 354 1068 376 1070
rect 384 1068 406 1070
rect 414 1068 436 1070
rect 444 1068 466 1070
rect 474 1068 496 1070
rect 504 1068 526 1070
rect 534 1068 560 1070
rect 40 1060 56 1068
rect 64 1060 76 1068
rect 94 1060 106 1068
rect 124 1060 136 1068
rect 154 1060 166 1068
rect 184 1060 196 1068
rect 214 1060 226 1068
rect 244 1060 256 1068
rect 274 1060 286 1068
rect 304 1060 316 1068
rect 334 1060 346 1068
rect 364 1060 376 1068
rect 394 1060 406 1068
rect 424 1060 436 1068
rect 454 1060 466 1068
rect 484 1060 496 1068
rect 514 1060 526 1068
rect 544 1060 560 1068
rect 40 1058 76 1060
rect 84 1058 106 1060
rect 114 1058 136 1060
rect 144 1058 166 1060
rect 174 1058 196 1060
rect 204 1058 226 1060
rect 234 1058 256 1060
rect 264 1058 286 1060
rect 294 1058 316 1060
rect 324 1058 346 1060
rect 354 1058 376 1060
rect 384 1058 406 1060
rect 414 1058 436 1060
rect 444 1058 466 1060
rect 474 1058 496 1060
rect 504 1058 526 1060
rect 534 1058 560 1060
rect 40 1050 46 1058
rect 54 1050 66 1058
rect 84 1050 96 1058
rect 114 1050 126 1058
rect 144 1050 156 1058
rect 174 1050 186 1058
rect 204 1050 216 1058
rect 234 1050 246 1058
rect 264 1050 276 1058
rect 294 1050 306 1058
rect 324 1050 336 1058
rect 354 1050 366 1058
rect 384 1050 396 1058
rect 414 1050 426 1058
rect 444 1050 456 1058
rect 474 1050 486 1058
rect 504 1050 516 1058
rect 534 1050 546 1058
rect 554 1050 560 1058
rect 40 1048 76 1050
rect 84 1048 106 1050
rect 114 1048 136 1050
rect 144 1048 166 1050
rect 174 1048 196 1050
rect 204 1048 226 1050
rect 234 1048 256 1050
rect 264 1048 286 1050
rect 294 1048 316 1050
rect 324 1048 346 1050
rect 354 1048 376 1050
rect 384 1048 406 1050
rect 414 1048 436 1050
rect 444 1048 466 1050
rect 474 1048 496 1050
rect 504 1048 526 1050
rect 534 1048 560 1050
rect 40 1040 56 1048
rect 64 1040 76 1048
rect 94 1040 106 1048
rect 124 1040 136 1048
rect 154 1040 166 1048
rect 184 1040 196 1048
rect 214 1040 226 1048
rect 244 1040 256 1048
rect 274 1040 286 1048
rect 304 1040 316 1048
rect 334 1040 346 1048
rect 364 1040 376 1048
rect 394 1040 406 1048
rect 424 1040 436 1048
rect 454 1040 466 1048
rect 484 1040 496 1048
rect 40 1038 76 1040
rect 40 1030 46 1038
rect 54 1030 66 1038
rect 40 1028 76 1030
rect 84 1028 506 1040
rect 40 1020 56 1028
rect 64 1020 76 1028
rect 94 1020 106 1028
rect 124 1020 136 1028
rect 154 1020 166 1028
rect 184 1020 196 1028
rect 214 1020 226 1028
rect 244 1020 256 1028
rect 274 1020 286 1028
rect 304 1020 316 1028
rect 334 1020 346 1028
rect 364 1020 376 1028
rect 394 1020 406 1028
rect 424 1020 436 1028
rect 454 1020 466 1028
rect 484 1020 496 1028
rect 514 1020 526 1048
rect 544 1040 560 1048
rect 534 1038 560 1040
rect 534 1030 546 1038
rect 554 1030 560 1038
rect 534 1028 560 1030
rect 544 1020 560 1028
rect 40 1018 76 1020
rect 84 1018 106 1020
rect 114 1018 136 1020
rect 144 1018 166 1020
rect 174 1018 196 1020
rect 204 1018 226 1020
rect 234 1018 256 1020
rect 264 1018 286 1020
rect 294 1018 316 1020
rect 324 1018 346 1020
rect 354 1018 376 1020
rect 384 1018 406 1020
rect 414 1018 436 1020
rect 444 1018 466 1020
rect 474 1018 496 1020
rect 504 1018 526 1020
rect 534 1018 560 1020
rect 40 1010 46 1018
rect 54 1010 66 1018
rect 84 1010 96 1018
rect 114 1010 126 1018
rect 144 1010 156 1018
rect 174 1010 186 1018
rect 204 1010 216 1018
rect 234 1010 246 1018
rect 264 1010 276 1018
rect 294 1010 306 1018
rect 324 1010 336 1018
rect 354 1010 366 1018
rect 384 1010 396 1018
rect 414 1010 426 1018
rect 444 1010 456 1018
rect 474 1010 486 1018
rect 504 1010 516 1018
rect 534 1010 546 1018
rect 554 1010 560 1018
rect 40 1008 76 1010
rect 84 1008 106 1010
rect 114 1008 136 1010
rect 144 1008 166 1010
rect 174 1008 196 1010
rect 204 1008 226 1010
rect 234 1008 256 1010
rect 264 1008 286 1010
rect 294 1008 316 1010
rect 324 1008 346 1010
rect 354 1008 376 1010
rect 384 1008 406 1010
rect 414 1008 436 1010
rect 444 1008 466 1010
rect 474 1008 496 1010
rect 504 1008 526 1010
rect 534 1008 560 1010
rect 40 1000 56 1008
rect 64 1000 76 1008
rect 94 1000 106 1008
rect 124 1000 136 1008
rect 154 1000 166 1008
rect 184 1000 196 1008
rect 214 1000 226 1008
rect 244 1000 256 1008
rect 274 1000 286 1008
rect 304 1000 316 1008
rect 334 1000 346 1008
rect 364 1000 376 1008
rect 394 1000 406 1008
rect 424 1000 436 1008
rect 454 1000 466 1008
rect 484 1000 496 1008
rect 514 1000 526 1008
rect 544 1000 560 1008
rect 40 998 76 1000
rect 84 998 106 1000
rect 114 998 136 1000
rect 144 998 166 1000
rect 174 998 196 1000
rect 204 998 226 1000
rect 234 998 256 1000
rect 264 998 286 1000
rect 294 998 316 1000
rect 324 998 346 1000
rect 354 998 376 1000
rect 384 998 406 1000
rect 414 998 436 1000
rect 444 998 466 1000
rect 474 998 496 1000
rect 504 998 526 1000
rect 534 998 560 1000
rect 40 990 46 998
rect 54 990 66 998
rect 84 990 96 998
rect 114 990 126 998
rect 144 990 156 998
rect 174 990 186 998
rect 204 990 216 998
rect 234 990 246 998
rect 264 990 276 998
rect 294 990 306 998
rect 324 990 336 998
rect 354 990 366 998
rect 384 990 396 998
rect 414 990 426 998
rect 444 990 456 998
rect 474 990 486 998
rect 504 990 516 998
rect 534 990 546 998
rect 554 990 560 998
rect 40 988 76 990
rect 84 988 106 990
rect 114 988 136 990
rect 144 988 166 990
rect 174 988 196 990
rect 204 988 226 990
rect 234 988 256 990
rect 264 988 286 990
rect 294 988 316 990
rect 324 988 346 990
rect 354 988 376 990
rect 384 988 406 990
rect 414 988 436 990
rect 444 988 466 990
rect 474 988 496 990
rect 504 988 526 990
rect 534 988 560 990
rect 40 980 56 988
rect 64 980 76 988
rect 94 980 106 988
rect 124 980 136 988
rect 154 980 166 988
rect 184 980 196 988
rect 214 980 226 988
rect 244 980 256 988
rect 274 980 286 988
rect 304 980 316 988
rect 334 980 346 988
rect 364 980 376 988
rect 394 980 406 988
rect 424 980 436 988
rect 454 980 466 988
rect 484 980 496 988
rect 514 980 526 988
rect 544 980 560 988
rect 40 978 76 980
rect 84 978 106 980
rect 114 978 136 980
rect 144 978 166 980
rect 174 978 196 980
rect 204 978 226 980
rect 234 978 256 980
rect 264 978 286 980
rect 294 978 316 980
rect 324 978 346 980
rect 354 978 376 980
rect 384 978 406 980
rect 414 978 436 980
rect 444 978 466 980
rect 474 978 496 980
rect 504 978 526 980
rect 534 978 560 980
rect 40 970 46 978
rect 54 970 66 978
rect 84 970 96 978
rect 114 970 126 978
rect 144 970 156 978
rect 174 970 186 978
rect 204 970 216 978
rect 234 970 246 978
rect 264 970 276 978
rect 294 970 306 978
rect 324 970 336 978
rect 354 970 366 978
rect 384 970 396 978
rect 414 970 426 978
rect 444 970 456 978
rect 474 970 486 978
rect 504 970 516 978
rect 534 970 546 978
rect 554 970 560 978
rect 40 968 560 970
rect 40 960 536 968
rect 544 960 560 968
rect 40 958 560 960
rect 40 950 46 958
rect 54 950 66 958
rect 84 950 96 958
rect 114 950 126 958
rect 144 950 156 958
rect 174 950 186 958
rect 204 950 216 958
rect 234 950 246 958
rect 264 950 276 958
rect 294 950 306 958
rect 324 950 336 958
rect 354 950 366 958
rect 384 950 396 958
rect 414 950 426 958
rect 444 950 456 958
rect 474 950 486 958
rect 504 950 516 958
rect 534 950 546 958
rect 554 950 560 958
rect 40 948 76 950
rect 84 948 106 950
rect 114 948 136 950
rect 144 948 166 950
rect 174 948 196 950
rect 204 948 226 950
rect 234 948 256 950
rect 264 948 286 950
rect 294 948 316 950
rect 324 948 346 950
rect 354 948 376 950
rect 384 948 406 950
rect 414 948 436 950
rect 444 948 466 950
rect 474 948 496 950
rect 504 948 526 950
rect 534 948 560 950
rect 40 940 56 948
rect 64 940 76 948
rect 94 940 106 948
rect 124 940 136 948
rect 154 940 166 948
rect 184 940 196 948
rect 214 940 226 948
rect 244 940 256 948
rect 274 940 286 948
rect 304 940 316 948
rect 334 940 346 948
rect 364 940 376 948
rect 394 940 406 948
rect 424 940 436 948
rect 454 940 466 948
rect 484 940 496 948
rect 514 940 526 948
rect 544 940 560 948
rect 40 938 76 940
rect 84 938 106 940
rect 114 938 136 940
rect 144 938 166 940
rect 174 938 196 940
rect 204 938 226 940
rect 234 938 256 940
rect 264 938 286 940
rect 294 938 316 940
rect 324 938 346 940
rect 354 938 376 940
rect 384 938 406 940
rect 414 938 436 940
rect 444 938 466 940
rect 474 938 496 940
rect 504 938 526 940
rect 534 938 560 940
rect 40 930 46 938
rect 54 930 66 938
rect 84 930 96 938
rect 114 930 126 938
rect 144 930 156 938
rect 174 930 186 938
rect 204 930 216 938
rect 234 930 246 938
rect 264 930 276 938
rect 294 930 306 938
rect 324 930 336 938
rect 354 930 366 938
rect 384 930 396 938
rect 414 930 426 938
rect 444 930 456 938
rect 474 930 486 938
rect 504 930 516 938
rect 534 930 546 938
rect 554 930 560 938
rect 40 928 76 930
rect 84 928 106 930
rect 114 928 136 930
rect 144 928 166 930
rect 174 928 196 930
rect 204 928 226 930
rect 234 928 256 930
rect 264 928 286 930
rect 294 928 316 930
rect 324 928 346 930
rect 354 928 376 930
rect 384 928 406 930
rect 414 928 436 930
rect 444 928 466 930
rect 474 928 496 930
rect 504 928 526 930
rect 534 928 560 930
rect 40 920 56 928
rect 64 920 76 928
rect 94 920 106 928
rect 124 920 136 928
rect 154 920 166 928
rect 184 920 196 928
rect 214 920 226 928
rect 244 920 256 928
rect 274 920 286 928
rect 304 920 316 928
rect 334 920 346 928
rect 364 920 376 928
rect 394 920 406 928
rect 424 920 436 928
rect 454 920 466 928
rect 484 920 496 928
rect 514 920 526 928
rect 544 920 560 928
rect 40 918 76 920
rect 84 918 106 920
rect 114 918 136 920
rect 144 918 166 920
rect 174 918 196 920
rect 204 918 226 920
rect 234 918 256 920
rect 264 918 286 920
rect 294 918 316 920
rect 324 918 346 920
rect 354 918 376 920
rect 384 918 406 920
rect 414 918 436 920
rect 444 918 466 920
rect 474 918 496 920
rect 504 918 526 920
rect 534 918 560 920
rect 40 910 46 918
rect 54 910 66 918
rect 84 910 96 918
rect 114 910 126 918
rect 144 910 156 918
rect 174 910 186 918
rect 204 910 216 918
rect 234 910 246 918
rect 264 910 276 918
rect 294 910 306 918
rect 324 910 336 918
rect 354 910 366 918
rect 384 910 396 918
rect 414 910 426 918
rect 444 910 456 918
rect 474 910 486 918
rect 504 910 516 918
rect 534 910 546 918
rect 554 910 560 918
rect 40 908 76 910
rect 84 908 106 910
rect 114 908 136 910
rect 144 908 166 910
rect 174 908 196 910
rect 204 908 226 910
rect 234 908 256 910
rect 264 908 286 910
rect 294 908 316 910
rect 324 908 346 910
rect 354 908 376 910
rect 384 908 406 910
rect 414 908 436 910
rect 444 908 466 910
rect 474 908 496 910
rect 504 908 526 910
rect 534 908 560 910
rect 40 900 56 908
rect 64 900 76 908
rect 94 900 106 908
rect 124 900 136 908
rect 154 900 166 908
rect 184 900 196 908
rect 214 900 226 908
rect 244 900 256 908
rect 274 900 286 908
rect 304 900 316 908
rect 334 900 346 908
rect 364 900 376 908
rect 394 900 406 908
rect 424 900 436 908
rect 454 900 466 908
rect 484 900 496 908
rect 514 900 526 908
rect 544 900 560 908
rect 40 898 76 900
rect 84 898 106 900
rect 114 898 136 900
rect 144 898 166 900
rect 174 898 196 900
rect 204 898 226 900
rect 234 898 256 900
rect 264 898 286 900
rect 294 898 316 900
rect 324 898 346 900
rect 354 898 376 900
rect 384 898 406 900
rect 414 898 436 900
rect 444 898 466 900
rect 474 898 496 900
rect 504 898 526 900
rect 534 898 560 900
rect 40 890 46 898
rect 54 890 66 898
rect 84 890 96 898
rect 114 890 126 898
rect 144 890 156 898
rect 174 890 186 898
rect 204 890 216 898
rect 234 890 246 898
rect 264 890 276 898
rect 294 890 306 898
rect 324 890 336 898
rect 354 890 366 898
rect 384 890 396 898
rect 414 890 426 898
rect 444 890 456 898
rect 474 890 486 898
rect 504 890 516 898
rect 534 890 546 898
rect 554 890 560 898
rect 40 888 76 890
rect 84 888 106 890
rect 114 888 136 890
rect 144 888 166 890
rect 174 888 196 890
rect 204 888 226 890
rect 234 888 256 890
rect 264 888 286 890
rect 294 888 316 890
rect 324 888 346 890
rect 354 888 376 890
rect 384 888 406 890
rect 414 888 436 890
rect 444 888 466 890
rect 474 888 496 890
rect 504 888 526 890
rect 534 888 560 890
rect 40 878 56 888
rect 64 878 76 888
rect 94 878 106 888
rect 124 878 136 888
rect 154 878 166 888
rect 184 878 196 888
rect 214 878 226 888
rect 244 878 256 888
rect 274 878 286 888
rect 304 878 316 888
rect 334 878 346 888
rect 364 878 376 888
rect 394 878 406 888
rect 424 878 436 888
rect 454 878 466 888
rect 484 878 496 888
rect 514 878 526 888
rect 544 878 560 888
rect 40 870 46 878
rect 554 870 560 878
rect 40 864 560 870
rect 0 652 600 654
rect 0 644 4 652
rect 12 644 24 652
rect 42 644 54 652
rect 72 644 84 652
rect 102 644 114 652
rect 132 644 144 652
rect 162 644 174 652
rect 192 644 204 652
rect 222 644 234 652
rect 242 644 256 652
rect 264 644 276 652
rect 294 644 306 652
rect 324 644 336 652
rect 344 644 358 652
rect 366 644 378 652
rect 396 644 408 652
rect 426 644 438 652
rect 456 644 468 652
rect 486 644 498 652
rect 516 644 528 652
rect 546 644 558 652
rect 576 644 588 652
rect 596 644 600 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 192 642 214 644
rect 222 642 286 644
rect 294 642 316 644
rect 324 642 378 644
rect 386 642 408 644
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 0 634 14 642
rect 22 634 34 642
rect 52 634 64 642
rect 82 634 94 642
rect 112 634 124 642
rect 142 634 154 642
rect 172 634 184 642
rect 202 634 214 642
rect 232 634 244 642
rect 252 634 266 642
rect 274 634 286 642
rect 304 634 316 642
rect 334 634 348 642
rect 356 634 368 642
rect 386 634 398 642
rect 416 634 428 642
rect 446 634 458 642
rect 476 634 488 642
rect 506 634 518 642
rect 536 634 548 642
rect 566 634 578 642
rect 586 634 600 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 192 632 214 634
rect 222 632 286 634
rect 294 632 316 634
rect 324 632 378 634
rect 386 632 408 634
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 0 624 4 632
rect 12 624 24 632
rect 42 624 54 632
rect 72 624 84 632
rect 102 624 114 632
rect 132 624 144 632
rect 162 624 174 632
rect 192 624 204 632
rect 222 624 234 632
rect 242 624 256 632
rect 264 624 276 632
rect 294 624 306 632
rect 324 624 336 632
rect 344 624 358 632
rect 366 624 378 632
rect 396 624 408 632
rect 426 624 438 632
rect 456 624 468 632
rect 486 624 498 632
rect 516 624 528 632
rect 546 624 558 632
rect 576 624 588 632
rect 596 624 600 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 192 622 214 624
rect 222 622 286 624
rect 294 622 316 624
rect 324 622 378 624
rect 386 622 408 624
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 0 614 14 622
rect 22 614 34 622
rect 52 614 64 622
rect 82 614 94 622
rect 112 614 124 622
rect 142 614 154 622
rect 172 614 184 622
rect 202 614 214 622
rect 232 614 244 622
rect 252 614 266 622
rect 274 614 286 622
rect 304 614 316 622
rect 334 614 348 622
rect 356 614 368 622
rect 386 614 398 622
rect 416 614 428 622
rect 446 614 458 622
rect 476 614 488 622
rect 506 614 518 622
rect 536 614 548 622
rect 566 614 578 622
rect 586 614 600 622
rect 0 612 214 614
rect 0 604 4 612
rect 12 604 24 612
rect 32 604 214 612
rect 0 602 214 604
rect 222 612 286 614
rect 294 612 316 614
rect 324 612 378 614
rect 222 604 234 612
rect 242 604 256 612
rect 264 604 276 612
rect 294 604 306 612
rect 324 604 336 612
rect 344 604 358 612
rect 366 604 378 612
rect 222 602 286 604
rect 294 602 316 604
rect 324 602 378 604
rect 386 612 600 614
rect 386 604 568 612
rect 576 604 588 612
rect 596 604 600 612
rect 386 602 600 604
rect 0 594 14 602
rect 22 594 34 602
rect 52 594 64 602
rect 82 594 94 602
rect 112 594 124 602
rect 142 594 154 602
rect 172 594 184 602
rect 202 594 214 602
rect 232 594 244 602
rect 252 594 266 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 192 592 214 594
rect 222 592 266 594
rect 274 592 286 602
rect 304 592 316 602
rect 334 594 348 602
rect 356 594 368 602
rect 386 594 398 602
rect 416 594 428 602
rect 446 594 458 602
rect 476 594 488 602
rect 506 594 518 602
rect 536 594 548 602
rect 566 594 578 602
rect 586 594 600 602
rect 334 592 378 594
rect 386 592 408 594
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 0 584 4 592
rect 12 584 24 592
rect 42 584 54 592
rect 72 584 84 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 592
rect 132 582 144 592
rect 162 582 174 592
rect 192 582 204 592
rect 222 582 234 592
rect 242 582 256 592
rect 0 574 14 582
rect 22 574 34 582
rect 52 574 64 582
rect 82 574 94 582
rect 252 574 256 582
rect 344 582 358 592
rect 366 582 378 592
rect 396 582 408 592
rect 426 582 438 592
rect 456 582 468 592
rect 486 582 498 592
rect 516 584 528 592
rect 546 584 558 592
rect 576 584 588 592
rect 596 584 600 592
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 344 574 348 582
rect 506 574 518 582
rect 536 574 548 582
rect 566 574 578 582
rect 586 574 600 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 0 564 4 572
rect 12 564 24 572
rect 42 564 54 572
rect 72 564 84 572
rect 102 564 114 574
rect 132 564 144 574
rect 162 564 174 574
rect 192 564 204 574
rect 222 564 234 574
rect 242 564 256 574
rect 264 564 276 574
rect 294 564 306 574
rect 324 564 336 574
rect 344 564 358 574
rect 366 564 378 574
rect 396 564 408 574
rect 426 564 438 574
rect 456 564 468 574
rect 486 564 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 516 564 528 572
rect 546 564 558 572
rect 576 564 588 572
rect 596 564 600 572
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 192 562 214 564
rect 222 562 286 564
rect 294 562 316 564
rect 324 562 378 564
rect 386 562 408 564
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 0 554 14 562
rect 22 554 34 562
rect 52 554 64 562
rect 82 554 94 562
rect 112 554 124 562
rect 142 554 154 562
rect 172 554 184 562
rect 202 554 214 562
rect 232 554 244 562
rect 252 554 266 562
rect 274 554 286 562
rect 304 554 316 562
rect 334 554 348 562
rect 356 554 368 562
rect 386 554 398 562
rect 416 554 428 562
rect 446 554 458 562
rect 476 554 488 562
rect 506 554 518 562
rect 536 554 548 562
rect 566 554 578 562
rect 586 554 600 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 192 552 214 554
rect 222 552 286 554
rect 294 552 316 554
rect 324 552 378 554
rect 386 552 408 554
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 0 544 4 552
rect 12 544 24 552
rect 42 544 54 552
rect 72 544 84 552
rect 102 544 114 552
rect 132 544 144 552
rect 162 544 174 552
rect 192 544 204 552
rect 222 544 234 552
rect 242 544 256 552
rect 264 544 276 552
rect 294 544 306 552
rect 324 544 336 552
rect 344 544 358 552
rect 366 544 378 552
rect 396 544 408 552
rect 426 544 438 552
rect 456 544 468 552
rect 486 544 498 552
rect 516 544 528 552
rect 546 544 558 552
rect 576 544 588 552
rect 596 544 600 552
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 192 542 214 544
rect 222 542 286 544
rect 294 542 316 544
rect 324 542 378 544
rect 386 542 408 544
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 0 534 14 542
rect 22 534 34 542
rect 52 534 64 542
rect 82 534 94 542
rect 112 534 124 542
rect 142 534 154 542
rect 172 534 184 542
rect 202 534 214 542
rect 232 534 244 542
rect 252 534 266 542
rect 274 534 286 542
rect 304 534 316 542
rect 334 534 348 542
rect 356 534 368 542
rect 386 534 398 542
rect 416 534 428 542
rect 446 534 458 542
rect 476 534 488 542
rect 506 534 518 542
rect 536 534 548 542
rect 566 534 578 542
rect 586 534 600 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 192 532 214 534
rect 222 532 286 534
rect 294 532 316 534
rect 324 532 378 534
rect 386 532 408 534
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 0 524 4 532
rect 12 524 24 532
rect 42 524 54 532
rect 72 524 84 532
rect 102 524 114 532
rect 132 524 144 532
rect 162 524 174 532
rect 192 524 204 532
rect 222 524 234 532
rect 242 524 256 532
rect 264 524 276 532
rect 294 524 306 532
rect 324 524 336 532
rect 344 524 358 532
rect 366 524 378 532
rect 396 524 408 532
rect 426 524 438 532
rect 456 524 468 532
rect 486 524 498 532
rect 516 524 528 532
rect 546 524 558 532
rect 576 524 588 532
rect 596 524 600 532
rect 0 516 600 524
rect 0 512 24 516
rect 0 4 4 512
rect 12 508 24 512
rect 32 508 44 516
rect 52 508 64 516
rect 72 508 84 516
rect 92 508 104 516
rect 112 508 124 516
rect 132 508 144 516
rect 152 508 164 516
rect 172 508 184 516
rect 192 508 204 516
rect 212 508 224 516
rect 232 508 244 516
rect 252 508 264 516
rect 272 508 284 516
rect 292 508 318 516
rect 326 508 338 516
rect 346 508 358 516
rect 366 508 378 516
rect 386 508 398 516
rect 406 508 418 516
rect 426 508 438 516
rect 446 508 458 516
rect 466 508 478 516
rect 486 508 498 516
rect 506 508 518 516
rect 526 508 538 516
rect 546 508 558 516
rect 566 508 578 516
rect 586 512 600 516
rect 12 504 588 508
rect 12 16 16 504
rect 584 16 588 504
rect 12 12 588 16
rect 12 4 16 12
rect 584 4 588 12
rect 596 4 600 512
rect 0 0 600 4
<< psubstratepcontact >>
rect 4 1328 332 1336
rect 338 1328 596 1336
rect 4 828 12 1328
rect 24 828 42 836
rect 54 828 72 836
rect 84 828 102 836
rect 114 828 132 836
rect 144 828 162 836
rect 174 828 192 836
rect 204 828 222 836
rect 234 828 242 836
rect 256 828 264 836
rect 276 828 294 836
rect 306 828 324 836
rect 336 828 344 836
rect 358 828 366 836
rect 378 828 396 836
rect 408 828 426 836
rect 438 828 456 836
rect 468 828 486 836
rect 498 828 516 836
rect 528 828 546 836
rect 558 828 576 836
rect 588 828 596 1328
rect 34 826 42 828
rect 64 826 72 828
rect 94 826 102 828
rect 124 826 132 828
rect 154 826 162 828
rect 184 826 192 828
rect 214 826 222 828
rect 286 826 294 828
rect 316 826 324 828
rect 378 826 386 828
rect 408 826 416 828
rect 438 826 446 828
rect 468 826 476 828
rect 498 826 506 828
rect 528 826 536 828
rect 558 826 566 828
rect 14 818 22 826
rect 34 818 52 826
rect 64 818 82 826
rect 94 818 112 826
rect 124 818 142 826
rect 154 818 172 826
rect 184 818 202 826
rect 214 818 232 826
rect 244 818 252 826
rect 266 818 274 826
rect 286 818 304 826
rect 316 818 334 826
rect 348 818 356 826
rect 368 818 386 826
rect 398 818 416 826
rect 428 818 446 826
rect 458 818 476 826
rect 488 818 506 826
rect 518 818 536 826
rect 548 818 566 826
rect 578 818 586 826
rect 34 816 42 818
rect 64 816 72 818
rect 94 816 102 818
rect 124 816 132 818
rect 154 816 162 818
rect 184 816 192 818
rect 214 816 222 818
rect 286 816 294 818
rect 316 816 324 818
rect 378 816 386 818
rect 408 816 416 818
rect 438 816 446 818
rect 468 816 476 818
rect 498 816 506 818
rect 528 816 536 818
rect 558 816 566 818
rect 4 808 12 816
rect 24 808 42 816
rect 54 808 72 816
rect 84 808 102 816
rect 114 808 132 816
rect 144 808 162 816
rect 174 808 192 816
rect 204 808 222 816
rect 234 808 242 816
rect 256 808 264 816
rect 276 808 294 816
rect 306 808 324 816
rect 336 808 344 816
rect 358 808 366 816
rect 378 808 396 816
rect 408 808 426 816
rect 438 808 456 816
rect 468 808 486 816
rect 498 808 516 816
rect 528 808 546 816
rect 558 808 576 816
rect 588 808 596 816
rect 34 806 42 808
rect 64 806 72 808
rect 94 806 102 808
rect 124 806 132 808
rect 154 806 162 808
rect 184 806 192 808
rect 214 806 222 808
rect 286 806 294 808
rect 316 806 324 808
rect 378 806 386 808
rect 408 806 416 808
rect 438 806 446 808
rect 468 806 476 808
rect 498 806 506 808
rect 528 806 536 808
rect 558 806 566 808
rect 14 798 22 806
rect 34 798 52 806
rect 64 798 82 806
rect 94 798 112 806
rect 124 798 142 806
rect 154 798 172 806
rect 184 798 202 806
rect 214 798 232 806
rect 244 798 252 806
rect 266 798 274 806
rect 286 798 304 806
rect 316 798 334 806
rect 348 798 356 806
rect 368 798 386 806
rect 398 798 416 806
rect 428 798 446 806
rect 458 798 476 806
rect 488 798 506 806
rect 518 798 536 806
rect 548 798 566 806
rect 578 798 586 806
rect 34 796 42 798
rect 64 796 72 798
rect 94 796 102 798
rect 124 796 132 798
rect 154 796 162 798
rect 184 796 192 798
rect 214 796 222 798
rect 286 796 294 798
rect 316 796 324 798
rect 378 796 386 798
rect 408 796 416 798
rect 438 796 446 798
rect 468 796 476 798
rect 498 796 506 798
rect 528 796 536 798
rect 558 796 566 798
rect 4 788 12 796
rect 24 788 42 796
rect 54 788 72 796
rect 84 788 102 796
rect 114 788 132 796
rect 144 788 162 796
rect 174 788 192 796
rect 204 788 222 796
rect 234 788 242 796
rect 256 788 264 796
rect 276 788 294 796
rect 306 788 324 796
rect 336 788 344 796
rect 358 788 366 796
rect 378 788 396 796
rect 408 788 426 796
rect 438 788 456 796
rect 468 788 486 796
rect 498 788 516 796
rect 528 788 546 796
rect 558 788 576 796
rect 588 788 596 796
rect 34 786 42 788
rect 64 786 72 788
rect 94 786 102 788
rect 124 786 132 788
rect 154 786 162 788
rect 184 786 192 788
rect 214 786 222 788
rect 286 786 294 788
rect 316 786 324 788
rect 378 786 386 788
rect 408 786 416 788
rect 438 786 446 788
rect 468 786 476 788
rect 498 786 506 788
rect 528 786 536 788
rect 558 786 566 788
rect 14 778 22 786
rect 34 778 52 786
rect 64 778 82 786
rect 34 776 42 778
rect 64 776 72 778
rect 94 776 112 786
rect 124 776 142 786
rect 154 776 172 786
rect 184 776 202 786
rect 214 776 232 786
rect 244 776 252 786
rect 266 776 274 786
rect 286 776 304 786
rect 316 776 334 786
rect 348 776 356 786
rect 368 776 386 786
rect 398 776 416 786
rect 428 776 446 786
rect 458 776 476 786
rect 488 776 506 786
rect 518 778 536 786
rect 548 778 566 786
rect 578 778 586 786
rect 528 776 536 778
rect 558 776 566 778
rect 4 768 12 776
rect 24 768 42 776
rect 54 768 72 776
rect 84 768 252 776
rect 256 768 344 776
rect 348 768 516 776
rect 528 768 546 776
rect 558 768 576 776
rect 588 768 596 776
rect 34 766 42 768
rect 64 766 72 768
rect 14 758 22 766
rect 34 758 52 766
rect 64 758 82 766
rect 94 758 112 768
rect 124 758 142 768
rect 154 758 172 768
rect 184 758 202 768
rect 214 758 232 768
rect 244 758 252 768
rect 266 758 274 768
rect 286 758 304 768
rect 316 758 334 768
rect 348 758 356 768
rect 368 758 386 768
rect 398 758 416 768
rect 428 758 446 768
rect 458 758 476 768
rect 488 758 506 768
rect 528 766 536 768
rect 558 766 566 768
rect 518 758 536 766
rect 548 758 566 766
rect 578 758 586 766
rect 34 756 42 758
rect 64 756 72 758
rect 94 756 102 758
rect 124 756 132 758
rect 154 756 162 758
rect 184 756 192 758
rect 214 756 222 758
rect 286 756 294 758
rect 316 756 324 758
rect 378 756 386 758
rect 408 756 416 758
rect 438 756 446 758
rect 468 756 476 758
rect 498 756 506 758
rect 528 756 536 758
rect 558 756 566 758
rect 4 748 12 756
rect 24 748 42 756
rect 54 748 72 756
rect 84 748 102 756
rect 114 748 132 756
rect 144 748 162 756
rect 174 748 192 756
rect 204 748 222 756
rect 234 748 242 756
rect 256 748 264 756
rect 276 748 294 756
rect 306 748 324 756
rect 336 748 344 756
rect 358 748 366 756
rect 378 748 396 756
rect 408 748 426 756
rect 438 748 456 756
rect 468 748 486 756
rect 498 748 516 756
rect 528 748 546 756
rect 558 748 576 756
rect 588 748 596 756
rect 34 746 42 748
rect 64 746 72 748
rect 94 746 102 748
rect 124 746 132 748
rect 154 746 162 748
rect 184 746 192 748
rect 214 746 222 748
rect 286 746 294 748
rect 316 746 324 748
rect 378 746 386 748
rect 408 746 416 748
rect 438 746 446 748
rect 468 746 476 748
rect 498 746 506 748
rect 528 746 536 748
rect 558 746 566 748
rect 14 738 22 746
rect 34 738 52 746
rect 64 738 82 746
rect 94 738 112 746
rect 124 738 142 746
rect 154 738 172 746
rect 184 738 202 746
rect 214 738 232 746
rect 244 738 252 746
rect 266 738 274 746
rect 286 738 304 746
rect 316 738 334 746
rect 348 738 356 746
rect 368 738 386 746
rect 398 738 416 746
rect 428 738 446 746
rect 458 738 476 746
rect 488 738 506 746
rect 518 738 536 746
rect 548 738 566 746
rect 578 738 586 746
rect 4 728 12 736
rect 24 728 32 736
rect 214 726 222 738
rect 286 736 294 738
rect 316 736 324 738
rect 234 728 242 736
rect 256 728 264 736
rect 276 728 294 736
rect 306 728 324 736
rect 336 728 344 736
rect 358 728 366 736
rect 286 726 294 728
rect 316 726 324 728
rect 378 726 386 738
rect 568 728 576 736
rect 588 728 596 736
rect 14 718 22 726
rect 34 718 52 726
rect 64 718 82 726
rect 94 718 112 726
rect 124 718 142 726
rect 154 718 172 726
rect 184 718 202 726
rect 214 718 232 726
rect 244 718 252 726
rect 266 718 274 726
rect 286 718 304 726
rect 316 718 334 726
rect 348 718 356 726
rect 368 718 386 726
rect 398 718 416 726
rect 428 718 446 726
rect 458 718 476 726
rect 488 718 506 726
rect 518 718 536 726
rect 548 718 566 726
rect 578 718 586 726
rect 34 716 42 718
rect 64 716 72 718
rect 94 716 102 718
rect 124 716 132 718
rect 154 716 162 718
rect 184 716 192 718
rect 214 716 222 718
rect 286 716 294 718
rect 316 716 324 718
rect 378 716 386 718
rect 408 716 416 718
rect 438 716 446 718
rect 468 716 476 718
rect 498 716 506 718
rect 528 716 536 718
rect 558 716 566 718
rect 4 708 12 716
rect 24 708 42 716
rect 54 708 72 716
rect 84 708 102 716
rect 114 708 132 716
rect 144 708 162 716
rect 174 708 192 716
rect 204 708 222 716
rect 234 708 242 716
rect 256 708 264 716
rect 276 708 294 716
rect 306 708 324 716
rect 336 708 344 716
rect 358 708 366 716
rect 378 708 396 716
rect 408 708 426 716
rect 438 708 456 716
rect 468 708 486 716
rect 498 708 516 716
rect 528 708 546 716
rect 558 708 576 716
rect 588 708 596 716
rect 34 706 42 708
rect 64 706 72 708
rect 94 706 102 708
rect 124 706 132 708
rect 154 706 162 708
rect 184 706 192 708
rect 214 706 222 708
rect 286 706 294 708
rect 316 706 324 708
rect 378 706 386 708
rect 408 706 416 708
rect 438 706 446 708
rect 468 706 476 708
rect 498 706 506 708
rect 528 706 536 708
rect 558 706 566 708
rect 14 698 22 706
rect 34 698 52 706
rect 64 698 82 706
rect 94 698 112 706
rect 124 698 142 706
rect 154 698 172 706
rect 184 698 202 706
rect 214 698 232 706
rect 244 698 252 706
rect 266 698 274 706
rect 286 698 304 706
rect 316 698 334 706
rect 348 698 356 706
rect 368 698 386 706
rect 398 698 416 706
rect 428 698 446 706
rect 458 698 476 706
rect 488 698 506 706
rect 518 698 536 706
rect 548 698 566 706
rect 578 698 586 706
rect 34 696 42 698
rect 64 696 72 698
rect 94 696 102 698
rect 124 696 132 698
rect 154 696 162 698
rect 184 696 192 698
rect 214 696 222 698
rect 286 696 294 698
rect 316 696 324 698
rect 378 696 386 698
rect 408 696 416 698
rect 438 696 446 698
rect 468 696 476 698
rect 498 696 506 698
rect 528 696 536 698
rect 558 696 566 698
rect 4 688 12 696
rect 24 688 42 696
rect 54 688 72 696
rect 84 688 102 696
rect 114 688 132 696
rect 144 688 162 696
rect 174 688 192 696
rect 204 688 222 696
rect 234 688 242 696
rect 256 688 264 696
rect 276 688 294 696
rect 306 688 324 696
rect 336 688 344 696
rect 358 688 366 696
rect 378 688 396 696
rect 408 688 426 696
rect 438 688 456 696
rect 468 688 486 696
rect 498 688 516 696
rect 528 688 546 696
rect 558 688 576 696
rect 588 688 596 696
rect 32 460 570 488
rect 42 450 50 460
rect 62 450 80 460
rect 92 450 110 460
rect 122 450 140 460
rect 152 450 170 460
rect 182 450 200 460
rect 212 450 230 460
rect 242 450 260 460
rect 272 450 290 460
rect 302 450 320 460
rect 332 450 350 460
rect 362 450 380 460
rect 392 450 410 460
rect 422 450 440 460
rect 452 450 470 460
rect 482 450 500 460
rect 512 450 530 460
rect 542 450 560 460
rect 62 448 70 450
rect 92 448 100 450
rect 122 448 130 450
rect 152 448 160 450
rect 182 448 190 450
rect 212 448 220 450
rect 242 448 250 450
rect 272 448 280 450
rect 302 448 310 450
rect 332 448 340 450
rect 362 448 370 450
rect 392 448 400 450
rect 422 448 430 450
rect 452 448 460 450
rect 482 448 490 450
rect 512 448 520 450
rect 542 448 550 450
rect 32 440 40 448
rect 52 440 70 448
rect 82 440 100 448
rect 112 440 130 448
rect 142 440 160 448
rect 172 440 190 448
rect 202 440 220 448
rect 232 440 250 448
rect 262 440 280 448
rect 292 440 310 448
rect 322 440 340 448
rect 352 440 370 448
rect 382 440 400 448
rect 412 440 430 448
rect 442 440 460 448
rect 472 440 490 448
rect 502 440 520 448
rect 532 440 550 448
rect 562 440 570 448
rect 62 438 70 440
rect 92 438 100 440
rect 122 438 130 440
rect 152 438 160 440
rect 182 438 190 440
rect 212 438 220 440
rect 242 438 250 440
rect 272 438 280 440
rect 302 438 310 440
rect 332 438 340 440
rect 362 438 370 440
rect 392 438 400 440
rect 422 438 430 440
rect 452 438 460 440
rect 482 438 490 440
rect 512 438 520 440
rect 542 438 550 440
rect 42 430 50 438
rect 62 430 80 438
rect 92 430 110 438
rect 122 430 140 438
rect 152 430 170 438
rect 182 430 200 438
rect 212 430 230 438
rect 242 430 260 438
rect 272 430 290 438
rect 302 430 320 438
rect 332 430 350 438
rect 362 430 380 438
rect 392 430 410 438
rect 422 430 440 438
rect 452 430 470 438
rect 482 430 500 438
rect 512 430 530 438
rect 542 430 560 438
rect 62 428 70 430
rect 92 428 100 430
rect 122 428 130 430
rect 152 428 160 430
rect 182 428 190 430
rect 212 428 220 430
rect 242 428 250 430
rect 272 428 280 430
rect 302 428 310 430
rect 332 428 340 430
rect 362 428 370 430
rect 392 428 400 430
rect 422 428 430 430
rect 452 428 460 430
rect 482 428 490 430
rect 512 428 520 430
rect 542 428 550 430
rect 32 420 40 428
rect 52 420 70 428
rect 82 420 100 428
rect 112 420 130 428
rect 142 420 160 428
rect 172 420 190 428
rect 202 420 220 428
rect 232 420 250 428
rect 262 420 280 428
rect 292 420 310 428
rect 322 420 340 428
rect 352 420 370 428
rect 382 420 400 428
rect 412 420 430 428
rect 442 420 460 428
rect 472 420 490 428
rect 502 420 520 428
rect 532 420 550 428
rect 562 420 570 428
rect 62 418 70 420
rect 92 418 100 420
rect 122 418 130 420
rect 152 418 160 420
rect 182 418 190 420
rect 212 418 220 420
rect 242 418 250 420
rect 272 418 280 420
rect 302 418 310 420
rect 332 418 340 420
rect 362 418 370 420
rect 392 418 400 420
rect 422 418 430 420
rect 452 418 460 420
rect 482 418 490 420
rect 512 418 520 420
rect 542 418 550 420
rect 42 410 50 418
rect 62 410 80 418
rect 92 410 110 418
rect 122 410 140 418
rect 152 410 170 418
rect 182 410 200 418
rect 212 410 230 418
rect 242 410 260 418
rect 272 410 290 418
rect 302 410 320 418
rect 332 410 350 418
rect 362 410 380 418
rect 392 410 410 418
rect 422 410 440 418
rect 452 410 470 418
rect 482 410 500 418
rect 512 410 530 418
rect 542 410 560 418
rect 62 408 70 410
rect 92 408 100 410
rect 122 408 130 410
rect 152 408 160 410
rect 182 408 190 410
rect 212 408 220 410
rect 242 408 250 410
rect 272 408 280 410
rect 302 408 310 410
rect 332 408 340 410
rect 362 408 370 410
rect 392 408 400 410
rect 422 408 430 410
rect 452 408 460 410
rect 482 408 490 410
rect 512 408 520 410
rect 542 408 550 410
rect 32 400 40 408
rect 52 400 70 408
rect 82 400 100 408
rect 112 400 130 408
rect 142 400 160 408
rect 172 400 190 408
rect 202 400 220 408
rect 232 400 250 408
rect 262 400 280 408
rect 292 400 310 408
rect 322 400 340 408
rect 352 400 370 408
rect 382 400 400 408
rect 412 400 430 408
rect 442 400 460 408
rect 472 400 490 408
rect 502 400 520 408
rect 532 400 550 408
rect 562 400 570 408
rect 62 398 70 400
rect 92 398 100 400
rect 122 398 130 400
rect 152 398 160 400
rect 182 398 190 400
rect 212 398 220 400
rect 242 398 250 400
rect 272 398 280 400
rect 302 398 310 400
rect 332 398 340 400
rect 362 398 370 400
rect 392 398 400 400
rect 422 398 430 400
rect 452 398 460 400
rect 482 398 490 400
rect 512 398 520 400
rect 542 398 550 400
rect 42 370 50 398
rect 62 370 80 398
rect 92 390 110 398
rect 122 390 140 398
rect 152 390 170 398
rect 182 390 200 398
rect 212 390 230 398
rect 242 390 260 398
rect 272 390 290 398
rect 302 390 320 398
rect 332 390 350 398
rect 362 390 380 398
rect 392 390 410 398
rect 422 390 440 398
rect 452 390 470 398
rect 482 390 500 398
rect 512 390 530 398
rect 542 390 560 398
rect 92 378 100 390
rect 512 378 520 390
rect 542 388 550 390
rect 532 380 550 388
rect 562 380 570 388
rect 542 378 550 380
rect 92 370 110 378
rect 122 370 140 378
rect 152 370 170 378
rect 182 370 200 378
rect 212 370 230 378
rect 242 370 260 378
rect 272 370 290 378
rect 302 370 320 378
rect 332 370 350 378
rect 362 370 380 378
rect 392 370 410 378
rect 422 370 440 378
rect 452 370 470 378
rect 482 370 500 378
rect 512 370 530 378
rect 542 370 560 378
rect 62 368 70 370
rect 92 368 100 370
rect 122 368 130 370
rect 152 368 160 370
rect 182 368 190 370
rect 212 368 220 370
rect 242 368 250 370
rect 272 368 280 370
rect 302 368 310 370
rect 332 368 340 370
rect 362 368 370 370
rect 392 368 400 370
rect 422 368 430 370
rect 452 368 460 370
rect 482 368 490 370
rect 512 368 520 370
rect 542 368 550 370
rect 32 360 40 368
rect 52 360 70 368
rect 82 360 100 368
rect 112 360 130 368
rect 142 360 160 368
rect 172 360 190 368
rect 202 360 220 368
rect 232 360 250 368
rect 262 360 280 368
rect 292 360 310 368
rect 322 360 340 368
rect 352 360 370 368
rect 382 360 400 368
rect 412 360 430 368
rect 442 360 460 368
rect 472 360 490 368
rect 502 360 520 368
rect 532 360 550 368
rect 562 360 570 368
rect 62 358 70 360
rect 92 358 100 360
rect 122 358 130 360
rect 152 358 160 360
rect 182 358 190 360
rect 212 358 220 360
rect 242 358 250 360
rect 272 358 280 360
rect 302 358 310 360
rect 332 358 340 360
rect 362 358 370 360
rect 392 358 400 360
rect 422 358 430 360
rect 452 358 460 360
rect 482 358 490 360
rect 512 358 520 360
rect 542 358 550 360
rect 42 350 50 358
rect 62 350 80 358
rect 92 350 110 358
rect 122 350 140 358
rect 152 350 170 358
rect 182 350 200 358
rect 212 350 230 358
rect 242 350 260 358
rect 272 350 290 358
rect 302 350 320 358
rect 332 350 350 358
rect 362 350 380 358
rect 392 350 410 358
rect 422 350 440 358
rect 452 350 470 358
rect 482 350 500 358
rect 512 350 530 358
rect 542 350 560 358
rect 62 348 70 350
rect 92 348 100 350
rect 122 348 130 350
rect 152 348 160 350
rect 182 348 190 350
rect 212 348 220 350
rect 242 348 250 350
rect 272 348 280 350
rect 302 348 310 350
rect 332 348 340 350
rect 362 348 370 350
rect 392 348 400 350
rect 422 348 430 350
rect 452 348 460 350
rect 482 348 490 350
rect 512 348 520 350
rect 542 348 550 350
rect 32 340 40 348
rect 52 340 70 348
rect 82 340 100 348
rect 112 340 130 348
rect 142 340 160 348
rect 172 340 190 348
rect 202 340 220 348
rect 232 340 250 348
rect 262 340 280 348
rect 292 340 310 348
rect 322 340 340 348
rect 352 340 370 348
rect 382 340 400 348
rect 412 340 430 348
rect 442 340 460 348
rect 472 340 490 348
rect 502 340 520 348
rect 532 340 550 348
rect 562 340 570 348
rect 62 338 70 340
rect 92 338 100 340
rect 122 338 130 340
rect 152 338 160 340
rect 182 338 190 340
rect 212 338 220 340
rect 242 338 250 340
rect 272 338 280 340
rect 302 338 310 340
rect 332 338 340 340
rect 362 338 370 340
rect 392 338 400 340
rect 422 338 430 340
rect 452 338 460 340
rect 482 338 490 340
rect 512 338 520 340
rect 542 338 550 340
rect 42 330 50 338
rect 62 330 80 338
rect 92 330 110 338
rect 122 330 140 338
rect 152 330 170 338
rect 182 330 200 338
rect 212 330 230 338
rect 242 330 260 338
rect 272 330 290 338
rect 302 330 320 338
rect 332 330 350 338
rect 362 330 380 338
rect 392 330 410 338
rect 422 330 440 338
rect 452 330 470 338
rect 482 330 500 338
rect 512 330 530 338
rect 542 330 560 338
rect 62 328 70 330
rect 92 328 100 330
rect 122 328 130 330
rect 152 328 160 330
rect 182 328 190 330
rect 212 328 220 330
rect 242 328 250 330
rect 272 328 280 330
rect 302 328 310 330
rect 332 328 340 330
rect 362 328 370 330
rect 392 328 400 330
rect 422 328 430 330
rect 452 328 460 330
rect 482 328 490 330
rect 512 328 520 330
rect 542 328 550 330
rect 32 320 40 328
rect 52 320 70 328
rect 82 320 100 328
rect 112 320 130 328
rect 142 320 160 328
rect 172 320 190 328
rect 202 320 220 328
rect 232 320 250 328
rect 262 320 280 328
rect 292 320 310 328
rect 322 320 340 328
rect 352 320 370 328
rect 382 320 400 328
rect 412 320 430 328
rect 442 320 460 328
rect 472 320 490 328
rect 502 320 520 328
rect 532 320 550 328
rect 562 320 570 328
rect 62 318 70 320
rect 92 318 100 320
rect 122 318 130 320
rect 152 318 160 320
rect 182 318 190 320
rect 212 318 220 320
rect 242 318 250 320
rect 272 318 280 320
rect 302 318 310 320
rect 332 318 340 320
rect 362 318 370 320
rect 392 318 400 320
rect 422 318 430 320
rect 452 318 460 320
rect 482 318 490 320
rect 512 318 520 320
rect 542 318 550 320
rect 42 310 50 318
rect 62 310 80 318
rect 92 310 110 318
rect 122 310 140 318
rect 152 310 170 318
rect 182 310 200 318
rect 212 310 230 318
rect 242 310 260 318
rect 272 310 290 318
rect 302 310 320 318
rect 332 310 350 318
rect 362 310 380 318
rect 392 310 410 318
rect 422 310 440 318
rect 452 310 470 318
rect 482 310 500 318
rect 512 310 530 318
rect 542 310 560 318
rect 62 308 70 310
rect 512 308 520 310
rect 542 308 550 310
rect 32 300 40 308
rect 52 300 70 308
rect 82 300 90 308
rect 502 300 520 308
rect 532 300 550 308
rect 562 300 570 308
rect 62 298 70 300
rect 512 298 520 300
rect 542 298 550 300
rect 42 290 50 298
rect 62 290 80 298
rect 92 290 110 298
rect 122 290 140 298
rect 152 290 170 298
rect 182 290 200 298
rect 212 290 230 298
rect 242 290 260 298
rect 272 290 290 298
rect 302 290 320 298
rect 332 290 350 298
rect 362 290 380 298
rect 392 290 410 298
rect 422 290 440 298
rect 452 290 470 298
rect 482 290 500 298
rect 512 290 530 298
rect 542 290 560 298
rect 62 288 70 290
rect 92 288 100 290
rect 122 288 130 290
rect 152 288 160 290
rect 182 288 190 290
rect 212 288 220 290
rect 242 288 250 290
rect 272 288 280 290
rect 302 288 310 290
rect 332 288 340 290
rect 362 288 370 290
rect 392 288 400 290
rect 422 288 430 290
rect 452 288 460 290
rect 482 288 490 290
rect 512 288 520 290
rect 542 288 550 290
rect 32 280 40 288
rect 52 280 70 288
rect 82 280 100 288
rect 112 280 130 288
rect 142 280 160 288
rect 172 280 190 288
rect 202 280 220 288
rect 232 280 250 288
rect 262 280 280 288
rect 292 280 310 288
rect 322 280 340 288
rect 352 280 370 288
rect 382 280 400 288
rect 412 280 430 288
rect 442 280 460 288
rect 472 280 490 288
rect 502 280 520 288
rect 532 280 550 288
rect 562 280 570 288
rect 62 278 70 280
rect 92 278 100 280
rect 122 278 130 280
rect 152 278 160 280
rect 182 278 190 280
rect 212 278 220 280
rect 242 278 250 280
rect 272 278 280 280
rect 302 278 310 280
rect 332 278 340 280
rect 362 278 370 280
rect 392 278 400 280
rect 422 278 430 280
rect 452 278 460 280
rect 482 278 490 280
rect 512 278 520 280
rect 542 278 550 280
rect 42 270 50 278
rect 62 270 80 278
rect 92 270 110 278
rect 122 270 140 278
rect 152 270 170 278
rect 182 270 200 278
rect 212 270 230 278
rect 242 270 260 278
rect 272 270 290 278
rect 302 270 320 278
rect 332 270 350 278
rect 362 270 380 278
rect 392 270 410 278
rect 422 270 440 278
rect 452 270 470 278
rect 482 270 500 278
rect 512 270 530 278
rect 542 270 560 278
rect 62 268 70 270
rect 92 268 100 270
rect 122 268 130 270
rect 152 268 160 270
rect 182 268 190 270
rect 212 268 220 270
rect 242 268 250 270
rect 272 268 280 270
rect 302 268 310 270
rect 332 268 340 270
rect 362 268 370 270
rect 392 268 400 270
rect 422 268 430 270
rect 452 268 460 270
rect 482 268 490 270
rect 512 268 520 270
rect 542 268 550 270
rect 32 260 40 268
rect 52 260 70 268
rect 82 260 100 268
rect 112 260 130 268
rect 142 260 160 268
rect 172 260 190 268
rect 202 260 220 268
rect 232 260 250 268
rect 262 260 280 268
rect 292 260 310 268
rect 322 260 340 268
rect 352 260 370 268
rect 382 260 400 268
rect 412 260 430 268
rect 442 260 460 268
rect 472 260 490 268
rect 502 260 520 268
rect 532 260 550 268
rect 562 260 570 268
rect 62 258 70 260
rect 92 258 100 260
rect 122 258 130 260
rect 152 258 160 260
rect 182 258 190 260
rect 212 258 220 260
rect 242 258 250 260
rect 272 258 280 260
rect 302 258 310 260
rect 332 258 340 260
rect 362 258 370 260
rect 392 258 400 260
rect 422 258 430 260
rect 452 258 460 260
rect 482 258 490 260
rect 512 258 520 260
rect 542 258 550 260
rect 42 250 50 258
rect 62 250 80 258
rect 92 250 110 258
rect 122 250 140 258
rect 152 250 170 258
rect 182 250 200 258
rect 212 250 230 258
rect 242 250 260 258
rect 272 250 290 258
rect 302 250 320 258
rect 332 250 350 258
rect 362 250 380 258
rect 392 250 410 258
rect 422 250 440 258
rect 452 250 470 258
rect 482 250 500 258
rect 512 250 530 258
rect 542 250 560 258
rect 62 248 70 250
rect 92 248 100 250
rect 122 248 130 250
rect 152 248 160 250
rect 182 248 190 250
rect 212 248 220 250
rect 242 248 250 250
rect 272 248 280 250
rect 302 248 310 250
rect 332 248 340 250
rect 362 248 370 250
rect 392 248 400 250
rect 422 248 430 250
rect 452 248 460 250
rect 482 248 490 250
rect 512 248 520 250
rect 542 248 550 250
rect 32 240 40 248
rect 52 240 70 248
rect 42 230 50 238
rect 62 228 70 240
rect 32 220 40 228
rect 52 220 70 228
rect 82 240 100 248
rect 112 240 130 248
rect 142 240 160 248
rect 172 240 190 248
rect 202 240 220 248
rect 232 240 250 248
rect 262 240 280 248
rect 292 240 310 248
rect 322 240 340 248
rect 352 240 370 248
rect 382 240 400 248
rect 412 240 430 248
rect 442 240 460 248
rect 472 240 490 248
rect 502 240 520 248
rect 532 240 550 248
rect 562 240 570 248
rect 82 228 90 240
rect 502 228 510 240
rect 542 238 550 240
rect 522 230 530 238
rect 542 230 560 238
rect 542 228 550 230
rect 82 220 100 228
rect 112 220 130 228
rect 142 220 160 228
rect 172 220 190 228
rect 202 220 220 228
rect 232 220 250 228
rect 262 220 280 228
rect 292 220 310 228
rect 322 220 340 228
rect 352 220 370 228
rect 382 220 400 228
rect 412 220 430 228
rect 442 220 460 228
rect 472 220 490 228
rect 502 220 520 228
rect 532 220 550 228
rect 562 220 570 228
rect 62 218 70 220
rect 92 218 100 220
rect 122 218 130 220
rect 152 218 160 220
rect 182 218 190 220
rect 212 218 220 220
rect 242 218 250 220
rect 272 218 280 220
rect 302 218 310 220
rect 332 218 340 220
rect 362 218 370 220
rect 392 218 400 220
rect 422 218 430 220
rect 452 218 460 220
rect 482 218 490 220
rect 512 218 520 220
rect 542 218 550 220
rect 42 210 50 218
rect 62 210 80 218
rect 92 210 110 218
rect 122 210 140 218
rect 152 210 170 218
rect 182 210 200 218
rect 212 210 230 218
rect 242 210 260 218
rect 272 210 290 218
rect 302 210 320 218
rect 332 210 350 218
rect 362 210 380 218
rect 392 210 410 218
rect 422 210 440 218
rect 452 210 470 218
rect 482 210 500 218
rect 512 210 530 218
rect 542 210 560 218
rect 62 208 70 210
rect 92 208 100 210
rect 122 208 130 210
rect 152 208 160 210
rect 182 208 190 210
rect 212 208 220 210
rect 242 208 250 210
rect 272 208 280 210
rect 302 208 310 210
rect 332 208 340 210
rect 362 208 370 210
rect 392 208 400 210
rect 422 208 430 210
rect 452 208 460 210
rect 482 208 490 210
rect 512 208 520 210
rect 542 208 550 210
rect 32 200 40 208
rect 52 200 70 208
rect 82 200 100 208
rect 112 200 130 208
rect 142 200 160 208
rect 172 200 190 208
rect 202 200 220 208
rect 232 200 250 208
rect 262 200 280 208
rect 292 200 310 208
rect 322 200 340 208
rect 352 200 370 208
rect 382 200 400 208
rect 412 200 430 208
rect 442 200 460 208
rect 472 200 490 208
rect 502 200 520 208
rect 532 200 550 208
rect 562 200 570 208
rect 62 198 70 200
rect 92 198 100 200
rect 122 198 130 200
rect 152 198 160 200
rect 182 198 190 200
rect 212 198 220 200
rect 242 198 250 200
rect 272 198 280 200
rect 302 198 310 200
rect 332 198 340 200
rect 362 198 370 200
rect 392 198 400 200
rect 422 198 430 200
rect 452 198 460 200
rect 482 198 490 200
rect 512 198 520 200
rect 542 198 550 200
rect 42 190 50 198
rect 62 190 80 198
rect 92 190 110 198
rect 122 190 140 198
rect 152 190 170 198
rect 182 190 200 198
rect 212 190 230 198
rect 242 190 260 198
rect 272 190 290 198
rect 302 190 320 198
rect 332 190 350 198
rect 362 190 380 198
rect 392 190 410 198
rect 422 190 440 198
rect 452 190 470 198
rect 482 190 500 198
rect 512 190 530 198
rect 542 190 560 198
rect 62 188 70 190
rect 92 188 100 190
rect 122 188 130 190
rect 152 188 160 190
rect 182 188 190 190
rect 212 188 220 190
rect 242 188 250 190
rect 272 188 280 190
rect 302 188 310 190
rect 332 188 340 190
rect 362 188 370 190
rect 392 188 400 190
rect 422 188 430 190
rect 452 188 460 190
rect 482 188 490 190
rect 512 188 520 190
rect 542 188 550 190
rect 32 180 40 188
rect 52 180 70 188
rect 82 180 100 188
rect 112 180 130 188
rect 142 180 160 188
rect 172 180 190 188
rect 202 180 220 188
rect 232 180 250 188
rect 262 180 280 188
rect 292 180 310 188
rect 322 180 340 188
rect 352 180 370 188
rect 382 180 400 188
rect 412 180 430 188
rect 442 180 460 188
rect 472 180 490 188
rect 502 180 520 188
rect 532 180 550 188
rect 562 180 570 188
rect 62 178 70 180
rect 92 178 100 180
rect 122 178 130 180
rect 152 178 160 180
rect 182 178 190 180
rect 212 178 220 180
rect 242 178 250 180
rect 272 178 280 180
rect 302 178 310 180
rect 332 178 340 180
rect 362 178 370 180
rect 392 178 400 180
rect 422 178 430 180
rect 452 178 460 180
rect 482 178 490 180
rect 512 178 520 180
rect 542 178 550 180
rect 42 170 50 178
rect 62 170 80 178
rect 92 170 110 178
rect 122 170 140 178
rect 152 170 170 178
rect 182 170 200 178
rect 212 170 230 178
rect 242 170 260 178
rect 272 170 290 178
rect 302 170 320 178
rect 332 170 350 178
rect 362 170 380 178
rect 392 170 410 178
rect 422 170 440 178
rect 452 170 470 178
rect 482 170 500 178
rect 512 170 530 178
rect 542 170 560 178
rect 62 168 70 170
rect 92 168 100 170
rect 122 168 130 170
rect 152 168 160 170
rect 182 168 190 170
rect 212 168 220 170
rect 242 168 250 170
rect 272 168 280 170
rect 302 168 310 170
rect 332 168 340 170
rect 362 168 370 170
rect 392 168 400 170
rect 422 168 430 170
rect 452 168 460 170
rect 482 168 490 170
rect 512 168 520 170
rect 542 168 550 170
rect 32 160 40 168
rect 52 160 70 168
rect 82 160 100 168
rect 112 160 130 168
rect 142 160 160 168
rect 172 160 190 168
rect 202 160 220 168
rect 232 160 250 168
rect 262 160 280 168
rect 292 160 310 168
rect 322 160 340 168
rect 352 160 370 168
rect 382 160 400 168
rect 412 160 430 168
rect 442 160 460 168
rect 472 160 490 168
rect 502 160 520 168
rect 532 160 550 168
rect 562 160 570 168
rect 62 158 70 160
rect 42 150 50 158
rect 62 150 80 158
rect 62 148 70 150
rect 92 148 100 160
rect 502 148 510 160
rect 542 158 550 160
rect 522 150 530 158
rect 542 150 560 158
rect 542 148 550 150
rect 32 140 40 148
rect 52 140 70 148
rect 82 140 100 148
rect 112 140 130 148
rect 142 140 160 148
rect 172 140 190 148
rect 202 140 220 148
rect 232 140 250 148
rect 262 140 280 148
rect 292 140 310 148
rect 322 140 340 148
rect 352 140 370 148
rect 382 140 400 148
rect 412 140 430 148
rect 442 140 460 148
rect 472 140 490 148
rect 502 140 520 148
rect 532 140 550 148
rect 562 140 570 148
rect 62 138 70 140
rect 92 138 100 140
rect 122 138 130 140
rect 152 138 160 140
rect 182 138 190 140
rect 212 138 220 140
rect 242 138 250 140
rect 272 138 280 140
rect 302 138 310 140
rect 332 138 340 140
rect 362 138 370 140
rect 392 138 400 140
rect 422 138 430 140
rect 452 138 460 140
rect 482 138 490 140
rect 512 138 520 140
rect 542 138 550 140
rect 42 130 50 138
rect 62 130 80 138
rect 92 130 110 138
rect 122 130 140 138
rect 152 130 170 138
rect 182 130 200 138
rect 212 130 230 138
rect 242 130 260 138
rect 272 130 290 138
rect 302 130 320 138
rect 332 130 350 138
rect 362 130 380 138
rect 392 130 410 138
rect 422 130 440 138
rect 452 130 470 138
rect 482 130 500 138
rect 512 130 530 138
rect 542 130 560 138
rect 62 128 70 130
rect 92 128 100 130
rect 122 128 130 130
rect 152 128 160 130
rect 182 128 190 130
rect 212 128 220 130
rect 242 128 250 130
rect 272 128 280 130
rect 302 128 310 130
rect 332 128 340 130
rect 362 128 370 130
rect 392 128 400 130
rect 422 128 430 130
rect 452 128 460 130
rect 482 128 490 130
rect 512 128 520 130
rect 542 128 550 130
rect 32 120 40 128
rect 52 120 70 128
rect 82 120 100 128
rect 112 120 130 128
rect 142 120 160 128
rect 172 120 190 128
rect 202 120 220 128
rect 232 120 250 128
rect 262 120 280 128
rect 292 120 310 128
rect 322 120 340 128
rect 352 120 370 128
rect 382 120 400 128
rect 412 120 430 128
rect 442 120 460 128
rect 472 120 490 128
rect 502 120 520 128
rect 532 120 550 128
rect 562 120 570 128
rect 62 118 70 120
rect 92 118 100 120
rect 122 118 130 120
rect 152 118 160 120
rect 182 118 190 120
rect 212 118 220 120
rect 242 118 250 120
rect 272 118 280 120
rect 302 118 310 120
rect 332 118 340 120
rect 362 118 370 120
rect 392 118 400 120
rect 422 118 430 120
rect 452 118 460 120
rect 482 118 490 120
rect 512 118 520 120
rect 542 118 550 120
rect 42 110 50 118
rect 62 110 80 118
rect 92 110 110 118
rect 122 110 140 118
rect 152 110 170 118
rect 182 110 200 118
rect 212 110 230 118
rect 242 110 260 118
rect 272 110 290 118
rect 302 110 320 118
rect 332 110 350 118
rect 362 110 380 118
rect 392 110 410 118
rect 422 110 440 118
rect 452 110 470 118
rect 482 110 500 118
rect 512 110 530 118
rect 542 110 560 118
rect 62 108 70 110
rect 92 108 100 110
rect 122 108 130 110
rect 152 108 160 110
rect 182 108 190 110
rect 212 108 220 110
rect 242 108 250 110
rect 272 108 280 110
rect 302 108 310 110
rect 332 108 340 110
rect 362 108 370 110
rect 392 108 400 110
rect 422 108 430 110
rect 452 108 460 110
rect 482 108 490 110
rect 512 108 520 110
rect 542 108 550 110
rect 32 100 40 108
rect 52 100 70 108
rect 82 100 100 108
rect 112 100 130 108
rect 142 100 160 108
rect 172 100 190 108
rect 202 100 220 108
rect 232 100 250 108
rect 262 100 280 108
rect 292 100 310 108
rect 322 100 340 108
rect 352 100 370 108
rect 382 100 400 108
rect 412 100 430 108
rect 442 100 460 108
rect 472 100 490 108
rect 502 100 520 108
rect 532 100 550 108
rect 562 100 570 108
rect 62 98 70 100
rect 92 98 100 100
rect 122 98 130 100
rect 152 98 160 100
rect 182 98 190 100
rect 212 98 220 100
rect 242 98 250 100
rect 272 98 280 100
rect 302 98 310 100
rect 332 98 340 100
rect 362 98 370 100
rect 392 98 400 100
rect 422 98 430 100
rect 452 98 460 100
rect 482 98 490 100
rect 512 98 520 100
rect 542 98 550 100
rect 42 90 50 98
rect 62 90 80 98
rect 92 90 110 98
rect 122 90 140 98
rect 152 90 170 98
rect 182 90 200 98
rect 212 90 230 98
rect 242 90 260 98
rect 272 90 290 98
rect 302 90 320 98
rect 332 90 350 98
rect 362 90 380 98
rect 392 90 410 98
rect 422 90 440 98
rect 452 90 470 98
rect 482 90 500 98
rect 512 90 530 98
rect 542 90 560 98
rect 62 88 70 90
rect 92 88 100 90
rect 122 88 130 90
rect 152 88 160 90
rect 182 88 190 90
rect 212 88 220 90
rect 242 88 250 90
rect 272 88 280 90
rect 302 88 310 90
rect 332 88 340 90
rect 362 88 370 90
rect 392 88 400 90
rect 422 88 430 90
rect 452 88 460 90
rect 482 88 490 90
rect 512 88 520 90
rect 542 88 550 90
rect 32 80 40 88
rect 52 80 70 88
rect 82 80 100 88
rect 112 80 130 88
rect 142 80 160 88
rect 172 80 190 88
rect 202 80 220 88
rect 232 80 250 88
rect 262 80 280 88
rect 292 80 310 88
rect 322 80 340 88
rect 352 80 370 88
rect 382 80 400 88
rect 412 80 430 88
rect 442 80 460 88
rect 472 80 490 88
rect 502 80 520 88
rect 532 80 550 88
rect 562 80 570 88
rect 62 78 70 80
rect 92 78 100 80
rect 122 78 130 80
rect 152 78 160 80
rect 182 78 190 80
rect 212 78 220 80
rect 242 78 250 80
rect 272 78 280 80
rect 302 78 310 80
rect 332 78 340 80
rect 362 78 370 80
rect 392 78 400 80
rect 422 78 430 80
rect 452 78 460 80
rect 482 78 490 80
rect 512 78 520 80
rect 542 78 550 80
rect 42 70 50 78
rect 62 70 80 78
rect 92 70 110 78
rect 122 70 140 78
rect 152 70 170 78
rect 182 70 200 78
rect 212 70 230 78
rect 242 70 260 78
rect 272 70 290 78
rect 302 70 320 78
rect 332 70 350 78
rect 362 70 380 78
rect 392 70 410 78
rect 422 70 440 78
rect 452 70 470 78
rect 482 70 500 78
rect 512 70 530 78
rect 542 70 560 78
rect 62 68 70 70
rect 92 68 100 70
rect 122 68 130 70
rect 152 68 160 70
rect 182 68 190 70
rect 212 68 220 70
rect 242 68 250 70
rect 272 68 280 70
rect 302 68 310 70
rect 332 68 340 70
rect 362 68 370 70
rect 392 68 400 70
rect 422 68 430 70
rect 452 68 460 70
rect 482 68 490 70
rect 512 68 520 70
rect 542 68 550 70
rect 32 60 40 68
rect 52 60 70 68
rect 82 60 100 68
rect 112 60 130 68
rect 142 60 160 68
rect 172 60 190 68
rect 202 60 220 68
rect 232 60 250 68
rect 262 60 280 68
rect 292 60 310 68
rect 322 60 340 68
rect 352 60 370 68
rect 382 60 400 68
rect 412 60 430 68
rect 442 60 460 68
rect 472 60 490 68
rect 502 60 520 68
rect 532 60 550 68
rect 562 60 570 68
rect 62 58 70 60
rect 92 58 100 60
rect 122 58 130 60
rect 152 58 160 60
rect 182 58 190 60
rect 212 58 220 60
rect 242 58 250 60
rect 272 58 280 60
rect 302 58 310 60
rect 332 58 340 60
rect 362 58 370 60
rect 392 58 400 60
rect 422 58 430 60
rect 452 58 460 60
rect 482 58 490 60
rect 512 58 520 60
rect 542 58 550 60
rect 42 50 50 58
rect 62 50 80 58
rect 92 50 110 58
rect 122 50 140 58
rect 152 50 170 58
rect 182 50 200 58
rect 212 50 230 58
rect 242 50 260 58
rect 272 50 290 58
rect 302 50 320 58
rect 332 50 350 58
rect 362 50 380 58
rect 392 50 410 58
rect 422 50 440 58
rect 452 50 470 58
rect 482 50 500 58
rect 512 50 530 58
rect 542 50 560 58
rect 62 48 70 50
rect 92 48 100 50
rect 122 48 130 50
rect 152 48 160 50
rect 182 48 190 50
rect 212 48 220 50
rect 242 48 250 50
rect 272 48 280 50
rect 302 48 310 50
rect 332 48 340 50
rect 362 48 370 50
rect 392 48 400 50
rect 422 48 430 50
rect 452 48 460 50
rect 482 48 490 50
rect 512 48 520 50
rect 542 48 550 50
rect 32 40 40 48
rect 52 40 70 48
rect 82 40 100 48
rect 112 40 130 48
rect 142 40 160 48
rect 172 40 190 48
rect 202 40 220 48
rect 232 40 250 48
rect 262 40 280 48
rect 292 40 310 48
rect 322 40 340 48
rect 352 40 370 48
rect 382 40 400 48
rect 412 40 430 48
rect 442 40 460 48
rect 472 40 490 48
rect 502 40 520 48
rect 532 40 550 48
rect 562 40 570 48
rect 62 38 70 40
rect 92 38 100 40
rect 122 38 130 40
rect 152 38 160 40
rect 182 38 190 40
rect 212 38 220 40
rect 242 38 250 40
rect 272 38 280 40
rect 302 38 310 40
rect 332 38 340 40
rect 362 38 370 40
rect 392 38 400 40
rect 422 38 430 40
rect 452 38 460 40
rect 482 38 490 40
rect 512 38 520 40
rect 542 38 550 40
rect 42 30 50 38
rect 62 30 80 38
rect 92 30 110 38
rect 122 30 140 38
rect 152 30 170 38
rect 182 30 200 38
rect 212 30 230 38
rect 242 30 260 38
rect 272 30 290 38
rect 302 30 320 38
rect 332 30 350 38
rect 362 30 380 38
rect 392 30 410 38
rect 422 30 440 38
rect 452 30 470 38
rect 482 30 500 38
rect 512 30 530 38
rect 542 30 560 38
<< nsubstratencontact >>
rect 46 1290 54 1298
rect 66 1290 84 1298
rect 96 1290 114 1298
rect 126 1290 144 1298
rect 156 1290 174 1298
rect 186 1290 204 1298
rect 216 1290 234 1298
rect 246 1290 264 1298
rect 276 1290 294 1298
rect 306 1290 324 1298
rect 336 1290 354 1298
rect 366 1290 384 1298
rect 396 1290 414 1298
rect 426 1290 444 1298
rect 456 1290 474 1298
rect 486 1290 504 1298
rect 516 1290 534 1298
rect 546 1290 554 1298
rect 76 1288 84 1290
rect 106 1288 114 1290
rect 136 1288 144 1290
rect 166 1288 174 1290
rect 196 1288 204 1290
rect 226 1288 234 1290
rect 256 1288 264 1290
rect 286 1288 294 1290
rect 316 1288 324 1290
rect 346 1288 354 1290
rect 376 1288 384 1290
rect 406 1288 414 1290
rect 436 1288 444 1290
rect 466 1288 474 1290
rect 496 1288 504 1290
rect 526 1288 534 1290
rect 56 1280 64 1288
rect 76 1280 94 1288
rect 106 1280 124 1288
rect 136 1280 154 1288
rect 166 1280 184 1288
rect 196 1280 214 1288
rect 226 1280 244 1288
rect 256 1280 274 1288
rect 286 1280 304 1288
rect 316 1280 334 1288
rect 346 1280 364 1288
rect 376 1280 394 1288
rect 406 1280 424 1288
rect 436 1280 454 1288
rect 466 1280 484 1288
rect 496 1280 514 1288
rect 526 1280 544 1288
rect 76 1278 84 1280
rect 106 1278 114 1280
rect 136 1278 144 1280
rect 166 1278 174 1280
rect 196 1278 204 1280
rect 226 1278 234 1280
rect 256 1278 264 1280
rect 286 1278 294 1280
rect 316 1278 324 1280
rect 346 1278 354 1280
rect 376 1278 384 1280
rect 406 1278 414 1280
rect 436 1278 444 1280
rect 466 1278 474 1280
rect 496 1278 504 1280
rect 526 1278 534 1280
rect 46 1270 54 1278
rect 66 1270 84 1278
rect 96 1270 114 1278
rect 126 1270 144 1278
rect 156 1270 174 1278
rect 186 1270 204 1278
rect 216 1270 234 1278
rect 246 1270 264 1278
rect 276 1270 294 1278
rect 306 1270 324 1278
rect 336 1270 354 1278
rect 366 1270 384 1278
rect 396 1270 414 1278
rect 426 1270 444 1278
rect 456 1270 474 1278
rect 486 1270 504 1278
rect 516 1270 534 1278
rect 546 1270 554 1278
rect 76 1268 84 1270
rect 106 1268 114 1270
rect 136 1268 144 1270
rect 166 1268 174 1270
rect 196 1268 204 1270
rect 226 1268 234 1270
rect 256 1268 264 1270
rect 286 1268 294 1270
rect 316 1268 324 1270
rect 346 1268 354 1270
rect 376 1268 384 1270
rect 406 1268 414 1270
rect 436 1268 444 1270
rect 466 1268 474 1270
rect 496 1268 504 1270
rect 526 1268 534 1270
rect 56 1260 64 1268
rect 76 1260 94 1268
rect 106 1260 124 1268
rect 136 1260 154 1268
rect 166 1260 184 1268
rect 196 1260 214 1268
rect 226 1260 244 1268
rect 256 1260 274 1268
rect 286 1260 304 1268
rect 316 1260 334 1268
rect 346 1260 364 1268
rect 376 1260 394 1268
rect 406 1260 424 1268
rect 436 1260 454 1268
rect 466 1260 484 1268
rect 496 1260 514 1268
rect 526 1260 544 1268
rect 76 1258 84 1260
rect 106 1258 114 1260
rect 136 1258 144 1260
rect 166 1258 174 1260
rect 196 1258 204 1260
rect 226 1258 234 1260
rect 256 1258 264 1260
rect 286 1258 294 1260
rect 316 1258 324 1260
rect 346 1258 354 1260
rect 376 1258 384 1260
rect 406 1258 414 1260
rect 436 1258 444 1260
rect 466 1258 474 1260
rect 496 1258 504 1260
rect 526 1258 534 1260
rect 46 1250 54 1258
rect 66 1250 84 1258
rect 96 1250 114 1258
rect 126 1250 144 1258
rect 156 1250 174 1258
rect 186 1250 204 1258
rect 216 1250 234 1258
rect 246 1250 264 1258
rect 276 1250 294 1258
rect 306 1250 324 1258
rect 336 1250 354 1258
rect 366 1250 384 1258
rect 396 1250 414 1258
rect 426 1250 444 1258
rect 456 1250 474 1258
rect 486 1250 504 1258
rect 516 1250 534 1258
rect 546 1250 554 1258
rect 76 1248 84 1250
rect 106 1248 114 1250
rect 136 1248 144 1250
rect 166 1248 174 1250
rect 196 1248 204 1250
rect 226 1248 234 1250
rect 256 1248 264 1250
rect 286 1248 294 1250
rect 316 1248 324 1250
rect 346 1248 354 1250
rect 376 1248 384 1250
rect 406 1248 414 1250
rect 436 1248 444 1250
rect 466 1248 474 1250
rect 496 1248 504 1250
rect 526 1248 534 1250
rect 56 1240 64 1248
rect 76 1240 94 1248
rect 106 1240 124 1248
rect 136 1240 154 1248
rect 166 1240 184 1248
rect 196 1240 214 1248
rect 226 1240 244 1248
rect 256 1240 274 1248
rect 286 1240 304 1248
rect 316 1240 334 1248
rect 346 1240 364 1248
rect 376 1240 394 1248
rect 406 1240 424 1248
rect 436 1240 454 1248
rect 466 1240 484 1248
rect 496 1240 514 1248
rect 526 1240 544 1248
rect 76 1238 84 1240
rect 106 1238 114 1240
rect 136 1238 144 1240
rect 166 1238 174 1240
rect 196 1238 204 1240
rect 226 1238 234 1240
rect 256 1238 264 1240
rect 286 1238 294 1240
rect 316 1238 324 1240
rect 346 1238 354 1240
rect 376 1238 384 1240
rect 406 1238 414 1240
rect 436 1238 444 1240
rect 466 1238 474 1240
rect 496 1238 504 1240
rect 526 1238 534 1240
rect 46 1230 54 1238
rect 66 1230 84 1238
rect 96 1230 114 1238
rect 126 1230 144 1238
rect 156 1230 174 1238
rect 186 1230 204 1238
rect 216 1230 234 1238
rect 246 1230 264 1238
rect 276 1230 294 1238
rect 306 1230 324 1238
rect 336 1230 354 1238
rect 366 1230 384 1238
rect 396 1230 414 1238
rect 426 1230 444 1238
rect 456 1230 474 1238
rect 486 1230 504 1238
rect 516 1230 534 1238
rect 546 1230 554 1238
rect 76 1228 84 1230
rect 106 1228 114 1230
rect 136 1228 144 1230
rect 166 1228 174 1230
rect 196 1228 204 1230
rect 226 1228 234 1230
rect 256 1228 264 1230
rect 286 1228 294 1230
rect 316 1228 324 1230
rect 346 1228 354 1230
rect 376 1228 384 1230
rect 406 1228 414 1230
rect 436 1228 444 1230
rect 466 1228 474 1230
rect 496 1228 504 1230
rect 526 1228 534 1230
rect 56 1220 64 1228
rect 76 1220 94 1228
rect 106 1220 124 1228
rect 136 1220 154 1228
rect 166 1220 184 1228
rect 196 1220 214 1228
rect 226 1220 244 1228
rect 256 1220 274 1228
rect 286 1220 304 1228
rect 316 1220 334 1228
rect 346 1220 364 1228
rect 376 1220 394 1228
rect 406 1220 424 1228
rect 436 1220 454 1228
rect 466 1220 484 1228
rect 496 1220 514 1228
rect 526 1220 544 1228
rect 76 1218 84 1220
rect 106 1218 114 1220
rect 136 1218 144 1220
rect 166 1218 174 1220
rect 196 1218 204 1220
rect 226 1218 234 1220
rect 256 1218 264 1220
rect 286 1218 294 1220
rect 316 1218 324 1220
rect 346 1218 354 1220
rect 376 1218 384 1220
rect 406 1218 414 1220
rect 436 1218 444 1220
rect 466 1218 474 1220
rect 496 1218 504 1220
rect 526 1218 534 1220
rect 46 1210 54 1218
rect 66 1210 84 1218
rect 96 1210 114 1218
rect 126 1210 144 1218
rect 156 1210 174 1218
rect 186 1210 204 1218
rect 216 1210 234 1218
rect 246 1210 264 1218
rect 276 1210 294 1218
rect 306 1210 324 1218
rect 336 1210 354 1218
rect 366 1210 384 1218
rect 396 1210 414 1218
rect 426 1210 444 1218
rect 456 1210 474 1218
rect 486 1210 504 1218
rect 516 1210 534 1218
rect 546 1210 554 1218
rect 76 1208 84 1210
rect 106 1208 114 1210
rect 136 1208 144 1210
rect 166 1208 174 1210
rect 196 1208 204 1210
rect 226 1208 234 1210
rect 256 1208 264 1210
rect 286 1208 294 1210
rect 316 1208 324 1210
rect 346 1208 354 1210
rect 376 1208 384 1210
rect 406 1208 414 1210
rect 436 1208 444 1210
rect 466 1208 474 1210
rect 496 1208 504 1210
rect 526 1208 534 1210
rect 56 1200 64 1208
rect 76 1200 94 1208
rect 106 1200 124 1208
rect 136 1200 154 1208
rect 166 1200 184 1208
rect 196 1200 214 1208
rect 226 1200 244 1208
rect 256 1200 274 1208
rect 286 1200 304 1208
rect 316 1200 334 1208
rect 346 1200 364 1208
rect 376 1200 394 1208
rect 406 1200 424 1208
rect 436 1200 454 1208
rect 466 1200 484 1208
rect 496 1200 514 1208
rect 526 1200 544 1208
rect 76 1198 84 1200
rect 106 1198 114 1200
rect 136 1198 144 1200
rect 166 1198 174 1200
rect 196 1198 204 1200
rect 226 1198 234 1200
rect 256 1198 264 1200
rect 286 1198 294 1200
rect 316 1198 324 1200
rect 346 1198 354 1200
rect 376 1198 384 1200
rect 406 1198 414 1200
rect 436 1198 444 1200
rect 466 1198 474 1200
rect 496 1198 504 1200
rect 526 1198 534 1200
rect 46 1190 54 1198
rect 66 1190 84 1198
rect 96 1190 114 1198
rect 126 1190 144 1198
rect 156 1190 174 1198
rect 186 1190 204 1198
rect 216 1190 234 1198
rect 246 1190 264 1198
rect 276 1190 294 1198
rect 306 1190 324 1198
rect 336 1190 354 1198
rect 366 1190 384 1198
rect 396 1190 414 1198
rect 426 1190 444 1198
rect 456 1190 474 1198
rect 486 1190 504 1198
rect 516 1190 534 1198
rect 546 1190 554 1198
rect 76 1188 84 1190
rect 526 1188 534 1190
rect 56 1180 64 1188
rect 76 1180 94 1188
rect 506 1180 514 1188
rect 526 1180 544 1188
rect 76 1178 84 1180
rect 526 1178 534 1180
rect 46 1170 54 1178
rect 66 1170 84 1178
rect 96 1170 114 1178
rect 126 1170 144 1178
rect 156 1170 174 1178
rect 186 1170 204 1178
rect 216 1170 234 1178
rect 246 1170 264 1178
rect 276 1170 294 1178
rect 306 1170 324 1178
rect 336 1170 354 1178
rect 366 1170 384 1178
rect 396 1170 414 1178
rect 426 1170 444 1178
rect 456 1170 474 1178
rect 486 1170 504 1178
rect 516 1170 534 1178
rect 546 1170 554 1178
rect 76 1168 84 1170
rect 106 1168 114 1170
rect 136 1168 144 1170
rect 166 1168 174 1170
rect 196 1168 204 1170
rect 226 1168 234 1170
rect 256 1168 264 1170
rect 286 1168 294 1170
rect 316 1168 324 1170
rect 346 1168 354 1170
rect 376 1168 384 1170
rect 406 1168 414 1170
rect 436 1168 444 1170
rect 466 1168 474 1170
rect 496 1168 504 1170
rect 526 1168 534 1170
rect 56 1160 64 1168
rect 76 1160 94 1168
rect 106 1160 124 1168
rect 136 1160 154 1168
rect 166 1160 184 1168
rect 196 1160 214 1168
rect 226 1160 244 1168
rect 256 1160 274 1168
rect 286 1160 304 1168
rect 316 1160 334 1168
rect 346 1160 364 1168
rect 376 1160 394 1168
rect 406 1160 424 1168
rect 436 1160 454 1168
rect 466 1160 484 1168
rect 496 1160 514 1168
rect 526 1160 544 1168
rect 76 1158 84 1160
rect 106 1158 114 1160
rect 136 1158 144 1160
rect 166 1158 174 1160
rect 196 1158 204 1160
rect 226 1158 234 1160
rect 256 1158 264 1160
rect 286 1158 294 1160
rect 316 1158 324 1160
rect 346 1158 354 1160
rect 376 1158 384 1160
rect 406 1158 414 1160
rect 436 1158 444 1160
rect 466 1158 474 1160
rect 496 1158 504 1160
rect 526 1158 534 1160
rect 46 1150 54 1158
rect 66 1150 84 1158
rect 96 1150 114 1158
rect 126 1150 144 1158
rect 156 1150 174 1158
rect 186 1150 204 1158
rect 216 1150 234 1158
rect 246 1150 264 1158
rect 276 1150 294 1158
rect 306 1150 324 1158
rect 336 1150 354 1158
rect 366 1150 384 1158
rect 396 1150 414 1158
rect 426 1150 444 1158
rect 456 1150 474 1158
rect 486 1150 504 1158
rect 516 1150 534 1158
rect 546 1150 554 1158
rect 76 1148 84 1150
rect 106 1148 114 1150
rect 136 1148 144 1150
rect 166 1148 174 1150
rect 196 1148 204 1150
rect 226 1148 234 1150
rect 256 1148 264 1150
rect 286 1148 294 1150
rect 316 1148 324 1150
rect 346 1148 354 1150
rect 376 1148 384 1150
rect 406 1148 414 1150
rect 436 1148 444 1150
rect 466 1148 474 1150
rect 496 1148 504 1150
rect 526 1148 534 1150
rect 56 1140 64 1148
rect 76 1140 94 1148
rect 106 1140 124 1148
rect 136 1140 154 1148
rect 166 1140 184 1148
rect 196 1140 214 1148
rect 226 1140 244 1148
rect 256 1140 274 1148
rect 286 1140 304 1148
rect 316 1140 334 1148
rect 346 1140 364 1148
rect 376 1140 394 1148
rect 406 1140 424 1148
rect 436 1140 454 1148
rect 466 1140 484 1148
rect 496 1140 514 1148
rect 526 1140 544 1148
rect 76 1138 84 1140
rect 106 1138 114 1140
rect 136 1138 144 1140
rect 166 1138 174 1140
rect 196 1138 204 1140
rect 226 1138 234 1140
rect 256 1138 264 1140
rect 286 1138 294 1140
rect 316 1138 324 1140
rect 346 1138 354 1140
rect 376 1138 384 1140
rect 406 1138 414 1140
rect 436 1138 444 1140
rect 466 1138 474 1140
rect 496 1138 504 1140
rect 526 1138 534 1140
rect 46 1130 54 1138
rect 66 1130 84 1138
rect 96 1130 114 1138
rect 126 1130 144 1138
rect 156 1130 174 1138
rect 186 1130 204 1138
rect 216 1130 234 1138
rect 246 1130 264 1138
rect 276 1130 294 1138
rect 306 1130 324 1138
rect 336 1130 354 1138
rect 366 1130 384 1138
rect 396 1130 414 1138
rect 426 1130 444 1138
rect 456 1130 474 1138
rect 486 1130 504 1138
rect 516 1130 534 1138
rect 546 1130 554 1138
rect 76 1128 84 1130
rect 106 1128 114 1130
rect 136 1128 144 1130
rect 166 1128 174 1130
rect 196 1128 204 1130
rect 226 1128 234 1130
rect 256 1128 264 1130
rect 286 1128 294 1130
rect 316 1128 324 1130
rect 346 1128 354 1130
rect 376 1128 384 1130
rect 406 1128 414 1130
rect 436 1128 444 1130
rect 466 1128 474 1130
rect 496 1128 504 1130
rect 526 1128 534 1130
rect 56 1120 64 1128
rect 76 1120 94 1128
rect 106 1120 124 1128
rect 136 1120 154 1128
rect 166 1120 184 1128
rect 196 1120 214 1128
rect 226 1120 244 1128
rect 256 1120 274 1128
rect 286 1120 304 1128
rect 316 1120 334 1128
rect 346 1120 364 1128
rect 376 1120 394 1128
rect 406 1120 424 1128
rect 436 1120 454 1128
rect 466 1120 484 1128
rect 496 1120 514 1128
rect 46 1110 54 1118
rect 66 1110 74 1118
rect 86 1108 94 1120
rect 506 1108 514 1120
rect 56 1100 64 1108
rect 76 1100 94 1108
rect 106 1100 124 1108
rect 136 1100 154 1108
rect 166 1100 184 1108
rect 196 1100 214 1108
rect 226 1100 244 1108
rect 256 1100 274 1108
rect 286 1100 304 1108
rect 316 1100 334 1108
rect 346 1100 364 1108
rect 376 1100 394 1108
rect 406 1100 424 1108
rect 436 1100 454 1108
rect 466 1100 484 1108
rect 496 1100 514 1108
rect 526 1120 544 1128
rect 526 1108 534 1120
rect 546 1110 554 1118
rect 526 1100 544 1108
rect 76 1098 84 1100
rect 106 1098 114 1100
rect 136 1098 144 1100
rect 166 1098 174 1100
rect 196 1098 204 1100
rect 226 1098 234 1100
rect 256 1098 264 1100
rect 286 1098 294 1100
rect 316 1098 324 1100
rect 346 1098 354 1100
rect 376 1098 384 1100
rect 406 1098 414 1100
rect 436 1098 444 1100
rect 466 1098 474 1100
rect 496 1098 504 1100
rect 526 1098 534 1100
rect 46 1090 54 1098
rect 66 1090 84 1098
rect 96 1090 114 1098
rect 126 1090 144 1098
rect 156 1090 174 1098
rect 186 1090 204 1098
rect 216 1090 234 1098
rect 246 1090 264 1098
rect 276 1090 294 1098
rect 306 1090 324 1098
rect 336 1090 354 1098
rect 366 1090 384 1098
rect 396 1090 414 1098
rect 426 1090 444 1098
rect 456 1090 474 1098
rect 486 1090 504 1098
rect 516 1090 534 1098
rect 546 1090 554 1098
rect 76 1088 84 1090
rect 106 1088 114 1090
rect 136 1088 144 1090
rect 166 1088 174 1090
rect 196 1088 204 1090
rect 226 1088 234 1090
rect 256 1088 264 1090
rect 286 1088 294 1090
rect 316 1088 324 1090
rect 346 1088 354 1090
rect 376 1088 384 1090
rect 406 1088 414 1090
rect 436 1088 444 1090
rect 466 1088 474 1090
rect 496 1088 504 1090
rect 526 1088 534 1090
rect 56 1080 64 1088
rect 76 1080 94 1088
rect 106 1080 124 1088
rect 136 1080 154 1088
rect 166 1080 184 1088
rect 196 1080 214 1088
rect 226 1080 244 1088
rect 256 1080 274 1088
rect 286 1080 304 1088
rect 316 1080 334 1088
rect 346 1080 364 1088
rect 376 1080 394 1088
rect 406 1080 424 1088
rect 436 1080 454 1088
rect 466 1080 484 1088
rect 496 1080 514 1088
rect 526 1080 544 1088
rect 76 1078 84 1080
rect 106 1078 114 1080
rect 136 1078 144 1080
rect 166 1078 174 1080
rect 196 1078 204 1080
rect 226 1078 234 1080
rect 256 1078 264 1080
rect 286 1078 294 1080
rect 316 1078 324 1080
rect 346 1078 354 1080
rect 376 1078 384 1080
rect 406 1078 414 1080
rect 436 1078 444 1080
rect 466 1078 474 1080
rect 496 1078 504 1080
rect 526 1078 534 1080
rect 46 1070 54 1078
rect 66 1070 84 1078
rect 96 1070 114 1078
rect 126 1070 144 1078
rect 156 1070 174 1078
rect 186 1070 204 1078
rect 216 1070 234 1078
rect 246 1070 264 1078
rect 276 1070 294 1078
rect 306 1070 324 1078
rect 336 1070 354 1078
rect 366 1070 384 1078
rect 396 1070 414 1078
rect 426 1070 444 1078
rect 456 1070 474 1078
rect 486 1070 504 1078
rect 516 1070 534 1078
rect 546 1070 554 1078
rect 76 1068 84 1070
rect 106 1068 114 1070
rect 136 1068 144 1070
rect 166 1068 174 1070
rect 196 1068 204 1070
rect 226 1068 234 1070
rect 256 1068 264 1070
rect 286 1068 294 1070
rect 316 1068 324 1070
rect 346 1068 354 1070
rect 376 1068 384 1070
rect 406 1068 414 1070
rect 436 1068 444 1070
rect 466 1068 474 1070
rect 496 1068 504 1070
rect 526 1068 534 1070
rect 56 1060 64 1068
rect 76 1060 94 1068
rect 106 1060 124 1068
rect 136 1060 154 1068
rect 166 1060 184 1068
rect 196 1060 214 1068
rect 226 1060 244 1068
rect 256 1060 274 1068
rect 286 1060 304 1068
rect 316 1060 334 1068
rect 346 1060 364 1068
rect 376 1060 394 1068
rect 406 1060 424 1068
rect 436 1060 454 1068
rect 466 1060 484 1068
rect 496 1060 514 1068
rect 526 1060 544 1068
rect 76 1058 84 1060
rect 106 1058 114 1060
rect 136 1058 144 1060
rect 166 1058 174 1060
rect 196 1058 204 1060
rect 226 1058 234 1060
rect 256 1058 264 1060
rect 286 1058 294 1060
rect 316 1058 324 1060
rect 346 1058 354 1060
rect 376 1058 384 1060
rect 406 1058 414 1060
rect 436 1058 444 1060
rect 466 1058 474 1060
rect 496 1058 504 1060
rect 526 1058 534 1060
rect 46 1050 54 1058
rect 66 1050 84 1058
rect 96 1050 114 1058
rect 126 1050 144 1058
rect 156 1050 174 1058
rect 186 1050 204 1058
rect 216 1050 234 1058
rect 246 1050 264 1058
rect 276 1050 294 1058
rect 306 1050 324 1058
rect 336 1050 354 1058
rect 366 1050 384 1058
rect 396 1050 414 1058
rect 426 1050 444 1058
rect 456 1050 474 1058
rect 486 1050 504 1058
rect 516 1050 534 1058
rect 546 1050 554 1058
rect 76 1048 84 1050
rect 106 1048 114 1050
rect 136 1048 144 1050
rect 166 1048 174 1050
rect 196 1048 204 1050
rect 226 1048 234 1050
rect 256 1048 264 1050
rect 286 1048 294 1050
rect 316 1048 324 1050
rect 346 1048 354 1050
rect 376 1048 384 1050
rect 406 1048 414 1050
rect 436 1048 444 1050
rect 466 1048 474 1050
rect 496 1048 504 1050
rect 526 1048 534 1050
rect 56 1040 64 1048
rect 76 1040 94 1048
rect 106 1040 124 1048
rect 136 1040 154 1048
rect 166 1040 184 1048
rect 196 1040 214 1048
rect 226 1040 244 1048
rect 256 1040 274 1048
rect 286 1040 304 1048
rect 316 1040 334 1048
rect 346 1040 364 1048
rect 376 1040 394 1048
rect 406 1040 424 1048
rect 436 1040 454 1048
rect 466 1040 484 1048
rect 496 1040 514 1048
rect 76 1038 84 1040
rect 46 1030 54 1038
rect 66 1030 84 1038
rect 76 1028 84 1030
rect 506 1028 514 1040
rect 56 1020 64 1028
rect 76 1020 94 1028
rect 106 1020 124 1028
rect 136 1020 154 1028
rect 166 1020 184 1028
rect 196 1020 214 1028
rect 226 1020 244 1028
rect 256 1020 274 1028
rect 286 1020 304 1028
rect 316 1020 334 1028
rect 346 1020 364 1028
rect 376 1020 394 1028
rect 406 1020 424 1028
rect 436 1020 454 1028
rect 466 1020 484 1028
rect 496 1020 514 1028
rect 526 1040 544 1048
rect 526 1028 534 1040
rect 546 1030 554 1038
rect 526 1020 544 1028
rect 76 1018 84 1020
rect 106 1018 114 1020
rect 136 1018 144 1020
rect 166 1018 174 1020
rect 196 1018 204 1020
rect 226 1018 234 1020
rect 256 1018 264 1020
rect 286 1018 294 1020
rect 316 1018 324 1020
rect 346 1018 354 1020
rect 376 1018 384 1020
rect 406 1018 414 1020
rect 436 1018 444 1020
rect 466 1018 474 1020
rect 496 1018 504 1020
rect 526 1018 534 1020
rect 46 1010 54 1018
rect 66 1010 84 1018
rect 96 1010 114 1018
rect 126 1010 144 1018
rect 156 1010 174 1018
rect 186 1010 204 1018
rect 216 1010 234 1018
rect 246 1010 264 1018
rect 276 1010 294 1018
rect 306 1010 324 1018
rect 336 1010 354 1018
rect 366 1010 384 1018
rect 396 1010 414 1018
rect 426 1010 444 1018
rect 456 1010 474 1018
rect 486 1010 504 1018
rect 516 1010 534 1018
rect 546 1010 554 1018
rect 76 1008 84 1010
rect 106 1008 114 1010
rect 136 1008 144 1010
rect 166 1008 174 1010
rect 196 1008 204 1010
rect 226 1008 234 1010
rect 256 1008 264 1010
rect 286 1008 294 1010
rect 316 1008 324 1010
rect 346 1008 354 1010
rect 376 1008 384 1010
rect 406 1008 414 1010
rect 436 1008 444 1010
rect 466 1008 474 1010
rect 496 1008 504 1010
rect 526 1008 534 1010
rect 56 1000 64 1008
rect 76 1000 94 1008
rect 106 1000 124 1008
rect 136 1000 154 1008
rect 166 1000 184 1008
rect 196 1000 214 1008
rect 226 1000 244 1008
rect 256 1000 274 1008
rect 286 1000 304 1008
rect 316 1000 334 1008
rect 346 1000 364 1008
rect 376 1000 394 1008
rect 406 1000 424 1008
rect 436 1000 454 1008
rect 466 1000 484 1008
rect 496 1000 514 1008
rect 526 1000 544 1008
rect 76 998 84 1000
rect 106 998 114 1000
rect 136 998 144 1000
rect 166 998 174 1000
rect 196 998 204 1000
rect 226 998 234 1000
rect 256 998 264 1000
rect 286 998 294 1000
rect 316 998 324 1000
rect 346 998 354 1000
rect 376 998 384 1000
rect 406 998 414 1000
rect 436 998 444 1000
rect 466 998 474 1000
rect 496 998 504 1000
rect 526 998 534 1000
rect 46 990 54 998
rect 66 990 84 998
rect 96 990 114 998
rect 126 990 144 998
rect 156 990 174 998
rect 186 990 204 998
rect 216 990 234 998
rect 246 990 264 998
rect 276 990 294 998
rect 306 990 324 998
rect 336 990 354 998
rect 366 990 384 998
rect 396 990 414 998
rect 426 990 444 998
rect 456 990 474 998
rect 486 990 504 998
rect 516 990 534 998
rect 546 990 554 998
rect 76 988 84 990
rect 106 988 114 990
rect 136 988 144 990
rect 166 988 174 990
rect 196 988 204 990
rect 226 988 234 990
rect 256 988 264 990
rect 286 988 294 990
rect 316 988 324 990
rect 346 988 354 990
rect 376 988 384 990
rect 406 988 414 990
rect 436 988 444 990
rect 466 988 474 990
rect 496 988 504 990
rect 526 988 534 990
rect 56 980 64 988
rect 76 980 94 988
rect 106 980 124 988
rect 136 980 154 988
rect 166 980 184 988
rect 196 980 214 988
rect 226 980 244 988
rect 256 980 274 988
rect 286 980 304 988
rect 316 980 334 988
rect 346 980 364 988
rect 376 980 394 988
rect 406 980 424 988
rect 436 980 454 988
rect 466 980 484 988
rect 496 980 514 988
rect 526 980 544 988
rect 76 978 84 980
rect 106 978 114 980
rect 136 978 144 980
rect 166 978 174 980
rect 196 978 204 980
rect 226 978 234 980
rect 256 978 264 980
rect 286 978 294 980
rect 316 978 324 980
rect 346 978 354 980
rect 376 978 384 980
rect 406 978 414 980
rect 436 978 444 980
rect 466 978 474 980
rect 496 978 504 980
rect 526 978 534 980
rect 46 970 54 978
rect 66 970 84 978
rect 96 970 114 978
rect 126 970 144 978
rect 156 970 174 978
rect 186 970 204 978
rect 216 970 234 978
rect 246 970 264 978
rect 276 970 294 978
rect 306 970 324 978
rect 336 970 354 978
rect 366 970 384 978
rect 396 970 414 978
rect 426 970 444 978
rect 456 970 474 978
rect 486 970 504 978
rect 516 970 534 978
rect 546 970 554 978
rect 536 960 544 968
rect 46 950 54 958
rect 66 950 84 958
rect 96 950 114 958
rect 126 950 144 958
rect 156 950 174 958
rect 186 950 204 958
rect 216 950 234 958
rect 246 950 264 958
rect 276 950 294 958
rect 306 950 324 958
rect 336 950 354 958
rect 366 950 384 958
rect 396 950 414 958
rect 426 950 444 958
rect 456 950 474 958
rect 486 950 504 958
rect 516 950 534 958
rect 546 950 554 958
rect 76 948 84 950
rect 106 948 114 950
rect 136 948 144 950
rect 166 948 174 950
rect 196 948 204 950
rect 226 948 234 950
rect 256 948 264 950
rect 286 948 294 950
rect 316 948 324 950
rect 346 948 354 950
rect 376 948 384 950
rect 406 948 414 950
rect 436 948 444 950
rect 466 948 474 950
rect 496 948 504 950
rect 526 948 534 950
rect 56 940 64 948
rect 76 940 94 948
rect 106 940 124 948
rect 136 940 154 948
rect 166 940 184 948
rect 196 940 214 948
rect 226 940 244 948
rect 256 940 274 948
rect 286 940 304 948
rect 316 940 334 948
rect 346 940 364 948
rect 376 940 394 948
rect 406 940 424 948
rect 436 940 454 948
rect 466 940 484 948
rect 496 940 514 948
rect 526 940 544 948
rect 76 938 84 940
rect 106 938 114 940
rect 136 938 144 940
rect 166 938 174 940
rect 196 938 204 940
rect 226 938 234 940
rect 256 938 264 940
rect 286 938 294 940
rect 316 938 324 940
rect 346 938 354 940
rect 376 938 384 940
rect 406 938 414 940
rect 436 938 444 940
rect 466 938 474 940
rect 496 938 504 940
rect 526 938 534 940
rect 46 930 54 938
rect 66 930 84 938
rect 96 930 114 938
rect 126 930 144 938
rect 156 930 174 938
rect 186 930 204 938
rect 216 930 234 938
rect 246 930 264 938
rect 276 930 294 938
rect 306 930 324 938
rect 336 930 354 938
rect 366 930 384 938
rect 396 930 414 938
rect 426 930 444 938
rect 456 930 474 938
rect 486 930 504 938
rect 516 930 534 938
rect 546 930 554 938
rect 76 928 84 930
rect 106 928 114 930
rect 136 928 144 930
rect 166 928 174 930
rect 196 928 204 930
rect 226 928 234 930
rect 256 928 264 930
rect 286 928 294 930
rect 316 928 324 930
rect 346 928 354 930
rect 376 928 384 930
rect 406 928 414 930
rect 436 928 444 930
rect 466 928 474 930
rect 496 928 504 930
rect 526 928 534 930
rect 56 920 64 928
rect 76 920 94 928
rect 106 920 124 928
rect 136 920 154 928
rect 166 920 184 928
rect 196 920 214 928
rect 226 920 244 928
rect 256 920 274 928
rect 286 920 304 928
rect 316 920 334 928
rect 346 920 364 928
rect 376 920 394 928
rect 406 920 424 928
rect 436 920 454 928
rect 466 920 484 928
rect 496 920 514 928
rect 526 920 544 928
rect 76 918 84 920
rect 106 918 114 920
rect 136 918 144 920
rect 166 918 174 920
rect 196 918 204 920
rect 226 918 234 920
rect 256 918 264 920
rect 286 918 294 920
rect 316 918 324 920
rect 346 918 354 920
rect 376 918 384 920
rect 406 918 414 920
rect 436 918 444 920
rect 466 918 474 920
rect 496 918 504 920
rect 526 918 534 920
rect 46 910 54 918
rect 66 910 84 918
rect 96 910 114 918
rect 126 910 144 918
rect 156 910 174 918
rect 186 910 204 918
rect 216 910 234 918
rect 246 910 264 918
rect 276 910 294 918
rect 306 910 324 918
rect 336 910 354 918
rect 366 910 384 918
rect 396 910 414 918
rect 426 910 444 918
rect 456 910 474 918
rect 486 910 504 918
rect 516 910 534 918
rect 546 910 554 918
rect 76 908 84 910
rect 106 908 114 910
rect 136 908 144 910
rect 166 908 174 910
rect 196 908 204 910
rect 226 908 234 910
rect 256 908 264 910
rect 286 908 294 910
rect 316 908 324 910
rect 346 908 354 910
rect 376 908 384 910
rect 406 908 414 910
rect 436 908 444 910
rect 466 908 474 910
rect 496 908 504 910
rect 526 908 534 910
rect 56 900 64 908
rect 76 900 94 908
rect 106 900 124 908
rect 136 900 154 908
rect 166 900 184 908
rect 196 900 214 908
rect 226 900 244 908
rect 256 900 274 908
rect 286 900 304 908
rect 316 900 334 908
rect 346 900 364 908
rect 376 900 394 908
rect 406 900 424 908
rect 436 900 454 908
rect 466 900 484 908
rect 496 900 514 908
rect 526 900 544 908
rect 76 898 84 900
rect 106 898 114 900
rect 136 898 144 900
rect 166 898 174 900
rect 196 898 204 900
rect 226 898 234 900
rect 256 898 264 900
rect 286 898 294 900
rect 316 898 324 900
rect 346 898 354 900
rect 376 898 384 900
rect 406 898 414 900
rect 436 898 444 900
rect 466 898 474 900
rect 496 898 504 900
rect 526 898 534 900
rect 46 890 54 898
rect 66 890 84 898
rect 96 890 114 898
rect 126 890 144 898
rect 156 890 174 898
rect 186 890 204 898
rect 216 890 234 898
rect 246 890 264 898
rect 276 890 294 898
rect 306 890 324 898
rect 336 890 354 898
rect 366 890 384 898
rect 396 890 414 898
rect 426 890 444 898
rect 456 890 474 898
rect 486 890 504 898
rect 516 890 534 898
rect 546 890 554 898
rect 76 888 84 890
rect 106 888 114 890
rect 136 888 144 890
rect 166 888 174 890
rect 196 888 204 890
rect 226 888 234 890
rect 256 888 264 890
rect 286 888 294 890
rect 316 888 324 890
rect 346 888 354 890
rect 376 888 384 890
rect 406 888 414 890
rect 436 888 444 890
rect 466 888 474 890
rect 496 888 504 890
rect 526 888 534 890
rect 56 878 64 888
rect 76 878 94 888
rect 106 878 124 888
rect 136 878 154 888
rect 166 878 184 888
rect 196 878 214 888
rect 226 878 244 888
rect 256 878 274 888
rect 286 878 304 888
rect 316 878 334 888
rect 346 878 364 888
rect 376 878 394 888
rect 406 878 424 888
rect 436 878 454 888
rect 466 878 484 888
rect 496 878 514 888
rect 526 878 544 888
rect 46 870 554 878
rect 4 644 12 652
rect 24 644 42 652
rect 54 644 72 652
rect 84 644 102 652
rect 114 644 132 652
rect 144 644 162 652
rect 174 644 192 652
rect 204 644 222 652
rect 234 644 242 652
rect 256 644 264 652
rect 276 644 294 652
rect 306 644 324 652
rect 336 644 344 652
rect 358 644 366 652
rect 378 644 396 652
rect 408 644 426 652
rect 438 644 456 652
rect 468 644 486 652
rect 498 644 516 652
rect 528 644 546 652
rect 558 644 576 652
rect 588 644 596 652
rect 34 642 42 644
rect 64 642 72 644
rect 94 642 102 644
rect 124 642 132 644
rect 154 642 162 644
rect 184 642 192 644
rect 214 642 222 644
rect 286 642 294 644
rect 316 642 324 644
rect 378 642 386 644
rect 408 642 416 644
rect 438 642 446 644
rect 468 642 476 644
rect 498 642 506 644
rect 528 642 536 644
rect 558 642 566 644
rect 14 634 22 642
rect 34 634 52 642
rect 64 634 82 642
rect 94 634 112 642
rect 124 634 142 642
rect 154 634 172 642
rect 184 634 202 642
rect 214 634 232 642
rect 244 634 252 642
rect 266 634 274 642
rect 286 634 304 642
rect 316 634 334 642
rect 348 634 356 642
rect 368 634 386 642
rect 398 634 416 642
rect 428 634 446 642
rect 458 634 476 642
rect 488 634 506 642
rect 518 634 536 642
rect 548 634 566 642
rect 578 634 586 642
rect 34 632 42 634
rect 64 632 72 634
rect 94 632 102 634
rect 124 632 132 634
rect 154 632 162 634
rect 184 632 192 634
rect 214 632 222 634
rect 286 632 294 634
rect 316 632 324 634
rect 378 632 386 634
rect 408 632 416 634
rect 438 632 446 634
rect 468 632 476 634
rect 498 632 506 634
rect 528 632 536 634
rect 558 632 566 634
rect 4 624 12 632
rect 24 624 42 632
rect 54 624 72 632
rect 84 624 102 632
rect 114 624 132 632
rect 144 624 162 632
rect 174 624 192 632
rect 204 624 222 632
rect 234 624 242 632
rect 256 624 264 632
rect 276 624 294 632
rect 306 624 324 632
rect 336 624 344 632
rect 358 624 366 632
rect 378 624 396 632
rect 408 624 426 632
rect 438 624 456 632
rect 468 624 486 632
rect 498 624 516 632
rect 528 624 546 632
rect 558 624 576 632
rect 588 624 596 632
rect 34 622 42 624
rect 64 622 72 624
rect 94 622 102 624
rect 124 622 132 624
rect 154 622 162 624
rect 184 622 192 624
rect 214 622 222 624
rect 286 622 294 624
rect 316 622 324 624
rect 378 622 386 624
rect 408 622 416 624
rect 438 622 446 624
rect 468 622 476 624
rect 498 622 506 624
rect 528 622 536 624
rect 558 622 566 624
rect 14 614 22 622
rect 34 614 52 622
rect 64 614 82 622
rect 94 614 112 622
rect 124 614 142 622
rect 154 614 172 622
rect 184 614 202 622
rect 214 614 232 622
rect 244 614 252 622
rect 266 614 274 622
rect 286 614 304 622
rect 316 614 334 622
rect 348 614 356 622
rect 368 614 386 622
rect 398 614 416 622
rect 428 614 446 622
rect 458 614 476 622
rect 488 614 506 622
rect 518 614 536 622
rect 548 614 566 622
rect 578 614 586 622
rect 4 604 12 612
rect 24 604 32 612
rect 214 602 222 614
rect 286 612 294 614
rect 316 612 324 614
rect 234 604 242 612
rect 256 604 264 612
rect 276 604 294 612
rect 306 604 324 612
rect 336 604 344 612
rect 358 604 366 612
rect 286 602 294 604
rect 316 602 324 604
rect 378 602 386 614
rect 568 604 576 612
rect 588 604 596 612
rect 14 594 22 602
rect 34 594 52 602
rect 64 594 82 602
rect 94 594 112 602
rect 124 594 142 602
rect 154 594 172 602
rect 184 594 202 602
rect 214 594 232 602
rect 244 594 252 602
rect 34 592 42 594
rect 64 592 72 594
rect 94 592 102 594
rect 124 592 132 594
rect 154 592 162 594
rect 184 592 192 594
rect 214 592 222 594
rect 266 592 274 602
rect 286 592 304 602
rect 316 592 334 602
rect 348 594 356 602
rect 368 594 386 602
rect 398 594 416 602
rect 428 594 446 602
rect 458 594 476 602
rect 488 594 506 602
rect 518 594 536 602
rect 548 594 566 602
rect 578 594 586 602
rect 378 592 386 594
rect 408 592 416 594
rect 438 592 446 594
rect 468 592 476 594
rect 498 592 506 594
rect 528 592 536 594
rect 558 592 566 594
rect 4 584 12 592
rect 24 584 42 592
rect 54 584 72 592
rect 84 584 102 592
rect 34 582 42 584
rect 64 582 72 584
rect 94 582 102 584
rect 114 582 132 592
rect 144 582 162 592
rect 174 582 192 592
rect 204 582 222 592
rect 234 582 242 592
rect 14 574 22 582
rect 34 574 52 582
rect 64 574 82 582
rect 94 574 252 582
rect 256 574 344 592
rect 358 582 366 592
rect 378 582 396 592
rect 408 582 426 592
rect 438 582 456 592
rect 468 582 486 592
rect 498 584 516 592
rect 528 584 546 592
rect 558 584 576 592
rect 588 584 596 592
rect 498 582 506 584
rect 528 582 536 584
rect 558 582 566 584
rect 348 574 506 582
rect 518 574 536 582
rect 548 574 566 582
rect 578 574 586 582
rect 34 572 42 574
rect 64 572 72 574
rect 94 572 102 574
rect 4 564 12 572
rect 24 564 42 572
rect 54 564 72 572
rect 84 564 102 572
rect 114 564 132 574
rect 144 564 162 574
rect 174 564 192 574
rect 204 564 222 574
rect 234 564 242 574
rect 256 564 264 574
rect 276 564 294 574
rect 306 564 324 574
rect 336 564 344 574
rect 358 564 366 574
rect 378 564 396 574
rect 408 564 426 574
rect 438 564 456 574
rect 468 564 486 574
rect 498 572 506 574
rect 528 572 536 574
rect 558 572 566 574
rect 498 564 516 572
rect 528 564 546 572
rect 558 564 576 572
rect 588 564 596 572
rect 34 562 42 564
rect 64 562 72 564
rect 94 562 102 564
rect 124 562 132 564
rect 154 562 162 564
rect 184 562 192 564
rect 214 562 222 564
rect 286 562 294 564
rect 316 562 324 564
rect 378 562 386 564
rect 408 562 416 564
rect 438 562 446 564
rect 468 562 476 564
rect 498 562 506 564
rect 528 562 536 564
rect 558 562 566 564
rect 14 554 22 562
rect 34 554 52 562
rect 64 554 82 562
rect 94 554 112 562
rect 124 554 142 562
rect 154 554 172 562
rect 184 554 202 562
rect 214 554 232 562
rect 244 554 252 562
rect 266 554 274 562
rect 286 554 304 562
rect 316 554 334 562
rect 348 554 356 562
rect 368 554 386 562
rect 398 554 416 562
rect 428 554 446 562
rect 458 554 476 562
rect 488 554 506 562
rect 518 554 536 562
rect 548 554 566 562
rect 578 554 586 562
rect 34 552 42 554
rect 64 552 72 554
rect 94 552 102 554
rect 124 552 132 554
rect 154 552 162 554
rect 184 552 192 554
rect 214 552 222 554
rect 286 552 294 554
rect 316 552 324 554
rect 378 552 386 554
rect 408 552 416 554
rect 438 552 446 554
rect 468 552 476 554
rect 498 552 506 554
rect 528 552 536 554
rect 558 552 566 554
rect 4 544 12 552
rect 24 544 42 552
rect 54 544 72 552
rect 84 544 102 552
rect 114 544 132 552
rect 144 544 162 552
rect 174 544 192 552
rect 204 544 222 552
rect 234 544 242 552
rect 256 544 264 552
rect 276 544 294 552
rect 306 544 324 552
rect 336 544 344 552
rect 358 544 366 552
rect 378 544 396 552
rect 408 544 426 552
rect 438 544 456 552
rect 468 544 486 552
rect 498 544 516 552
rect 528 544 546 552
rect 558 544 576 552
rect 588 544 596 552
rect 34 542 42 544
rect 64 542 72 544
rect 94 542 102 544
rect 124 542 132 544
rect 154 542 162 544
rect 184 542 192 544
rect 214 542 222 544
rect 286 542 294 544
rect 316 542 324 544
rect 378 542 386 544
rect 408 542 416 544
rect 438 542 446 544
rect 468 542 476 544
rect 498 542 506 544
rect 528 542 536 544
rect 558 542 566 544
rect 14 534 22 542
rect 34 534 52 542
rect 64 534 82 542
rect 94 534 112 542
rect 124 534 142 542
rect 154 534 172 542
rect 184 534 202 542
rect 214 534 232 542
rect 244 534 252 542
rect 266 534 274 542
rect 286 534 304 542
rect 316 534 334 542
rect 348 534 356 542
rect 368 534 386 542
rect 398 534 416 542
rect 428 534 446 542
rect 458 534 476 542
rect 488 534 506 542
rect 518 534 536 542
rect 548 534 566 542
rect 578 534 586 542
rect 34 532 42 534
rect 64 532 72 534
rect 94 532 102 534
rect 124 532 132 534
rect 154 532 162 534
rect 184 532 192 534
rect 214 532 222 534
rect 286 532 294 534
rect 316 532 324 534
rect 378 532 386 534
rect 408 532 416 534
rect 438 532 446 534
rect 468 532 476 534
rect 498 532 506 534
rect 528 532 536 534
rect 558 532 566 534
rect 4 524 12 532
rect 24 524 42 532
rect 54 524 72 532
rect 84 524 102 532
rect 114 524 132 532
rect 144 524 162 532
rect 174 524 192 532
rect 204 524 222 532
rect 234 524 242 532
rect 256 524 264 532
rect 276 524 294 532
rect 306 524 324 532
rect 336 524 344 532
rect 358 524 366 532
rect 378 524 396 532
rect 408 524 426 532
rect 438 524 456 532
rect 468 524 486 532
rect 498 524 516 532
rect 528 524 546 532
rect 558 524 576 532
rect 588 524 596 532
rect 4 4 12 512
rect 24 508 32 516
rect 44 508 52 516
rect 64 508 72 516
rect 84 508 92 516
rect 104 508 112 516
rect 124 508 132 516
rect 144 508 152 516
rect 164 508 172 516
rect 184 508 192 516
rect 204 508 212 516
rect 224 508 232 516
rect 244 508 252 516
rect 264 508 272 516
rect 284 508 292 516
rect 318 508 326 516
rect 338 508 346 516
rect 358 508 366 516
rect 378 508 386 516
rect 398 508 406 516
rect 418 508 426 516
rect 438 508 446 516
rect 458 508 466 516
rect 478 508 486 516
rect 498 508 506 516
rect 518 508 526 516
rect 538 508 546 516
rect 558 508 566 516
rect 578 512 586 516
rect 578 508 596 512
rect 16 4 584 12
rect 588 4 596 508
<< metal1 >>
rect 0 1336 600 1340
rect 0 828 4 1336
rect 332 1328 338 1336
rect 12 1326 588 1328
rect 12 838 14 1326
rect 100 1298 560 1300
rect 42 1290 46 1298
rect 54 1290 56 1298
rect 64 1290 66 1298
rect 84 1290 86 1298
rect 94 1290 96 1298
rect 114 1290 116 1298
rect 124 1290 126 1298
rect 144 1290 146 1298
rect 154 1290 156 1298
rect 174 1290 176 1298
rect 184 1290 186 1298
rect 204 1290 206 1298
rect 214 1290 216 1298
rect 234 1290 236 1298
rect 244 1290 246 1298
rect 264 1290 266 1298
rect 274 1290 276 1298
rect 294 1290 296 1298
rect 304 1290 306 1298
rect 324 1290 326 1298
rect 334 1290 336 1298
rect 354 1290 356 1298
rect 364 1290 366 1298
rect 384 1290 386 1298
rect 394 1290 396 1298
rect 414 1290 416 1298
rect 424 1290 426 1298
rect 444 1290 446 1298
rect 454 1290 456 1298
rect 474 1290 476 1298
rect 484 1290 486 1298
rect 504 1290 506 1298
rect 514 1290 516 1298
rect 534 1290 536 1298
rect 544 1290 546 1298
rect 554 1290 560 1298
rect 42 1288 76 1290
rect 84 1288 106 1290
rect 114 1288 136 1290
rect 144 1288 166 1290
rect 174 1288 196 1290
rect 204 1288 226 1290
rect 234 1288 256 1290
rect 264 1288 286 1290
rect 294 1288 316 1290
rect 324 1288 346 1290
rect 354 1288 376 1290
rect 384 1288 406 1290
rect 414 1288 436 1290
rect 444 1288 466 1290
rect 474 1288 496 1290
rect 504 1288 526 1290
rect 534 1288 560 1290
rect 42 1280 46 1288
rect 54 1280 56 1288
rect 64 1280 66 1288
rect 74 1280 76 1288
rect 94 1280 96 1288
rect 104 1280 106 1288
rect 124 1280 126 1288
rect 134 1280 136 1288
rect 154 1280 156 1288
rect 164 1280 166 1288
rect 184 1280 186 1288
rect 194 1280 196 1288
rect 214 1280 216 1288
rect 224 1280 226 1288
rect 244 1280 246 1288
rect 254 1280 256 1288
rect 274 1280 276 1288
rect 284 1280 286 1288
rect 304 1280 306 1288
rect 314 1280 316 1288
rect 334 1280 336 1288
rect 344 1280 346 1288
rect 364 1280 366 1288
rect 374 1280 376 1288
rect 394 1280 396 1288
rect 404 1280 406 1288
rect 424 1280 426 1288
rect 434 1280 436 1288
rect 454 1280 456 1288
rect 464 1280 466 1288
rect 484 1280 486 1288
rect 494 1280 496 1288
rect 514 1280 516 1288
rect 524 1280 526 1288
rect 544 1280 546 1288
rect 554 1280 560 1288
rect 42 1278 76 1280
rect 84 1278 106 1280
rect 114 1278 136 1280
rect 144 1278 166 1280
rect 174 1278 196 1280
rect 204 1278 226 1280
rect 234 1278 256 1280
rect 264 1278 286 1280
rect 294 1278 316 1280
rect 324 1278 346 1280
rect 354 1278 376 1280
rect 384 1278 406 1280
rect 414 1278 436 1280
rect 444 1278 466 1280
rect 474 1278 496 1280
rect 504 1278 526 1280
rect 534 1278 560 1280
rect 42 1270 46 1278
rect 54 1270 56 1278
rect 64 1270 66 1278
rect 84 1270 86 1278
rect 94 1270 96 1278
rect 114 1270 116 1278
rect 124 1270 126 1278
rect 144 1270 146 1278
rect 154 1270 156 1278
rect 174 1270 176 1278
rect 184 1270 186 1278
rect 204 1270 206 1278
rect 214 1270 216 1278
rect 234 1270 236 1278
rect 244 1270 246 1278
rect 264 1270 266 1278
rect 274 1270 276 1278
rect 294 1270 296 1278
rect 304 1270 306 1278
rect 324 1270 326 1278
rect 334 1270 336 1278
rect 354 1270 356 1278
rect 364 1270 366 1278
rect 384 1270 386 1278
rect 394 1270 396 1278
rect 414 1270 416 1278
rect 424 1270 426 1278
rect 444 1270 446 1278
rect 454 1270 456 1278
rect 474 1270 476 1278
rect 484 1270 486 1278
rect 504 1270 506 1278
rect 514 1270 516 1278
rect 534 1270 536 1278
rect 544 1270 546 1278
rect 554 1270 560 1278
rect 42 1268 76 1270
rect 84 1268 106 1270
rect 114 1268 136 1270
rect 144 1268 166 1270
rect 174 1268 196 1270
rect 204 1268 226 1270
rect 234 1268 256 1270
rect 264 1268 286 1270
rect 294 1268 316 1270
rect 324 1268 346 1270
rect 354 1268 376 1270
rect 384 1268 406 1270
rect 414 1268 436 1270
rect 444 1268 466 1270
rect 474 1268 496 1270
rect 504 1268 526 1270
rect 534 1268 560 1270
rect 42 1260 46 1268
rect 54 1260 56 1268
rect 64 1260 66 1268
rect 74 1260 76 1268
rect 94 1260 96 1268
rect 104 1260 106 1268
rect 124 1260 126 1268
rect 134 1260 136 1268
rect 154 1260 156 1268
rect 164 1260 166 1268
rect 184 1260 186 1268
rect 194 1260 196 1268
rect 214 1260 216 1268
rect 224 1260 226 1268
rect 244 1260 246 1268
rect 254 1260 256 1268
rect 274 1260 276 1268
rect 284 1260 286 1268
rect 304 1260 306 1268
rect 314 1260 316 1268
rect 334 1260 336 1268
rect 344 1260 346 1268
rect 364 1260 366 1268
rect 374 1260 376 1268
rect 394 1260 396 1268
rect 404 1260 406 1268
rect 424 1260 426 1268
rect 434 1260 436 1268
rect 454 1260 456 1268
rect 464 1260 466 1268
rect 484 1260 486 1268
rect 494 1260 496 1268
rect 514 1260 516 1268
rect 524 1260 526 1268
rect 544 1260 546 1268
rect 554 1260 560 1268
rect 42 1258 76 1260
rect 84 1258 106 1260
rect 114 1258 136 1260
rect 144 1258 166 1260
rect 174 1258 196 1260
rect 204 1258 226 1260
rect 234 1258 256 1260
rect 264 1258 286 1260
rect 294 1258 316 1260
rect 324 1258 346 1260
rect 354 1258 376 1260
rect 384 1258 406 1260
rect 414 1258 436 1260
rect 444 1258 466 1260
rect 474 1258 496 1260
rect 504 1258 526 1260
rect 534 1258 560 1260
rect 42 1250 46 1258
rect 54 1250 56 1258
rect 64 1250 66 1258
rect 84 1250 86 1258
rect 94 1250 96 1258
rect 114 1250 116 1258
rect 124 1250 126 1258
rect 144 1250 146 1258
rect 154 1250 156 1258
rect 174 1250 176 1258
rect 184 1250 186 1258
rect 204 1250 206 1258
rect 214 1250 216 1258
rect 234 1250 236 1258
rect 244 1250 246 1258
rect 264 1250 266 1258
rect 274 1250 276 1258
rect 294 1250 296 1258
rect 304 1250 306 1258
rect 324 1250 326 1258
rect 334 1250 336 1258
rect 354 1250 356 1258
rect 364 1250 366 1258
rect 384 1250 386 1258
rect 394 1250 396 1258
rect 414 1250 416 1258
rect 424 1250 426 1258
rect 444 1250 446 1258
rect 454 1250 456 1258
rect 474 1250 476 1258
rect 484 1250 486 1258
rect 504 1250 506 1258
rect 514 1250 516 1258
rect 534 1250 536 1258
rect 544 1250 546 1258
rect 554 1250 560 1258
rect 42 1248 76 1250
rect 84 1248 106 1250
rect 114 1248 136 1250
rect 144 1248 166 1250
rect 174 1248 196 1250
rect 204 1248 226 1250
rect 234 1248 256 1250
rect 264 1248 286 1250
rect 294 1248 316 1250
rect 324 1248 346 1250
rect 354 1248 376 1250
rect 384 1248 406 1250
rect 414 1248 436 1250
rect 444 1248 466 1250
rect 474 1248 496 1250
rect 504 1248 526 1250
rect 534 1248 560 1250
rect 42 1240 46 1248
rect 54 1240 56 1248
rect 64 1240 66 1248
rect 74 1240 76 1248
rect 94 1240 96 1248
rect 104 1240 106 1248
rect 124 1240 126 1248
rect 134 1240 136 1248
rect 154 1240 156 1248
rect 164 1240 166 1248
rect 184 1240 186 1248
rect 194 1240 196 1248
rect 214 1240 216 1248
rect 224 1240 226 1248
rect 244 1240 246 1248
rect 254 1240 256 1248
rect 274 1240 276 1248
rect 284 1240 286 1248
rect 304 1240 306 1248
rect 314 1240 316 1248
rect 334 1240 336 1248
rect 344 1240 346 1248
rect 364 1240 366 1248
rect 374 1240 376 1248
rect 394 1240 396 1248
rect 404 1240 406 1248
rect 424 1240 426 1248
rect 434 1240 436 1248
rect 454 1240 456 1248
rect 464 1240 466 1248
rect 484 1240 486 1248
rect 494 1240 496 1248
rect 514 1240 516 1248
rect 524 1240 526 1248
rect 544 1240 546 1248
rect 554 1240 560 1248
rect 42 1238 76 1240
rect 84 1238 106 1240
rect 114 1238 136 1240
rect 144 1238 166 1240
rect 174 1238 196 1240
rect 204 1238 226 1240
rect 234 1238 256 1240
rect 264 1238 286 1240
rect 294 1238 316 1240
rect 324 1238 346 1240
rect 354 1238 376 1240
rect 384 1238 406 1240
rect 414 1238 436 1240
rect 444 1238 466 1240
rect 474 1238 496 1240
rect 504 1238 526 1240
rect 534 1238 560 1240
rect 42 1230 46 1238
rect 54 1230 56 1238
rect 64 1230 66 1238
rect 84 1230 86 1238
rect 94 1230 96 1238
rect 114 1230 116 1238
rect 124 1230 126 1238
rect 144 1230 146 1238
rect 154 1230 156 1238
rect 174 1230 176 1238
rect 184 1230 186 1238
rect 204 1230 206 1238
rect 214 1230 216 1238
rect 234 1230 236 1238
rect 244 1230 246 1238
rect 264 1230 266 1238
rect 274 1230 276 1238
rect 294 1230 296 1238
rect 304 1230 306 1238
rect 324 1230 326 1238
rect 334 1230 336 1238
rect 354 1230 356 1238
rect 364 1230 366 1238
rect 384 1230 386 1238
rect 394 1230 396 1238
rect 414 1230 416 1238
rect 424 1230 426 1238
rect 444 1230 446 1238
rect 454 1230 456 1238
rect 474 1230 476 1238
rect 484 1230 486 1238
rect 504 1230 506 1238
rect 514 1230 516 1238
rect 534 1230 536 1238
rect 544 1230 546 1238
rect 554 1230 560 1238
rect 42 1228 76 1230
rect 84 1228 106 1230
rect 114 1228 136 1230
rect 144 1228 166 1230
rect 174 1228 196 1230
rect 204 1228 226 1230
rect 234 1228 256 1230
rect 264 1228 286 1230
rect 294 1228 316 1230
rect 324 1228 346 1230
rect 354 1228 376 1230
rect 384 1228 406 1230
rect 414 1228 436 1230
rect 444 1228 466 1230
rect 474 1228 496 1230
rect 504 1228 526 1230
rect 534 1228 560 1230
rect 42 1220 46 1228
rect 54 1220 56 1228
rect 64 1220 66 1228
rect 74 1220 76 1228
rect 94 1220 96 1228
rect 104 1220 106 1228
rect 124 1220 126 1228
rect 134 1220 136 1228
rect 154 1220 156 1228
rect 164 1220 166 1228
rect 184 1220 186 1228
rect 194 1220 196 1228
rect 214 1220 216 1228
rect 224 1220 226 1228
rect 244 1220 246 1228
rect 254 1220 256 1228
rect 274 1220 276 1228
rect 284 1220 286 1228
rect 304 1220 306 1228
rect 314 1220 316 1228
rect 334 1220 336 1228
rect 344 1220 346 1228
rect 364 1220 366 1228
rect 374 1220 376 1228
rect 394 1220 396 1228
rect 404 1220 406 1228
rect 424 1220 426 1228
rect 434 1220 436 1228
rect 454 1220 456 1228
rect 464 1220 466 1228
rect 484 1220 486 1228
rect 494 1220 496 1228
rect 514 1220 516 1228
rect 524 1220 526 1228
rect 544 1220 546 1228
rect 554 1220 560 1228
rect 42 1218 76 1220
rect 84 1218 106 1220
rect 114 1218 136 1220
rect 144 1218 166 1220
rect 174 1218 196 1220
rect 204 1218 226 1220
rect 234 1218 256 1220
rect 264 1218 286 1220
rect 294 1218 316 1220
rect 324 1218 346 1220
rect 354 1218 376 1220
rect 384 1218 406 1220
rect 414 1218 436 1220
rect 444 1218 466 1220
rect 474 1218 496 1220
rect 504 1218 526 1220
rect 534 1218 560 1220
rect 42 1210 46 1218
rect 54 1210 56 1218
rect 64 1210 66 1218
rect 84 1210 86 1218
rect 94 1210 96 1218
rect 114 1210 116 1218
rect 124 1210 126 1218
rect 144 1210 146 1218
rect 154 1210 156 1218
rect 174 1210 176 1218
rect 184 1210 186 1218
rect 204 1210 206 1218
rect 214 1210 216 1218
rect 234 1210 236 1218
rect 244 1210 246 1218
rect 264 1210 266 1218
rect 274 1210 276 1218
rect 294 1210 296 1218
rect 304 1210 306 1218
rect 324 1210 326 1218
rect 334 1210 336 1218
rect 354 1210 356 1218
rect 364 1210 366 1218
rect 384 1210 386 1218
rect 394 1210 396 1218
rect 414 1210 416 1218
rect 424 1210 426 1218
rect 444 1210 446 1218
rect 454 1210 456 1218
rect 474 1210 476 1218
rect 484 1210 486 1218
rect 504 1210 506 1218
rect 514 1210 516 1218
rect 534 1210 536 1218
rect 544 1210 546 1218
rect 554 1210 560 1218
rect 42 1208 76 1210
rect 84 1208 106 1210
rect 114 1208 136 1210
rect 144 1208 166 1210
rect 174 1208 196 1210
rect 204 1208 226 1210
rect 234 1208 256 1210
rect 264 1208 286 1210
rect 294 1208 316 1210
rect 324 1208 346 1210
rect 354 1208 376 1210
rect 384 1208 406 1210
rect 414 1208 436 1210
rect 444 1208 466 1210
rect 474 1208 496 1210
rect 504 1208 526 1210
rect 534 1208 560 1210
rect 42 1200 46 1208
rect 54 1200 56 1208
rect 64 1200 66 1208
rect 74 1200 76 1208
rect 94 1200 96 1208
rect 104 1200 106 1208
rect 124 1200 126 1208
rect 134 1200 136 1208
rect 154 1200 156 1208
rect 164 1200 166 1208
rect 184 1200 186 1208
rect 194 1200 196 1208
rect 214 1200 216 1208
rect 224 1200 226 1208
rect 244 1200 246 1208
rect 254 1200 256 1208
rect 274 1200 276 1208
rect 284 1200 286 1208
rect 304 1200 306 1208
rect 314 1200 316 1208
rect 334 1200 336 1208
rect 344 1200 346 1208
rect 364 1200 366 1208
rect 374 1200 376 1208
rect 394 1200 396 1208
rect 404 1200 406 1208
rect 424 1200 426 1208
rect 434 1200 436 1208
rect 454 1200 456 1208
rect 464 1200 466 1208
rect 484 1200 486 1208
rect 494 1200 496 1208
rect 514 1200 516 1208
rect 524 1200 526 1208
rect 544 1200 546 1208
rect 554 1200 560 1208
rect 42 1198 76 1200
rect 84 1198 106 1200
rect 114 1198 136 1200
rect 144 1198 166 1200
rect 174 1198 196 1200
rect 204 1198 226 1200
rect 234 1198 256 1200
rect 264 1198 286 1200
rect 294 1198 316 1200
rect 324 1198 346 1200
rect 354 1198 376 1200
rect 384 1198 406 1200
rect 414 1198 436 1200
rect 444 1198 466 1200
rect 474 1198 496 1200
rect 504 1198 526 1200
rect 534 1198 560 1200
rect 42 1190 46 1198
rect 54 1190 56 1198
rect 64 1190 66 1198
rect 84 1190 86 1198
rect 94 1190 96 1198
rect 114 1190 116 1198
rect 124 1190 126 1198
rect 144 1190 146 1198
rect 154 1190 156 1198
rect 174 1190 176 1198
rect 184 1190 186 1198
rect 204 1190 206 1198
rect 214 1190 216 1198
rect 234 1190 236 1198
rect 244 1190 246 1198
rect 264 1190 266 1198
rect 274 1190 276 1198
rect 294 1190 296 1198
rect 304 1190 306 1198
rect 324 1190 326 1198
rect 334 1190 336 1198
rect 354 1190 356 1198
rect 364 1190 366 1198
rect 384 1190 386 1198
rect 394 1190 396 1198
rect 414 1190 416 1198
rect 424 1190 426 1198
rect 444 1190 446 1198
rect 454 1190 456 1198
rect 474 1190 476 1198
rect 484 1190 486 1198
rect 504 1190 506 1198
rect 514 1190 516 1198
rect 534 1190 536 1198
rect 544 1190 546 1198
rect 554 1190 560 1198
rect 42 1188 76 1190
rect 84 1188 526 1190
rect 534 1188 560 1190
rect 42 1180 46 1188
rect 54 1180 56 1188
rect 64 1180 66 1188
rect 74 1180 76 1188
rect 94 1180 506 1188
rect 514 1180 516 1188
rect 524 1180 526 1188
rect 544 1180 546 1188
rect 554 1180 560 1188
rect 42 1178 76 1180
rect 84 1178 526 1180
rect 534 1178 560 1180
rect 42 1170 46 1178
rect 54 1170 56 1178
rect 64 1170 66 1178
rect 84 1170 86 1178
rect 94 1170 96 1178
rect 114 1170 116 1178
rect 124 1170 126 1178
rect 144 1170 146 1178
rect 154 1170 156 1178
rect 174 1170 176 1178
rect 184 1170 186 1178
rect 204 1170 206 1178
rect 214 1170 216 1178
rect 234 1170 236 1178
rect 244 1170 246 1178
rect 264 1170 266 1178
rect 274 1170 276 1178
rect 294 1170 296 1178
rect 304 1170 306 1178
rect 324 1170 326 1178
rect 334 1170 336 1178
rect 354 1170 356 1178
rect 364 1170 366 1178
rect 384 1170 386 1178
rect 394 1170 396 1178
rect 414 1170 416 1178
rect 424 1170 426 1178
rect 444 1170 446 1178
rect 454 1170 456 1178
rect 474 1170 476 1178
rect 484 1170 486 1178
rect 504 1170 506 1178
rect 514 1170 516 1178
rect 534 1170 536 1178
rect 544 1170 546 1178
rect 554 1170 560 1178
rect 42 1168 76 1170
rect 84 1168 106 1170
rect 114 1168 136 1170
rect 144 1168 166 1170
rect 174 1168 196 1170
rect 204 1168 226 1170
rect 234 1168 256 1170
rect 264 1168 286 1170
rect 294 1168 316 1170
rect 324 1168 346 1170
rect 354 1168 376 1170
rect 384 1168 406 1170
rect 414 1168 436 1170
rect 444 1168 466 1170
rect 474 1168 496 1170
rect 504 1168 526 1170
rect 534 1168 560 1170
rect 42 1160 46 1168
rect 54 1160 56 1168
rect 64 1160 66 1168
rect 74 1160 76 1168
rect 94 1160 96 1168
rect 104 1160 106 1168
rect 124 1160 126 1168
rect 134 1160 136 1168
rect 154 1160 156 1168
rect 164 1160 166 1168
rect 184 1160 186 1168
rect 194 1160 196 1168
rect 214 1160 216 1168
rect 224 1160 226 1168
rect 244 1160 246 1168
rect 254 1160 256 1168
rect 274 1160 276 1168
rect 284 1160 286 1168
rect 304 1160 306 1168
rect 314 1160 316 1168
rect 334 1160 336 1168
rect 344 1160 346 1168
rect 364 1160 366 1168
rect 374 1160 376 1168
rect 394 1160 396 1168
rect 404 1160 406 1168
rect 424 1160 426 1168
rect 434 1160 436 1168
rect 454 1160 456 1168
rect 464 1160 466 1168
rect 484 1160 486 1168
rect 494 1160 496 1168
rect 514 1160 516 1168
rect 524 1160 526 1168
rect 544 1160 546 1168
rect 554 1160 560 1168
rect 42 1158 76 1160
rect 84 1158 106 1160
rect 114 1158 136 1160
rect 144 1158 166 1160
rect 174 1158 196 1160
rect 204 1158 226 1160
rect 234 1158 256 1160
rect 264 1158 286 1160
rect 294 1158 316 1160
rect 324 1158 346 1160
rect 354 1158 376 1160
rect 384 1158 406 1160
rect 414 1158 436 1160
rect 444 1158 466 1160
rect 474 1158 496 1160
rect 504 1158 526 1160
rect 534 1158 560 1160
rect 42 1150 46 1158
rect 54 1150 56 1158
rect 64 1150 66 1158
rect 84 1150 86 1158
rect 94 1150 96 1158
rect 114 1150 116 1158
rect 124 1150 126 1158
rect 144 1150 146 1158
rect 154 1150 156 1158
rect 174 1150 176 1158
rect 184 1150 186 1158
rect 204 1150 206 1158
rect 214 1150 216 1158
rect 234 1150 236 1158
rect 244 1150 246 1158
rect 264 1150 266 1158
rect 274 1150 276 1158
rect 294 1150 296 1158
rect 304 1150 306 1158
rect 324 1150 326 1158
rect 334 1150 336 1158
rect 354 1150 356 1158
rect 364 1150 366 1158
rect 384 1150 386 1158
rect 394 1150 396 1158
rect 414 1150 416 1158
rect 424 1150 426 1158
rect 444 1150 446 1158
rect 454 1150 456 1158
rect 474 1150 476 1158
rect 484 1150 486 1158
rect 504 1150 506 1158
rect 514 1150 516 1158
rect 534 1150 536 1158
rect 544 1150 546 1158
rect 554 1150 560 1158
rect 42 1148 76 1150
rect 84 1148 106 1150
rect 114 1148 136 1150
rect 144 1148 166 1150
rect 174 1148 196 1150
rect 204 1148 226 1150
rect 234 1148 256 1150
rect 264 1148 286 1150
rect 294 1148 316 1150
rect 324 1148 346 1150
rect 354 1148 376 1150
rect 384 1148 406 1150
rect 414 1148 436 1150
rect 444 1148 466 1150
rect 474 1148 496 1150
rect 504 1148 526 1150
rect 534 1148 560 1150
rect 42 1140 46 1148
rect 54 1140 56 1148
rect 64 1140 66 1148
rect 74 1140 76 1148
rect 94 1140 96 1148
rect 104 1140 106 1148
rect 124 1140 126 1148
rect 134 1140 136 1148
rect 154 1140 156 1148
rect 164 1140 166 1148
rect 184 1140 186 1148
rect 194 1140 196 1148
rect 214 1140 216 1148
rect 224 1140 226 1148
rect 244 1140 246 1148
rect 254 1140 256 1148
rect 274 1140 276 1148
rect 284 1140 286 1148
rect 304 1140 306 1148
rect 314 1140 316 1148
rect 334 1140 336 1148
rect 344 1140 346 1148
rect 364 1140 366 1148
rect 374 1140 376 1148
rect 394 1140 396 1148
rect 404 1140 406 1148
rect 424 1140 426 1148
rect 434 1140 436 1148
rect 454 1140 456 1148
rect 464 1140 466 1148
rect 484 1140 486 1148
rect 494 1140 496 1148
rect 514 1140 516 1148
rect 524 1140 526 1148
rect 544 1140 546 1148
rect 554 1140 560 1148
rect 42 1138 76 1140
rect 84 1138 106 1140
rect 114 1138 136 1140
rect 144 1138 166 1140
rect 174 1138 196 1140
rect 204 1138 226 1140
rect 234 1138 256 1140
rect 264 1138 286 1140
rect 294 1138 316 1140
rect 324 1138 346 1140
rect 354 1138 376 1140
rect 384 1138 406 1140
rect 414 1138 436 1140
rect 444 1138 466 1140
rect 474 1138 496 1140
rect 504 1138 526 1140
rect 534 1138 560 1140
rect 42 1130 46 1138
rect 54 1130 56 1138
rect 64 1130 66 1138
rect 84 1130 86 1138
rect 94 1130 96 1138
rect 114 1130 116 1138
rect 124 1130 126 1138
rect 144 1130 146 1138
rect 154 1130 156 1138
rect 174 1130 176 1138
rect 184 1130 186 1138
rect 204 1130 206 1138
rect 214 1130 216 1138
rect 234 1130 236 1138
rect 244 1130 246 1138
rect 264 1130 266 1138
rect 274 1130 276 1138
rect 294 1130 296 1138
rect 304 1130 306 1138
rect 324 1130 326 1138
rect 334 1130 336 1138
rect 354 1130 356 1138
rect 364 1130 366 1138
rect 384 1130 386 1138
rect 394 1130 396 1138
rect 414 1130 416 1138
rect 424 1130 426 1138
rect 444 1130 446 1138
rect 454 1130 456 1138
rect 474 1130 476 1138
rect 484 1130 486 1138
rect 504 1130 506 1138
rect 514 1130 516 1138
rect 534 1130 536 1138
rect 544 1130 546 1138
rect 554 1130 560 1138
rect 42 1128 76 1130
rect 84 1128 106 1130
rect 114 1128 136 1130
rect 144 1128 166 1130
rect 174 1128 196 1130
rect 204 1128 226 1130
rect 234 1128 256 1130
rect 264 1128 286 1130
rect 294 1128 316 1130
rect 324 1128 346 1130
rect 354 1128 376 1130
rect 384 1128 406 1130
rect 414 1128 436 1130
rect 444 1128 466 1130
rect 474 1128 496 1130
rect 504 1128 526 1130
rect 534 1128 560 1130
rect 42 1120 46 1128
rect 54 1120 56 1128
rect 64 1120 66 1128
rect 74 1120 76 1128
rect 94 1120 96 1128
rect 104 1120 106 1128
rect 124 1120 126 1128
rect 134 1120 136 1128
rect 154 1120 156 1128
rect 164 1120 166 1128
rect 184 1120 186 1128
rect 194 1120 196 1128
rect 214 1120 216 1128
rect 224 1120 226 1128
rect 244 1120 246 1128
rect 254 1120 256 1128
rect 274 1120 276 1128
rect 284 1120 286 1128
rect 304 1120 306 1128
rect 314 1120 316 1128
rect 334 1120 336 1128
rect 344 1120 346 1128
rect 364 1120 366 1128
rect 374 1120 376 1128
rect 394 1120 396 1128
rect 404 1120 406 1128
rect 424 1120 426 1128
rect 434 1120 436 1128
rect 454 1120 456 1128
rect 464 1120 466 1128
rect 484 1120 486 1128
rect 494 1120 496 1128
rect 42 1118 86 1120
rect 42 1110 46 1118
rect 54 1110 56 1118
rect 64 1110 66 1118
rect 74 1110 76 1118
rect 84 1110 86 1118
rect 42 1108 86 1110
rect 94 1110 100 1120
rect 500 1110 506 1120
rect 94 1108 506 1110
rect 42 1100 46 1108
rect 54 1100 56 1108
rect 64 1100 66 1108
rect 74 1100 76 1108
rect 94 1100 96 1108
rect 104 1100 106 1108
rect 124 1100 126 1108
rect 134 1100 136 1108
rect 154 1100 156 1108
rect 164 1100 166 1108
rect 184 1100 186 1108
rect 194 1100 196 1108
rect 214 1100 216 1108
rect 224 1100 226 1108
rect 244 1100 246 1108
rect 254 1100 256 1108
rect 274 1100 276 1108
rect 284 1100 286 1108
rect 304 1100 306 1108
rect 314 1100 316 1108
rect 334 1100 336 1108
rect 344 1100 346 1108
rect 364 1100 366 1108
rect 374 1100 376 1108
rect 394 1100 396 1108
rect 404 1100 406 1108
rect 424 1100 426 1108
rect 434 1100 436 1108
rect 454 1100 456 1108
rect 464 1100 466 1108
rect 484 1100 486 1108
rect 494 1100 496 1108
rect 514 1100 516 1128
rect 524 1100 526 1128
rect 544 1120 546 1128
rect 554 1120 560 1128
rect 534 1118 560 1120
rect 534 1110 536 1118
rect 544 1110 546 1118
rect 554 1110 560 1118
rect 534 1108 560 1110
rect 544 1100 546 1108
rect 554 1100 560 1108
rect 42 1098 76 1100
rect 84 1098 106 1100
rect 114 1098 136 1100
rect 144 1098 166 1100
rect 174 1098 196 1100
rect 204 1098 226 1100
rect 234 1098 256 1100
rect 264 1098 286 1100
rect 294 1098 316 1100
rect 324 1098 346 1100
rect 354 1098 376 1100
rect 384 1098 406 1100
rect 414 1098 436 1100
rect 444 1098 466 1100
rect 474 1098 496 1100
rect 504 1098 526 1100
rect 534 1098 560 1100
rect 42 1090 46 1098
rect 54 1090 56 1098
rect 64 1090 66 1098
rect 84 1090 86 1098
rect 94 1090 96 1098
rect 114 1090 116 1098
rect 124 1090 126 1098
rect 144 1090 146 1098
rect 154 1090 156 1098
rect 174 1090 176 1098
rect 184 1090 186 1098
rect 204 1090 206 1098
rect 214 1090 216 1098
rect 234 1090 236 1098
rect 244 1090 246 1098
rect 264 1090 266 1098
rect 274 1090 276 1098
rect 294 1090 296 1098
rect 304 1090 306 1098
rect 324 1090 326 1098
rect 334 1090 336 1098
rect 354 1090 356 1098
rect 364 1090 366 1098
rect 384 1090 386 1098
rect 394 1090 396 1098
rect 414 1090 416 1098
rect 424 1090 426 1098
rect 444 1090 446 1098
rect 454 1090 456 1098
rect 474 1090 476 1098
rect 484 1090 486 1098
rect 504 1090 506 1098
rect 514 1090 516 1098
rect 534 1090 536 1098
rect 544 1090 546 1098
rect 554 1090 560 1098
rect 42 1088 76 1090
rect 84 1088 106 1090
rect 114 1088 136 1090
rect 144 1088 166 1090
rect 174 1088 196 1090
rect 204 1088 226 1090
rect 234 1088 256 1090
rect 264 1088 286 1090
rect 294 1088 316 1090
rect 324 1088 346 1090
rect 354 1088 376 1090
rect 384 1088 406 1090
rect 414 1088 436 1090
rect 444 1088 466 1090
rect 474 1088 496 1090
rect 504 1088 526 1090
rect 534 1088 560 1090
rect 42 1080 46 1088
rect 54 1080 56 1088
rect 64 1080 66 1088
rect 74 1080 76 1088
rect 94 1080 96 1088
rect 104 1080 106 1088
rect 124 1080 126 1088
rect 134 1080 136 1088
rect 154 1080 156 1088
rect 164 1080 166 1088
rect 184 1080 186 1088
rect 194 1080 196 1088
rect 214 1080 216 1088
rect 224 1080 226 1088
rect 244 1080 246 1088
rect 254 1080 256 1088
rect 274 1080 276 1088
rect 284 1080 286 1088
rect 304 1080 306 1088
rect 314 1080 316 1088
rect 334 1080 336 1088
rect 344 1080 346 1088
rect 364 1080 366 1088
rect 374 1080 376 1088
rect 394 1080 396 1088
rect 404 1080 406 1088
rect 424 1080 426 1088
rect 434 1080 436 1088
rect 454 1080 456 1088
rect 464 1080 466 1088
rect 484 1080 486 1088
rect 494 1080 496 1088
rect 514 1080 516 1088
rect 524 1080 526 1088
rect 544 1080 546 1088
rect 554 1080 560 1088
rect 42 1078 76 1080
rect 84 1078 106 1080
rect 114 1078 136 1080
rect 144 1078 166 1080
rect 174 1078 196 1080
rect 204 1078 226 1080
rect 234 1078 256 1080
rect 264 1078 286 1080
rect 294 1078 316 1080
rect 324 1078 346 1080
rect 354 1078 376 1080
rect 384 1078 406 1080
rect 414 1078 436 1080
rect 444 1078 466 1080
rect 474 1078 496 1080
rect 504 1078 526 1080
rect 534 1078 560 1080
rect 42 1070 46 1078
rect 54 1070 56 1078
rect 64 1070 66 1078
rect 84 1070 86 1078
rect 94 1070 96 1078
rect 114 1070 116 1078
rect 124 1070 126 1078
rect 144 1070 146 1078
rect 154 1070 156 1078
rect 174 1070 176 1078
rect 184 1070 186 1078
rect 204 1070 206 1078
rect 214 1070 216 1078
rect 234 1070 236 1078
rect 244 1070 246 1078
rect 264 1070 266 1078
rect 274 1070 276 1078
rect 294 1070 296 1078
rect 304 1070 306 1078
rect 324 1070 326 1078
rect 334 1070 336 1078
rect 354 1070 356 1078
rect 364 1070 366 1078
rect 384 1070 386 1078
rect 394 1070 396 1078
rect 414 1070 416 1078
rect 424 1070 426 1078
rect 444 1070 446 1078
rect 454 1070 456 1078
rect 474 1070 476 1078
rect 484 1070 486 1078
rect 504 1070 506 1078
rect 514 1070 516 1078
rect 534 1070 536 1078
rect 544 1070 546 1078
rect 554 1070 560 1078
rect 42 1068 76 1070
rect 84 1068 106 1070
rect 114 1068 136 1070
rect 144 1068 166 1070
rect 174 1068 196 1070
rect 204 1068 226 1070
rect 234 1068 256 1070
rect 264 1068 286 1070
rect 294 1068 316 1070
rect 324 1068 346 1070
rect 354 1068 376 1070
rect 384 1068 406 1070
rect 414 1068 436 1070
rect 444 1068 466 1070
rect 474 1068 496 1070
rect 504 1068 526 1070
rect 534 1068 560 1070
rect 42 1060 46 1068
rect 54 1060 56 1068
rect 64 1060 66 1068
rect 74 1060 76 1068
rect 94 1060 96 1068
rect 104 1060 106 1068
rect 124 1060 126 1068
rect 134 1060 136 1068
rect 154 1060 156 1068
rect 164 1060 166 1068
rect 184 1060 186 1068
rect 194 1060 196 1068
rect 214 1060 216 1068
rect 224 1060 226 1068
rect 244 1060 246 1068
rect 254 1060 256 1068
rect 274 1060 276 1068
rect 284 1060 286 1068
rect 304 1060 306 1068
rect 314 1060 316 1068
rect 334 1060 336 1068
rect 344 1060 346 1068
rect 364 1060 366 1068
rect 374 1060 376 1068
rect 394 1060 396 1068
rect 404 1060 406 1068
rect 424 1060 426 1068
rect 434 1060 436 1068
rect 454 1060 456 1068
rect 464 1060 466 1068
rect 484 1060 486 1068
rect 494 1060 496 1068
rect 514 1060 516 1068
rect 524 1060 526 1068
rect 544 1060 546 1068
rect 554 1060 560 1068
rect 42 1058 76 1060
rect 84 1058 106 1060
rect 114 1058 136 1060
rect 144 1058 166 1060
rect 174 1058 196 1060
rect 204 1058 226 1060
rect 234 1058 256 1060
rect 264 1058 286 1060
rect 294 1058 316 1060
rect 324 1058 346 1060
rect 354 1058 376 1060
rect 384 1058 406 1060
rect 414 1058 436 1060
rect 444 1058 466 1060
rect 474 1058 496 1060
rect 504 1058 526 1060
rect 534 1058 560 1060
rect 42 1050 46 1058
rect 54 1050 56 1058
rect 64 1050 66 1058
rect 84 1050 86 1058
rect 94 1050 96 1058
rect 114 1050 116 1058
rect 124 1050 126 1058
rect 144 1050 146 1058
rect 154 1050 156 1058
rect 174 1050 176 1058
rect 184 1050 186 1058
rect 204 1050 206 1058
rect 214 1050 216 1058
rect 234 1050 236 1058
rect 244 1050 246 1058
rect 264 1050 266 1058
rect 274 1050 276 1058
rect 294 1050 296 1058
rect 304 1050 306 1058
rect 324 1050 326 1058
rect 334 1050 336 1058
rect 354 1050 356 1058
rect 364 1050 366 1058
rect 384 1050 386 1058
rect 394 1050 396 1058
rect 414 1050 416 1058
rect 424 1050 426 1058
rect 444 1050 446 1058
rect 454 1050 456 1058
rect 474 1050 476 1058
rect 484 1050 486 1058
rect 504 1050 506 1058
rect 514 1050 516 1058
rect 534 1050 536 1058
rect 544 1050 546 1058
rect 554 1050 560 1058
rect 42 1048 76 1050
rect 84 1048 106 1050
rect 114 1048 136 1050
rect 144 1048 166 1050
rect 174 1048 196 1050
rect 204 1048 226 1050
rect 234 1048 256 1050
rect 264 1048 286 1050
rect 294 1048 316 1050
rect 324 1048 346 1050
rect 354 1048 376 1050
rect 384 1048 406 1050
rect 414 1048 436 1050
rect 444 1048 466 1050
rect 474 1048 496 1050
rect 504 1048 526 1050
rect 534 1048 560 1050
rect 42 1040 46 1048
rect 54 1040 56 1048
rect 64 1040 66 1048
rect 74 1040 76 1048
rect 94 1040 96 1048
rect 104 1040 106 1048
rect 124 1040 126 1048
rect 134 1040 136 1048
rect 154 1040 156 1048
rect 164 1040 166 1048
rect 184 1040 186 1048
rect 194 1040 196 1048
rect 214 1040 216 1048
rect 224 1040 226 1048
rect 244 1040 246 1048
rect 254 1040 256 1048
rect 274 1040 276 1048
rect 284 1040 286 1048
rect 304 1040 306 1048
rect 314 1040 316 1048
rect 334 1040 336 1048
rect 344 1040 346 1048
rect 364 1040 366 1048
rect 374 1040 376 1048
rect 394 1040 396 1048
rect 404 1040 406 1048
rect 424 1040 426 1048
rect 434 1040 436 1048
rect 454 1040 456 1048
rect 464 1040 466 1048
rect 484 1040 486 1048
rect 494 1040 496 1048
rect 42 1038 76 1040
rect 84 1038 506 1040
rect 42 1030 46 1038
rect 54 1030 56 1038
rect 64 1030 66 1038
rect 84 1030 86 1038
rect 94 1030 506 1038
rect 42 1028 76 1030
rect 84 1028 506 1030
rect 42 1020 46 1028
rect 54 1020 56 1028
rect 64 1020 66 1028
rect 74 1020 76 1028
rect 94 1020 96 1028
rect 104 1020 106 1028
rect 124 1020 126 1028
rect 134 1020 136 1028
rect 154 1020 156 1028
rect 164 1020 166 1028
rect 184 1020 186 1028
rect 194 1020 196 1028
rect 214 1020 216 1028
rect 224 1020 226 1028
rect 244 1020 246 1028
rect 254 1020 256 1028
rect 274 1020 276 1028
rect 284 1020 286 1028
rect 304 1020 306 1028
rect 314 1020 316 1028
rect 334 1020 336 1028
rect 344 1020 346 1028
rect 364 1020 366 1028
rect 374 1020 376 1028
rect 394 1020 396 1028
rect 404 1020 406 1028
rect 424 1020 426 1028
rect 434 1020 436 1028
rect 454 1020 456 1028
rect 464 1020 466 1028
rect 484 1020 486 1028
rect 494 1020 496 1028
rect 514 1020 516 1048
rect 524 1020 526 1048
rect 544 1040 546 1048
rect 554 1040 560 1048
rect 534 1038 560 1040
rect 534 1030 536 1038
rect 544 1030 546 1038
rect 554 1030 560 1038
rect 534 1028 560 1030
rect 544 1020 546 1028
rect 554 1020 560 1028
rect 42 1018 76 1020
rect 84 1018 106 1020
rect 114 1018 136 1020
rect 144 1018 166 1020
rect 174 1018 196 1020
rect 204 1018 226 1020
rect 234 1018 256 1020
rect 264 1018 286 1020
rect 294 1018 316 1020
rect 324 1018 346 1020
rect 354 1018 376 1020
rect 384 1018 406 1020
rect 414 1018 436 1020
rect 444 1018 466 1020
rect 474 1018 496 1020
rect 504 1018 526 1020
rect 534 1018 560 1020
rect 42 1010 46 1018
rect 54 1010 56 1018
rect 64 1010 66 1018
rect 84 1010 86 1018
rect 94 1010 96 1018
rect 114 1010 116 1018
rect 124 1010 126 1018
rect 144 1010 146 1018
rect 154 1010 156 1018
rect 174 1010 176 1018
rect 184 1010 186 1018
rect 204 1010 206 1018
rect 214 1010 216 1018
rect 234 1010 236 1018
rect 244 1010 246 1018
rect 264 1010 266 1018
rect 274 1010 276 1018
rect 294 1010 296 1018
rect 304 1010 306 1018
rect 324 1010 326 1018
rect 334 1010 336 1018
rect 354 1010 356 1018
rect 364 1010 366 1018
rect 384 1010 386 1018
rect 394 1010 396 1018
rect 414 1010 416 1018
rect 424 1010 426 1018
rect 444 1010 446 1018
rect 454 1010 456 1018
rect 474 1010 476 1018
rect 484 1010 486 1018
rect 504 1010 506 1018
rect 514 1010 516 1018
rect 534 1010 536 1018
rect 544 1010 546 1018
rect 554 1010 560 1018
rect 42 1008 76 1010
rect 84 1008 106 1010
rect 114 1008 136 1010
rect 144 1008 166 1010
rect 174 1008 196 1010
rect 204 1008 226 1010
rect 234 1008 256 1010
rect 264 1008 286 1010
rect 294 1008 316 1010
rect 324 1008 346 1010
rect 354 1008 376 1010
rect 384 1008 406 1010
rect 414 1008 436 1010
rect 444 1008 466 1010
rect 474 1008 496 1010
rect 504 1008 526 1010
rect 534 1008 560 1010
rect 42 1000 46 1008
rect 54 1000 56 1008
rect 64 1000 66 1008
rect 74 1000 76 1008
rect 94 1000 96 1008
rect 104 1000 106 1008
rect 124 1000 126 1008
rect 134 1000 136 1008
rect 154 1000 156 1008
rect 164 1000 166 1008
rect 184 1000 186 1008
rect 194 1000 196 1008
rect 214 1000 216 1008
rect 224 1000 226 1008
rect 244 1000 246 1008
rect 254 1000 256 1008
rect 274 1000 276 1008
rect 284 1000 286 1008
rect 304 1000 306 1008
rect 314 1000 316 1008
rect 334 1000 336 1008
rect 344 1000 346 1008
rect 364 1000 366 1008
rect 374 1000 376 1008
rect 394 1000 396 1008
rect 404 1000 406 1008
rect 424 1000 426 1008
rect 434 1000 436 1008
rect 454 1000 456 1008
rect 464 1000 466 1008
rect 484 1000 486 1008
rect 494 1000 496 1008
rect 514 1000 516 1008
rect 524 1000 526 1008
rect 544 1000 546 1008
rect 554 1000 560 1008
rect 42 998 76 1000
rect 84 998 106 1000
rect 114 998 136 1000
rect 144 998 166 1000
rect 174 998 196 1000
rect 204 998 226 1000
rect 234 998 256 1000
rect 264 998 286 1000
rect 294 998 316 1000
rect 324 998 346 1000
rect 354 998 376 1000
rect 384 998 406 1000
rect 414 998 436 1000
rect 444 998 466 1000
rect 474 998 496 1000
rect 504 998 526 1000
rect 534 998 560 1000
rect 42 990 46 998
rect 54 990 56 998
rect 64 990 66 998
rect 84 990 86 998
rect 94 990 96 998
rect 114 990 116 998
rect 124 990 126 998
rect 144 990 146 998
rect 154 990 156 998
rect 174 990 176 998
rect 184 990 186 998
rect 204 990 206 998
rect 214 990 216 998
rect 234 990 236 998
rect 244 990 246 998
rect 264 990 266 998
rect 274 990 276 998
rect 294 990 296 998
rect 304 990 306 998
rect 324 990 326 998
rect 334 990 336 998
rect 354 990 356 998
rect 364 990 366 998
rect 384 990 386 998
rect 394 990 396 998
rect 414 990 416 998
rect 424 990 426 998
rect 444 990 446 998
rect 454 990 456 998
rect 474 990 476 998
rect 484 990 486 998
rect 504 990 506 998
rect 514 990 516 998
rect 534 990 536 998
rect 544 990 546 998
rect 554 990 560 998
rect 42 988 76 990
rect 84 988 106 990
rect 114 988 136 990
rect 144 988 166 990
rect 174 988 196 990
rect 204 988 226 990
rect 234 988 256 990
rect 264 988 286 990
rect 294 988 316 990
rect 324 988 346 990
rect 354 988 376 990
rect 384 988 406 990
rect 414 988 436 990
rect 444 988 466 990
rect 474 988 496 990
rect 504 988 526 990
rect 534 988 560 990
rect 42 980 46 988
rect 54 980 56 988
rect 64 980 66 988
rect 74 980 76 988
rect 94 980 96 988
rect 104 980 106 988
rect 124 980 126 988
rect 134 980 136 988
rect 154 980 156 988
rect 164 980 166 988
rect 184 980 186 988
rect 194 980 196 988
rect 214 980 216 988
rect 224 980 226 988
rect 244 980 246 988
rect 254 980 256 988
rect 274 980 276 988
rect 284 980 286 988
rect 304 980 306 988
rect 314 980 316 988
rect 334 980 336 988
rect 344 980 346 988
rect 364 980 366 988
rect 374 980 376 988
rect 394 980 396 988
rect 404 980 406 988
rect 424 980 426 988
rect 434 980 436 988
rect 454 980 456 988
rect 464 980 466 988
rect 484 980 486 988
rect 494 980 496 988
rect 514 980 516 988
rect 524 980 526 988
rect 544 980 546 988
rect 554 980 560 988
rect 42 978 76 980
rect 84 978 106 980
rect 114 978 136 980
rect 144 978 166 980
rect 174 978 196 980
rect 204 978 226 980
rect 234 978 256 980
rect 264 978 286 980
rect 294 978 316 980
rect 324 978 346 980
rect 354 978 376 980
rect 384 978 406 980
rect 414 978 436 980
rect 444 978 466 980
rect 474 978 496 980
rect 504 978 526 980
rect 534 978 560 980
rect 42 970 46 978
rect 54 970 56 978
rect 64 970 66 978
rect 84 970 86 978
rect 94 970 96 978
rect 114 970 116 978
rect 124 970 126 978
rect 144 970 146 978
rect 154 970 156 978
rect 174 970 176 978
rect 184 970 186 978
rect 204 970 206 978
rect 214 970 216 978
rect 234 970 236 978
rect 244 970 246 978
rect 264 970 266 978
rect 274 970 276 978
rect 294 970 296 978
rect 304 970 306 978
rect 324 970 326 978
rect 334 970 336 978
rect 354 970 356 978
rect 364 970 366 978
rect 384 970 386 978
rect 394 970 396 978
rect 414 970 416 978
rect 424 970 426 978
rect 444 970 446 978
rect 454 970 456 978
rect 474 970 476 978
rect 484 970 486 978
rect 504 970 506 978
rect 514 970 516 978
rect 534 970 536 978
rect 544 970 546 978
rect 554 970 560 978
rect 42 968 100 970
rect 42 960 46 968
rect 54 960 100 968
rect 500 968 560 970
rect 500 960 536 968
rect 544 960 546 968
rect 554 960 560 968
rect 42 958 560 960
rect 42 950 46 958
rect 54 950 56 958
rect 64 950 66 958
rect 84 950 86 958
rect 94 950 96 958
rect 114 950 116 958
rect 124 950 126 958
rect 144 950 146 958
rect 154 950 156 958
rect 174 950 176 958
rect 184 950 186 958
rect 204 950 206 958
rect 214 950 216 958
rect 234 950 236 958
rect 244 950 246 958
rect 264 950 266 958
rect 274 950 276 958
rect 294 950 296 958
rect 304 950 306 958
rect 324 950 326 958
rect 334 950 336 958
rect 354 950 356 958
rect 364 950 366 958
rect 384 950 386 958
rect 394 950 396 958
rect 414 950 416 958
rect 424 950 426 958
rect 444 950 446 958
rect 454 950 456 958
rect 474 950 476 958
rect 484 950 486 958
rect 504 950 506 958
rect 514 950 516 958
rect 534 950 536 958
rect 544 950 546 958
rect 554 950 560 958
rect 42 948 76 950
rect 84 948 106 950
rect 114 948 136 950
rect 144 948 166 950
rect 174 948 196 950
rect 204 948 226 950
rect 234 948 256 950
rect 264 948 286 950
rect 294 948 316 950
rect 324 948 346 950
rect 354 948 376 950
rect 384 948 406 950
rect 414 948 436 950
rect 444 948 466 950
rect 474 948 496 950
rect 504 948 526 950
rect 534 948 560 950
rect 42 940 46 948
rect 54 940 56 948
rect 64 940 66 948
rect 74 940 76 948
rect 94 940 96 948
rect 104 940 106 948
rect 124 940 126 948
rect 134 940 136 948
rect 154 940 156 948
rect 164 940 166 948
rect 184 940 186 948
rect 194 940 196 948
rect 214 940 216 948
rect 224 940 226 948
rect 244 940 246 948
rect 254 940 256 948
rect 274 940 276 948
rect 284 940 286 948
rect 304 940 306 948
rect 314 940 316 948
rect 334 940 336 948
rect 344 940 346 948
rect 364 940 366 948
rect 374 940 376 948
rect 394 940 396 948
rect 404 940 406 948
rect 424 940 426 948
rect 434 940 436 948
rect 454 940 456 948
rect 464 940 466 948
rect 484 940 486 948
rect 494 940 496 948
rect 514 940 516 948
rect 524 940 526 948
rect 544 940 546 948
rect 554 940 560 948
rect 42 938 76 940
rect 84 938 106 940
rect 114 938 136 940
rect 144 938 166 940
rect 174 938 196 940
rect 204 938 226 940
rect 234 938 256 940
rect 264 938 286 940
rect 294 938 316 940
rect 324 938 346 940
rect 354 938 376 940
rect 384 938 406 940
rect 414 938 436 940
rect 444 938 466 940
rect 474 938 496 940
rect 504 938 526 940
rect 534 938 560 940
rect 42 930 46 938
rect 54 930 56 938
rect 64 930 66 938
rect 84 930 86 938
rect 94 930 96 938
rect 114 930 116 938
rect 124 930 126 938
rect 144 930 146 938
rect 154 930 156 938
rect 174 930 176 938
rect 184 930 186 938
rect 204 930 206 938
rect 214 930 216 938
rect 234 930 236 938
rect 244 930 246 938
rect 264 930 266 938
rect 274 930 276 938
rect 294 930 296 938
rect 304 930 306 938
rect 324 930 326 938
rect 334 930 336 938
rect 354 930 356 938
rect 364 930 366 938
rect 384 930 386 938
rect 394 930 396 938
rect 414 930 416 938
rect 424 930 426 938
rect 444 930 446 938
rect 454 930 456 938
rect 474 930 476 938
rect 484 930 486 938
rect 504 930 506 938
rect 514 930 516 938
rect 534 930 536 938
rect 544 930 546 938
rect 554 930 560 938
rect 42 928 76 930
rect 84 928 106 930
rect 114 928 136 930
rect 144 928 166 930
rect 174 928 196 930
rect 204 928 226 930
rect 234 928 256 930
rect 264 928 286 930
rect 294 928 316 930
rect 324 928 346 930
rect 354 928 376 930
rect 384 928 406 930
rect 414 928 436 930
rect 444 928 466 930
rect 474 928 496 930
rect 504 928 526 930
rect 534 928 560 930
rect 42 920 46 928
rect 54 920 56 928
rect 64 920 66 928
rect 74 920 76 928
rect 94 920 96 928
rect 104 920 106 928
rect 124 920 126 928
rect 134 920 136 928
rect 154 920 156 928
rect 164 920 166 928
rect 184 920 186 928
rect 194 920 196 928
rect 214 920 216 928
rect 224 920 226 928
rect 244 920 246 928
rect 254 920 256 928
rect 274 920 276 928
rect 284 920 286 928
rect 304 920 306 928
rect 314 920 316 928
rect 334 920 336 928
rect 344 920 346 928
rect 364 920 366 928
rect 374 920 376 928
rect 394 920 396 928
rect 404 920 406 928
rect 424 920 426 928
rect 434 920 436 928
rect 454 920 456 928
rect 464 920 466 928
rect 484 920 486 928
rect 494 920 496 928
rect 514 920 516 928
rect 524 920 526 928
rect 544 920 546 928
rect 554 920 560 928
rect 42 918 76 920
rect 84 918 106 920
rect 114 918 136 920
rect 144 918 166 920
rect 174 918 196 920
rect 204 918 226 920
rect 234 918 256 920
rect 264 918 286 920
rect 294 918 316 920
rect 324 918 346 920
rect 354 918 376 920
rect 384 918 406 920
rect 414 918 436 920
rect 444 918 466 920
rect 474 918 496 920
rect 504 918 526 920
rect 534 918 560 920
rect 42 910 46 918
rect 54 910 56 918
rect 64 910 66 918
rect 84 910 86 918
rect 94 910 96 918
rect 114 910 116 918
rect 124 910 126 918
rect 144 910 146 918
rect 154 910 156 918
rect 174 910 176 918
rect 184 910 186 918
rect 204 910 206 918
rect 214 910 216 918
rect 234 910 236 918
rect 244 910 246 918
rect 264 910 266 918
rect 274 910 276 918
rect 294 910 296 918
rect 304 910 306 918
rect 324 910 326 918
rect 334 910 336 918
rect 354 910 356 918
rect 364 910 366 918
rect 384 910 386 918
rect 394 910 396 918
rect 414 910 416 918
rect 424 910 426 918
rect 444 910 446 918
rect 454 910 456 918
rect 474 910 476 918
rect 484 910 486 918
rect 504 910 506 918
rect 514 910 516 918
rect 534 910 536 918
rect 544 910 546 918
rect 554 910 560 918
rect 42 908 76 910
rect 84 908 106 910
rect 114 908 136 910
rect 144 908 166 910
rect 174 908 196 910
rect 204 908 226 910
rect 234 908 256 910
rect 264 908 286 910
rect 294 908 316 910
rect 324 908 346 910
rect 354 908 376 910
rect 384 908 406 910
rect 414 908 436 910
rect 444 908 466 910
rect 474 908 496 910
rect 504 908 526 910
rect 534 908 560 910
rect 42 900 46 908
rect 54 900 56 908
rect 64 900 66 908
rect 74 900 76 908
rect 94 900 96 908
rect 104 900 106 908
rect 124 900 126 908
rect 134 900 136 908
rect 154 900 156 908
rect 164 900 166 908
rect 184 900 186 908
rect 194 900 196 908
rect 214 900 216 908
rect 224 900 226 908
rect 244 900 246 908
rect 254 900 256 908
rect 274 900 276 908
rect 284 900 286 908
rect 304 900 306 908
rect 314 900 316 908
rect 334 900 336 908
rect 344 900 346 908
rect 364 900 366 908
rect 374 900 376 908
rect 394 900 396 908
rect 404 900 406 908
rect 424 900 426 908
rect 434 900 436 908
rect 454 900 456 908
rect 464 900 466 908
rect 484 900 486 908
rect 494 900 496 908
rect 514 900 516 908
rect 524 900 526 908
rect 544 900 546 908
rect 554 900 560 908
rect 42 898 76 900
rect 84 898 106 900
rect 114 898 136 900
rect 144 898 166 900
rect 174 898 196 900
rect 204 898 226 900
rect 234 898 256 900
rect 264 898 286 900
rect 294 898 316 900
rect 324 898 346 900
rect 354 898 376 900
rect 384 898 406 900
rect 414 898 436 900
rect 444 898 466 900
rect 474 898 496 900
rect 504 898 526 900
rect 534 898 560 900
rect 42 890 46 898
rect 54 890 56 898
rect 64 890 66 898
rect 84 890 86 898
rect 94 890 96 898
rect 114 890 116 898
rect 124 890 126 898
rect 144 890 146 898
rect 154 890 156 898
rect 174 890 176 898
rect 184 890 186 898
rect 204 890 206 898
rect 214 890 216 898
rect 234 890 236 898
rect 244 890 246 898
rect 264 890 266 898
rect 274 890 276 898
rect 294 890 296 898
rect 304 890 306 898
rect 324 890 326 898
rect 334 890 336 898
rect 354 890 356 898
rect 364 890 366 898
rect 384 890 386 898
rect 394 890 396 898
rect 414 890 416 898
rect 424 890 426 898
rect 444 890 446 898
rect 454 890 456 898
rect 474 890 476 898
rect 484 890 486 898
rect 504 890 506 898
rect 514 890 516 898
rect 534 890 536 898
rect 544 890 546 898
rect 554 890 560 898
rect 42 888 76 890
rect 84 888 106 890
rect 114 888 136 890
rect 144 888 166 890
rect 174 888 196 890
rect 204 888 226 890
rect 234 888 256 890
rect 264 888 286 890
rect 294 888 316 890
rect 324 888 346 890
rect 354 888 376 890
rect 384 888 406 890
rect 414 888 436 890
rect 444 888 466 890
rect 474 888 496 890
rect 504 888 526 890
rect 534 888 560 890
rect 42 880 46 888
rect 54 880 56 888
rect 42 878 56 880
rect 64 880 66 888
rect 74 880 76 888
rect 64 878 76 880
rect 94 880 96 888
rect 104 880 106 888
rect 94 878 106 880
rect 124 880 126 888
rect 134 880 136 888
rect 124 878 136 880
rect 154 880 156 888
rect 164 880 166 888
rect 154 878 166 880
rect 184 880 186 888
rect 194 880 196 888
rect 184 878 196 880
rect 214 880 216 888
rect 224 880 226 888
rect 214 878 226 880
rect 244 880 246 888
rect 254 880 256 888
rect 244 878 256 880
rect 274 880 276 888
rect 284 880 286 888
rect 274 878 286 880
rect 304 880 306 888
rect 314 880 316 888
rect 304 878 316 880
rect 334 880 336 888
rect 344 880 346 888
rect 334 878 346 880
rect 364 880 366 888
rect 374 880 376 888
rect 364 878 376 880
rect 394 880 396 888
rect 404 880 406 888
rect 394 878 406 880
rect 424 880 426 888
rect 434 880 436 888
rect 424 878 436 880
rect 454 880 456 888
rect 464 880 466 888
rect 454 878 466 880
rect 484 880 486 888
rect 494 880 496 888
rect 484 878 496 880
rect 514 880 516 888
rect 524 880 526 888
rect 514 878 526 880
rect 544 880 546 888
rect 554 880 560 888
rect 544 878 560 880
rect 42 870 46 878
rect 554 870 560 878
rect 42 866 560 870
rect 586 838 588 1326
rect 12 836 588 838
rect 12 828 14 836
rect 22 828 24 836
rect 42 828 44 836
rect 52 828 54 836
rect 72 828 74 836
rect 82 828 84 836
rect 102 828 104 836
rect 112 828 114 836
rect 132 828 134 836
rect 142 828 144 836
rect 162 828 164 836
rect 172 828 174 836
rect 192 828 194 836
rect 202 828 204 836
rect 222 828 224 836
rect 232 828 234 836
rect 242 828 244 836
rect 252 828 256 836
rect 264 828 266 836
rect 274 828 276 836
rect 294 828 296 836
rect 304 828 306 836
rect 324 828 326 836
rect 334 828 336 836
rect 344 828 348 836
rect 356 828 358 836
rect 366 828 368 836
rect 376 828 378 836
rect 396 828 398 836
rect 406 828 408 836
rect 426 828 428 836
rect 436 828 438 836
rect 456 828 458 836
rect 466 828 468 836
rect 486 828 488 836
rect 496 828 498 836
rect 516 828 518 836
rect 526 828 528 836
rect 546 828 548 836
rect 556 828 558 836
rect 576 828 578 836
rect 586 828 588 836
rect 596 828 600 1336
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 184 828
rect 192 826 214 828
rect 222 826 286 828
rect 294 826 316 828
rect 324 826 378 828
rect 386 826 408 828
rect 416 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 0 818 4 826
rect 12 818 14 826
rect 22 818 24 826
rect 32 818 34 826
rect 52 818 54 826
rect 62 818 64 826
rect 82 818 84 826
rect 92 818 94 826
rect 112 818 114 826
rect 122 818 124 826
rect 142 818 144 826
rect 152 818 154 826
rect 172 818 174 826
rect 182 818 184 826
rect 202 818 204 826
rect 212 818 214 826
rect 232 818 234 826
rect 242 818 244 826
rect 252 818 256 826
rect 264 818 266 826
rect 274 818 276 826
rect 284 818 286 826
rect 304 818 306 826
rect 314 818 316 826
rect 334 818 336 826
rect 344 818 348 826
rect 356 818 358 826
rect 366 818 368 826
rect 386 818 388 826
rect 396 818 398 826
rect 416 818 418 826
rect 426 818 428 826
rect 446 818 448 826
rect 456 818 458 826
rect 476 818 478 826
rect 486 818 488 826
rect 506 818 508 826
rect 516 818 518 826
rect 536 818 538 826
rect 546 818 548 826
rect 566 818 568 826
rect 576 818 578 826
rect 586 818 588 826
rect 596 818 600 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 184 818
rect 192 816 214 818
rect 222 816 286 818
rect 294 816 316 818
rect 324 816 378 818
rect 386 816 408 818
rect 416 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 0 808 4 816
rect 12 808 14 816
rect 22 808 24 816
rect 42 808 44 816
rect 52 808 54 816
rect 72 808 74 816
rect 82 808 84 816
rect 102 808 104 816
rect 112 808 114 816
rect 132 808 134 816
rect 142 808 144 816
rect 162 808 164 816
rect 172 808 174 816
rect 192 808 194 816
rect 202 808 204 816
rect 222 808 224 816
rect 232 808 234 816
rect 242 808 244 816
rect 252 808 256 816
rect 264 808 266 816
rect 274 808 276 816
rect 294 808 296 816
rect 304 808 306 816
rect 324 808 326 816
rect 334 808 336 816
rect 344 808 348 816
rect 356 808 358 816
rect 366 808 368 816
rect 376 808 378 816
rect 396 808 398 816
rect 406 808 408 816
rect 426 808 428 816
rect 436 808 438 816
rect 456 808 458 816
rect 466 808 468 816
rect 486 808 488 816
rect 496 808 498 816
rect 516 808 518 816
rect 526 808 528 816
rect 546 808 548 816
rect 556 808 558 816
rect 576 808 578 816
rect 586 808 588 816
rect 596 808 600 816
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 184 808
rect 192 806 214 808
rect 222 806 286 808
rect 294 806 316 808
rect 324 806 378 808
rect 386 806 408 808
rect 416 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 0 798 4 806
rect 12 798 14 806
rect 22 798 24 806
rect 32 798 34 806
rect 52 798 54 806
rect 62 798 64 806
rect 82 798 84 806
rect 92 798 94 806
rect 112 798 114 806
rect 122 798 124 806
rect 142 798 144 806
rect 152 798 154 806
rect 172 798 174 806
rect 182 798 184 806
rect 202 798 204 806
rect 212 798 214 806
rect 232 798 234 806
rect 242 798 244 806
rect 252 798 256 806
rect 264 798 266 806
rect 274 798 276 806
rect 284 798 286 806
rect 304 798 306 806
rect 314 798 316 806
rect 334 798 336 806
rect 344 798 348 806
rect 356 798 358 806
rect 366 798 368 806
rect 386 798 388 806
rect 396 798 398 806
rect 416 798 418 806
rect 426 798 428 806
rect 446 798 448 806
rect 456 798 458 806
rect 476 798 478 806
rect 486 798 488 806
rect 506 798 508 806
rect 516 798 518 806
rect 536 798 538 806
rect 546 798 548 806
rect 566 798 568 806
rect 576 798 578 806
rect 586 798 588 806
rect 596 798 600 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 184 798
rect 192 796 214 798
rect 222 796 286 798
rect 294 796 316 798
rect 324 796 378 798
rect 386 796 408 798
rect 416 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 0 788 4 796
rect 12 788 14 796
rect 22 788 24 796
rect 42 788 44 796
rect 52 788 54 796
rect 72 788 74 796
rect 82 788 84 796
rect 102 788 104 796
rect 112 788 114 796
rect 132 788 134 796
rect 142 788 144 796
rect 162 788 164 796
rect 172 788 174 796
rect 192 788 194 796
rect 202 788 204 796
rect 222 788 224 796
rect 232 788 234 796
rect 242 788 244 796
rect 252 788 256 796
rect 264 788 266 796
rect 274 788 276 796
rect 294 788 296 796
rect 304 788 306 796
rect 324 788 326 796
rect 334 788 336 796
rect 344 788 348 796
rect 356 788 358 796
rect 366 788 368 796
rect 376 788 378 796
rect 396 788 398 796
rect 406 788 408 796
rect 426 788 428 796
rect 436 788 438 796
rect 456 788 458 796
rect 466 788 468 796
rect 486 788 488 796
rect 496 788 498 796
rect 516 788 518 796
rect 526 788 528 796
rect 546 788 548 796
rect 556 788 558 796
rect 576 788 578 796
rect 586 788 588 796
rect 596 788 600 796
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 184 788
rect 192 786 214 788
rect 222 786 286 788
rect 294 786 316 788
rect 324 786 378 788
rect 386 786 408 788
rect 416 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 0 778 4 786
rect 12 778 14 786
rect 22 778 24 786
rect 32 778 34 786
rect 52 778 54 786
rect 62 778 64 786
rect 82 778 84 786
rect 92 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 778 114 786
rect 122 778 124 786
rect 112 776 124 778
rect 142 778 144 786
rect 152 778 154 786
rect 142 776 154 778
rect 172 778 174 786
rect 182 778 184 786
rect 172 776 184 778
rect 202 778 204 786
rect 212 778 214 786
rect 202 776 214 778
rect 232 778 234 786
rect 242 778 244 786
rect 232 776 244 778
rect 252 778 256 786
rect 264 778 266 786
rect 252 776 266 778
rect 274 778 276 786
rect 284 778 286 786
rect 274 776 286 778
rect 304 778 306 786
rect 314 778 316 786
rect 304 776 316 778
rect 334 778 336 786
rect 344 778 348 786
rect 334 776 348 778
rect 356 778 358 786
rect 366 778 368 786
rect 356 776 368 778
rect 386 778 388 786
rect 396 778 398 786
rect 386 776 398 778
rect 416 778 418 786
rect 426 778 428 786
rect 416 776 428 778
rect 446 778 448 786
rect 456 778 458 786
rect 446 776 458 778
rect 476 778 478 786
rect 486 778 488 786
rect 476 776 488 778
rect 506 778 508 786
rect 516 778 518 786
rect 536 778 538 786
rect 546 778 548 786
rect 566 778 568 786
rect 576 778 578 786
rect 586 778 588 786
rect 596 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 0 768 4 776
rect 12 768 14 776
rect 22 768 24 776
rect 42 768 44 776
rect 52 768 54 776
rect 72 768 74 776
rect 82 768 84 776
rect 252 768 256 776
rect 344 768 348 776
rect 516 768 518 776
rect 526 768 528 776
rect 546 768 548 776
rect 556 768 558 776
rect 576 768 578 776
rect 586 768 588 776
rect 596 768 600 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 4 766
rect 12 758 14 766
rect 22 758 24 766
rect 32 758 34 766
rect 52 758 54 766
rect 62 758 64 766
rect 82 758 84 766
rect 92 758 94 766
rect 112 766 124 768
rect 112 758 114 766
rect 122 758 124 766
rect 142 766 154 768
rect 142 758 144 766
rect 152 758 154 766
rect 172 766 184 768
rect 172 758 174 766
rect 182 758 184 766
rect 202 766 214 768
rect 202 758 204 766
rect 212 758 214 766
rect 232 766 244 768
rect 232 758 234 766
rect 242 758 244 766
rect 252 766 266 768
rect 252 758 256 766
rect 264 758 266 766
rect 274 766 286 768
rect 274 758 276 766
rect 284 758 286 766
rect 304 766 316 768
rect 304 758 306 766
rect 314 758 316 766
rect 334 766 348 768
rect 334 758 336 766
rect 344 758 348 766
rect 356 766 368 768
rect 356 758 358 766
rect 366 758 368 766
rect 386 766 398 768
rect 386 758 388 766
rect 396 758 398 766
rect 416 766 428 768
rect 416 758 418 766
rect 426 758 428 766
rect 446 766 458 768
rect 446 758 448 766
rect 456 758 458 766
rect 476 766 488 768
rect 476 758 478 766
rect 486 758 488 766
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 508 766
rect 516 758 518 766
rect 536 758 538 766
rect 546 758 548 766
rect 566 758 568 766
rect 576 758 578 766
rect 586 758 588 766
rect 596 758 600 766
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 184 758
rect 192 756 214 758
rect 222 756 286 758
rect 294 756 316 758
rect 324 756 378 758
rect 386 756 408 758
rect 416 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 0 748 4 756
rect 12 748 14 756
rect 22 748 24 756
rect 42 748 44 756
rect 52 748 54 756
rect 72 748 74 756
rect 82 748 84 756
rect 102 748 104 756
rect 112 748 114 756
rect 132 748 134 756
rect 142 748 144 756
rect 162 748 164 756
rect 172 748 174 756
rect 192 748 194 756
rect 202 748 204 756
rect 222 748 224 756
rect 232 748 234 756
rect 242 748 244 756
rect 252 748 256 756
rect 264 748 266 756
rect 274 748 276 756
rect 294 748 296 756
rect 304 748 306 756
rect 324 748 326 756
rect 334 748 336 756
rect 344 748 348 756
rect 356 748 358 756
rect 366 748 368 756
rect 376 748 378 756
rect 396 748 398 756
rect 406 748 408 756
rect 426 748 428 756
rect 436 748 438 756
rect 456 748 458 756
rect 466 748 468 756
rect 486 748 488 756
rect 496 748 498 756
rect 516 748 518 756
rect 526 748 528 756
rect 546 748 548 756
rect 556 748 558 756
rect 576 748 578 756
rect 586 748 588 756
rect 596 748 600 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 184 748
rect 192 746 214 748
rect 222 746 286 748
rect 294 746 316 748
rect 324 746 378 748
rect 386 746 408 748
rect 416 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 0 738 4 746
rect 12 738 14 746
rect 22 738 24 746
rect 32 738 34 746
rect 52 738 54 746
rect 62 738 64 746
rect 82 738 84 746
rect 92 738 94 746
rect 112 738 114 746
rect 122 738 124 746
rect 142 738 144 746
rect 152 738 154 746
rect 172 738 174 746
rect 182 738 184 746
rect 202 738 204 746
rect 212 738 214 746
rect 232 738 234 746
rect 242 738 244 746
rect 252 738 256 746
rect 264 738 266 746
rect 274 738 276 746
rect 284 738 286 746
rect 304 738 306 746
rect 314 738 316 746
rect 334 738 336 746
rect 344 738 348 746
rect 356 738 358 746
rect 366 738 368 746
rect 386 738 388 746
rect 396 738 398 746
rect 416 738 418 746
rect 426 738 428 746
rect 446 738 448 746
rect 456 738 458 746
rect 476 738 478 746
rect 486 738 488 746
rect 506 738 508 746
rect 516 738 518 746
rect 536 738 538 746
rect 546 738 548 746
rect 566 738 568 746
rect 576 738 578 746
rect 586 738 588 746
rect 596 738 600 746
rect 0 737 214 738
rect 0 736 42 737
rect 0 728 4 736
rect 12 728 14 736
rect 22 728 24 736
rect 32 728 42 736
rect 0 727 42 728
rect 0 726 214 727
rect 222 736 286 738
rect 294 736 316 738
rect 324 736 378 738
rect 222 728 224 736
rect 232 728 234 736
rect 242 728 244 736
rect 252 728 256 736
rect 264 728 266 736
rect 274 728 276 736
rect 294 728 296 736
rect 304 728 306 736
rect 324 728 326 736
rect 334 728 336 736
rect 344 728 348 736
rect 356 728 358 736
rect 366 728 368 736
rect 376 728 378 736
rect 222 726 286 728
rect 294 726 316 728
rect 324 726 378 728
rect 560 736 600 738
rect 560 728 568 736
rect 576 728 578 736
rect 586 728 588 736
rect 596 728 600 736
rect 386 726 600 728
rect 0 718 4 726
rect 12 718 14 726
rect 22 718 24 726
rect 32 718 34 726
rect 52 718 54 726
rect 62 718 64 726
rect 82 718 84 726
rect 92 718 94 726
rect 112 718 114 726
rect 122 718 124 726
rect 142 718 144 726
rect 152 718 154 726
rect 172 718 174 726
rect 182 718 184 726
rect 202 718 204 726
rect 212 718 214 726
rect 232 718 234 726
rect 242 718 244 726
rect 252 718 256 726
rect 264 718 266 726
rect 274 718 276 726
rect 284 718 286 726
rect 304 718 306 726
rect 314 718 316 726
rect 334 718 336 726
rect 344 718 348 726
rect 356 718 358 726
rect 366 718 368 726
rect 386 718 388 726
rect 396 718 398 726
rect 416 718 418 726
rect 426 718 428 726
rect 446 718 448 726
rect 456 718 458 726
rect 476 718 478 726
rect 486 718 488 726
rect 506 718 508 726
rect 516 718 518 726
rect 536 718 538 726
rect 546 718 548 726
rect 566 718 568 726
rect 576 718 578 726
rect 586 718 588 726
rect 596 718 600 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 184 718
rect 192 716 214 718
rect 222 716 286 718
rect 294 716 316 718
rect 324 716 378 718
rect 386 716 408 718
rect 416 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 0 708 4 716
rect 12 708 14 716
rect 22 708 24 716
rect 42 708 44 716
rect 52 708 54 716
rect 72 708 74 716
rect 82 708 84 716
rect 102 708 104 716
rect 112 708 114 716
rect 132 708 134 716
rect 142 708 144 716
rect 162 708 164 716
rect 172 708 174 716
rect 192 708 194 716
rect 202 708 204 716
rect 222 708 224 716
rect 232 708 234 716
rect 242 708 244 716
rect 252 708 256 716
rect 264 708 266 716
rect 274 708 276 716
rect 294 708 296 716
rect 304 708 306 716
rect 324 708 326 716
rect 334 708 336 716
rect 344 708 348 716
rect 356 708 358 716
rect 366 708 368 716
rect 376 708 378 716
rect 396 708 398 716
rect 406 708 408 716
rect 426 708 428 716
rect 436 708 438 716
rect 456 708 458 716
rect 466 708 468 716
rect 486 708 488 716
rect 496 708 498 716
rect 516 708 518 716
rect 526 708 528 716
rect 546 708 548 716
rect 556 708 558 716
rect 576 708 578 716
rect 586 708 588 716
rect 596 708 600 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 184 708
rect 192 706 214 708
rect 222 706 286 708
rect 294 706 316 708
rect 324 706 378 708
rect 386 706 408 708
rect 416 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 0 698 4 706
rect 12 698 14 706
rect 22 698 24 706
rect 32 698 34 706
rect 52 698 54 706
rect 62 698 64 706
rect 82 698 84 706
rect 92 698 94 706
rect 112 698 114 706
rect 122 698 124 706
rect 142 698 144 706
rect 152 698 154 706
rect 172 698 174 706
rect 182 698 184 706
rect 202 698 204 706
rect 212 698 214 706
rect 232 698 234 706
rect 242 698 244 706
rect 252 698 256 706
rect 264 698 266 706
rect 274 698 276 706
rect 284 698 286 706
rect 304 698 306 706
rect 314 698 316 706
rect 334 698 336 706
rect 344 698 348 706
rect 356 698 358 706
rect 366 698 368 706
rect 386 698 388 706
rect 396 698 398 706
rect 416 698 418 706
rect 426 698 428 706
rect 446 698 448 706
rect 456 698 458 706
rect 476 698 478 706
rect 486 698 488 706
rect 506 698 508 706
rect 516 698 518 706
rect 536 698 538 706
rect 546 698 548 706
rect 566 698 568 706
rect 576 698 578 706
rect 586 698 588 706
rect 596 698 600 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 184 698
rect 192 696 214 698
rect 222 696 286 698
rect 294 696 316 698
rect 324 696 378 698
rect 386 696 408 698
rect 416 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 0 688 4 696
rect 12 688 14 696
rect 22 688 24 696
rect 42 688 44 696
rect 52 688 54 696
rect 72 688 74 696
rect 82 688 84 696
rect 102 688 104 696
rect 112 688 114 696
rect 132 688 134 696
rect 142 688 144 696
rect 162 688 164 696
rect 172 688 174 696
rect 192 688 194 696
rect 202 688 204 696
rect 222 688 224 696
rect 232 688 234 696
rect 242 688 244 696
rect 252 688 256 696
rect 264 688 266 696
rect 274 688 276 696
rect 294 688 296 696
rect 304 688 306 696
rect 324 688 326 696
rect 334 688 336 696
rect 344 688 348 696
rect 356 688 358 696
rect 366 688 368 696
rect 376 688 378 696
rect 396 688 398 696
rect 406 688 408 696
rect 426 688 428 696
rect 436 688 438 696
rect 456 688 458 696
rect 466 688 468 696
rect 486 688 488 696
rect 496 688 498 696
rect 516 688 518 696
rect 526 688 528 696
rect 546 688 548 696
rect 556 688 558 696
rect 576 688 578 696
rect 586 688 588 696
rect 596 688 600 696
rect 0 644 4 652
rect 12 644 14 652
rect 22 644 24 652
rect 42 644 44 652
rect 52 644 54 652
rect 72 644 74 652
rect 82 644 84 652
rect 102 644 104 652
rect 112 644 114 652
rect 132 644 134 652
rect 142 644 144 652
rect 162 644 164 652
rect 172 644 174 652
rect 192 644 194 652
rect 202 644 204 652
rect 222 644 224 652
rect 232 644 234 652
rect 242 644 244 652
rect 252 644 256 652
rect 264 644 266 652
rect 274 644 276 652
rect 294 644 296 652
rect 304 644 306 652
rect 324 644 326 652
rect 334 644 336 652
rect 344 644 348 652
rect 356 644 358 652
rect 366 644 368 652
rect 376 644 378 652
rect 396 644 398 652
rect 406 644 408 652
rect 426 644 428 652
rect 436 644 438 652
rect 456 644 458 652
rect 466 644 468 652
rect 486 644 488 652
rect 496 644 498 652
rect 516 644 518 652
rect 526 644 528 652
rect 546 644 548 652
rect 556 644 558 652
rect 576 644 578 652
rect 586 644 588 652
rect 596 644 600 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 192 642 214 644
rect 222 642 286 644
rect 294 642 316 644
rect 324 642 378 644
rect 386 642 408 644
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 0 634 4 642
rect 12 634 14 642
rect 22 634 24 642
rect 32 634 34 642
rect 52 634 54 642
rect 62 634 64 642
rect 82 634 84 642
rect 92 634 94 642
rect 112 634 114 642
rect 122 634 124 642
rect 142 634 144 642
rect 152 634 154 642
rect 172 634 174 642
rect 182 634 184 642
rect 202 634 204 642
rect 212 634 214 642
rect 232 634 234 642
rect 242 634 244 642
rect 252 634 256 642
rect 264 634 266 642
rect 274 634 276 642
rect 284 634 286 642
rect 304 634 306 642
rect 314 634 316 642
rect 334 634 336 642
rect 344 634 348 642
rect 356 634 358 642
rect 366 634 368 642
rect 386 634 388 642
rect 396 634 398 642
rect 416 634 418 642
rect 426 634 428 642
rect 446 634 448 642
rect 456 634 458 642
rect 476 634 478 642
rect 486 634 488 642
rect 506 634 508 642
rect 516 634 518 642
rect 536 634 538 642
rect 546 634 548 642
rect 566 634 568 642
rect 576 634 578 642
rect 586 634 588 642
rect 596 634 600 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 192 632 214 634
rect 222 632 286 634
rect 294 632 316 634
rect 324 632 378 634
rect 386 632 408 634
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 0 624 4 632
rect 12 624 14 632
rect 22 624 24 632
rect 42 624 44 632
rect 52 624 54 632
rect 72 624 74 632
rect 82 624 84 632
rect 102 624 104 632
rect 112 624 114 632
rect 132 624 134 632
rect 142 624 144 632
rect 162 624 164 632
rect 172 624 174 632
rect 192 624 194 632
rect 202 624 204 632
rect 222 624 224 632
rect 232 624 234 632
rect 242 624 244 632
rect 252 624 256 632
rect 264 624 266 632
rect 274 624 276 632
rect 294 624 296 632
rect 304 624 306 632
rect 324 624 326 632
rect 334 624 336 632
rect 344 624 348 632
rect 356 624 358 632
rect 366 624 368 632
rect 376 624 378 632
rect 396 624 398 632
rect 406 624 408 632
rect 426 624 428 632
rect 436 624 438 632
rect 456 624 458 632
rect 466 624 468 632
rect 486 624 488 632
rect 496 624 498 632
rect 516 624 518 632
rect 526 624 528 632
rect 546 624 548 632
rect 556 624 558 632
rect 576 624 578 632
rect 586 624 588 632
rect 596 624 600 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 192 622 214 624
rect 222 622 286 624
rect 294 622 316 624
rect 324 622 378 624
rect 386 622 408 624
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 0 614 4 622
rect 12 614 14 622
rect 22 614 24 622
rect 32 614 34 622
rect 52 614 54 622
rect 62 614 64 622
rect 82 614 84 622
rect 92 614 94 622
rect 112 614 114 622
rect 122 614 124 622
rect 142 614 144 622
rect 152 614 154 622
rect 172 614 174 622
rect 182 614 184 622
rect 202 614 204 622
rect 212 614 214 622
rect 232 614 234 622
rect 242 614 244 622
rect 252 614 256 622
rect 264 614 266 622
rect 274 614 276 622
rect 284 614 286 622
rect 304 614 306 622
rect 314 614 316 622
rect 334 614 336 622
rect 344 614 348 622
rect 356 614 358 622
rect 366 614 368 622
rect 386 614 388 622
rect 396 614 398 622
rect 416 614 418 622
rect 426 614 428 622
rect 446 614 448 622
rect 456 614 458 622
rect 476 614 478 622
rect 486 614 488 622
rect 506 614 508 622
rect 516 614 518 622
rect 536 614 538 622
rect 546 614 548 622
rect 566 614 568 622
rect 576 614 578 622
rect 586 614 588 622
rect 596 614 600 622
rect 0 612 214 614
rect 0 604 4 612
rect 12 604 14 612
rect 22 604 24 612
rect 32 604 40 612
rect 0 602 40 604
rect 222 612 286 614
rect 294 612 316 614
rect 324 612 378 614
rect 222 604 224 612
rect 232 604 234 612
rect 242 604 244 612
rect 252 604 256 612
rect 264 604 266 612
rect 274 604 276 612
rect 294 604 296 612
rect 304 604 306 612
rect 324 604 326 612
rect 334 604 336 612
rect 344 604 348 612
rect 356 604 358 612
rect 366 604 368 612
rect 376 604 378 612
rect 222 602 286 604
rect 294 602 316 604
rect 324 602 378 604
rect 386 612 600 614
rect 560 604 568 612
rect 576 604 578 612
rect 586 604 588 612
rect 596 604 600 612
rect 560 602 600 604
rect 0 594 4 602
rect 12 594 14 602
rect 22 594 24 602
rect 32 594 34 602
rect 52 594 54 602
rect 62 594 64 602
rect 82 594 84 602
rect 92 594 94 602
rect 112 594 114 602
rect 122 594 124 602
rect 142 594 144 602
rect 152 594 154 602
rect 172 594 174 602
rect 182 594 184 602
rect 202 594 204 602
rect 212 594 214 602
rect 232 594 234 602
rect 242 594 244 602
rect 252 594 256 602
rect 264 594 266 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 192 592 214 594
rect 222 592 266 594
rect 274 594 276 602
rect 284 594 286 602
rect 274 592 286 594
rect 304 594 306 602
rect 314 594 316 602
rect 304 592 316 594
rect 334 594 336 602
rect 344 594 348 602
rect 356 594 358 602
rect 366 594 368 602
rect 386 594 388 602
rect 396 594 398 602
rect 416 594 418 602
rect 426 594 428 602
rect 446 594 448 602
rect 456 594 458 602
rect 476 594 478 602
rect 486 594 488 602
rect 506 594 508 602
rect 516 594 518 602
rect 536 594 538 602
rect 546 594 548 602
rect 566 594 568 602
rect 576 594 578 602
rect 586 594 588 602
rect 596 594 600 602
rect 334 592 378 594
rect 386 592 408 594
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 0 584 4 592
rect 12 584 14 592
rect 22 584 24 592
rect 42 584 44 592
rect 52 584 54 592
rect 72 584 74 592
rect 82 584 84 592
rect 102 584 104 592
rect 112 584 114 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 584
rect 132 584 134 592
rect 142 584 144 592
rect 132 582 144 584
rect 162 584 164 592
rect 172 584 174 592
rect 162 582 174 584
rect 192 584 194 592
rect 202 584 204 592
rect 192 582 204 584
rect 222 584 224 592
rect 232 584 234 592
rect 222 582 234 584
rect 242 584 244 592
rect 252 584 256 592
rect 242 582 256 584
rect 0 574 4 582
rect 12 574 14 582
rect 22 574 24 582
rect 32 574 34 582
rect 52 574 54 582
rect 62 574 64 582
rect 82 574 84 582
rect 92 574 94 582
rect 252 574 256 582
rect 344 584 348 592
rect 356 584 358 592
rect 344 582 358 584
rect 366 584 368 592
rect 376 584 378 592
rect 366 582 378 584
rect 396 584 398 592
rect 406 584 408 592
rect 396 582 408 584
rect 426 584 428 592
rect 436 584 438 592
rect 426 582 438 584
rect 456 584 458 592
rect 466 584 468 592
rect 456 582 468 584
rect 486 584 488 592
rect 496 584 498 592
rect 516 584 518 592
rect 526 584 528 592
rect 546 584 548 592
rect 556 584 558 592
rect 576 584 578 592
rect 586 584 588 592
rect 596 584 600 592
rect 486 582 498 584
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 344 574 348 582
rect 506 574 508 582
rect 516 574 518 582
rect 536 574 538 582
rect 546 574 548 582
rect 566 574 568 582
rect 576 574 578 582
rect 586 574 588 582
rect 596 574 600 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 102 572 114 574
rect 0 564 4 572
rect 12 564 14 572
rect 22 564 24 572
rect 42 564 44 572
rect 52 564 54 572
rect 72 564 74 572
rect 82 564 84 572
rect 102 564 104 572
rect 112 564 114 572
rect 132 572 144 574
rect 132 564 134 572
rect 142 564 144 572
rect 162 572 174 574
rect 162 564 164 572
rect 172 564 174 572
rect 192 572 204 574
rect 192 564 194 572
rect 202 564 204 572
rect 222 572 234 574
rect 222 564 224 572
rect 232 564 234 572
rect 242 572 256 574
rect 242 564 244 572
rect 252 564 256 572
rect 264 572 276 574
rect 264 564 266 572
rect 274 564 276 572
rect 294 572 306 574
rect 294 564 296 572
rect 304 564 306 572
rect 324 572 336 574
rect 324 564 326 572
rect 334 564 336 572
rect 344 572 358 574
rect 344 564 348 572
rect 356 564 358 572
rect 366 572 378 574
rect 366 564 368 572
rect 376 564 378 572
rect 396 572 408 574
rect 396 564 398 572
rect 406 564 408 572
rect 426 572 438 574
rect 426 564 428 572
rect 436 564 438 572
rect 456 572 468 574
rect 456 564 458 572
rect 466 564 468 572
rect 486 572 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 486 564 488 572
rect 496 564 498 572
rect 516 564 518 572
rect 526 564 528 572
rect 546 564 548 572
rect 556 564 558 572
rect 576 564 578 572
rect 586 564 588 572
rect 596 564 600 572
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 192 562 214 564
rect 222 562 286 564
rect 294 562 316 564
rect 324 562 378 564
rect 386 562 408 564
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 0 554 4 562
rect 12 554 14 562
rect 22 554 24 562
rect 32 554 34 562
rect 52 554 54 562
rect 62 554 64 562
rect 82 554 84 562
rect 92 554 94 562
rect 112 554 114 562
rect 122 554 124 562
rect 142 554 144 562
rect 152 554 154 562
rect 172 554 174 562
rect 182 554 184 562
rect 202 554 204 562
rect 212 554 214 562
rect 232 554 234 562
rect 242 554 244 562
rect 252 554 256 562
rect 264 554 266 562
rect 274 554 276 562
rect 284 554 286 562
rect 304 554 306 562
rect 314 554 316 562
rect 334 554 336 562
rect 344 554 348 562
rect 356 554 358 562
rect 366 554 368 562
rect 386 554 388 562
rect 396 554 398 562
rect 416 554 418 562
rect 426 554 428 562
rect 446 554 448 562
rect 456 554 458 562
rect 476 554 478 562
rect 486 554 488 562
rect 506 554 508 562
rect 516 554 518 562
rect 536 554 538 562
rect 546 554 548 562
rect 566 554 568 562
rect 576 554 578 562
rect 586 554 588 562
rect 596 554 600 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 192 552 214 554
rect 222 552 286 554
rect 294 552 316 554
rect 324 552 378 554
rect 386 552 408 554
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 0 544 4 552
rect 12 544 14 552
rect 22 544 24 552
rect 42 544 44 552
rect 52 544 54 552
rect 72 544 74 552
rect 82 544 84 552
rect 102 544 104 552
rect 112 544 114 552
rect 132 544 134 552
rect 142 544 144 552
rect 162 544 164 552
rect 172 544 174 552
rect 192 544 194 552
rect 202 544 204 552
rect 222 544 224 552
rect 232 544 234 552
rect 242 544 244 552
rect 252 544 256 552
rect 264 544 266 552
rect 274 544 276 552
rect 294 544 296 552
rect 304 544 306 552
rect 324 544 326 552
rect 334 544 336 552
rect 344 544 348 552
rect 356 544 358 552
rect 366 544 368 552
rect 376 544 378 552
rect 396 544 398 552
rect 406 544 408 552
rect 426 544 428 552
rect 436 544 438 552
rect 456 544 458 552
rect 466 544 468 552
rect 486 544 488 552
rect 496 544 498 552
rect 516 544 518 552
rect 526 544 528 552
rect 546 544 548 552
rect 556 544 558 552
rect 576 544 578 552
rect 586 544 588 552
rect 596 544 600 552
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 192 542 214 544
rect 222 542 286 544
rect 294 542 316 544
rect 324 542 378 544
rect 386 542 408 544
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 0 534 4 542
rect 12 534 14 542
rect 22 534 24 542
rect 32 534 34 542
rect 52 534 54 542
rect 62 534 64 542
rect 82 534 84 542
rect 92 534 94 542
rect 112 534 114 542
rect 122 534 124 542
rect 142 534 144 542
rect 152 534 154 542
rect 172 534 174 542
rect 182 534 184 542
rect 202 534 204 542
rect 212 534 214 542
rect 232 534 234 542
rect 242 534 244 542
rect 252 534 256 542
rect 264 534 266 542
rect 274 534 276 542
rect 284 534 286 542
rect 304 534 306 542
rect 314 534 316 542
rect 334 534 336 542
rect 344 534 348 542
rect 356 534 358 542
rect 366 534 368 542
rect 386 534 388 542
rect 396 534 398 542
rect 416 534 418 542
rect 426 534 428 542
rect 446 534 448 542
rect 456 534 458 542
rect 476 534 478 542
rect 486 534 488 542
rect 506 534 508 542
rect 516 534 518 542
rect 536 534 538 542
rect 546 534 548 542
rect 566 534 568 542
rect 576 534 578 542
rect 586 534 588 542
rect 596 534 600 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 192 532 214 534
rect 222 532 286 534
rect 294 532 316 534
rect 324 532 378 534
rect 386 532 408 534
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 0 524 4 532
rect 12 524 14 532
rect 22 524 24 532
rect 42 524 44 532
rect 52 524 54 532
rect 72 524 74 532
rect 82 524 84 532
rect 102 524 104 532
rect 112 524 114 532
rect 132 524 134 532
rect 142 524 144 532
rect 162 524 164 532
rect 172 524 174 532
rect 192 524 194 532
rect 202 524 204 532
rect 222 524 224 532
rect 232 524 234 532
rect 242 524 244 532
rect 252 524 256 532
rect 264 524 266 532
rect 274 524 276 532
rect 294 524 296 532
rect 304 524 306 532
rect 324 524 326 532
rect 334 524 336 532
rect 344 524 348 532
rect 356 524 358 532
rect 366 524 368 532
rect 376 524 378 532
rect 396 524 398 532
rect 406 524 408 532
rect 426 524 428 532
rect 436 524 438 532
rect 456 524 458 532
rect 466 524 468 532
rect 486 524 488 532
rect 496 524 498 532
rect 516 524 518 532
rect 526 524 528 532
rect 546 524 548 532
rect 556 524 558 532
rect 576 524 578 532
rect 586 524 588 532
rect 596 524 600 532
rect 0 516 600 524
rect 0 512 14 516
rect 0 4 4 512
rect 12 508 14 512
rect 22 508 24 516
rect 32 508 34 516
rect 42 508 44 516
rect 52 508 54 516
rect 62 508 64 516
rect 72 508 74 516
rect 82 508 84 516
rect 92 508 94 516
rect 102 508 104 516
rect 112 508 114 516
rect 122 508 124 516
rect 132 508 134 516
rect 142 508 144 516
rect 152 508 154 516
rect 162 508 164 516
rect 172 508 174 516
rect 182 508 184 516
rect 192 508 194 516
rect 202 508 204 516
rect 212 508 214 516
rect 222 508 224 516
rect 232 508 234 516
rect 242 508 244 516
rect 252 508 254 516
rect 262 508 264 516
rect 272 508 274 516
rect 282 508 284 516
rect 292 508 294 516
rect 302 508 308 516
rect 316 508 318 516
rect 326 508 328 516
rect 336 508 338 516
rect 346 508 348 516
rect 356 508 358 516
rect 366 508 368 516
rect 376 508 378 516
rect 386 508 388 516
rect 396 508 398 516
rect 406 508 408 516
rect 416 508 418 516
rect 426 508 428 516
rect 436 508 438 516
rect 446 508 448 516
rect 456 508 458 516
rect 466 508 468 516
rect 476 508 478 516
rect 486 508 488 516
rect 496 508 498 516
rect 506 508 508 516
rect 516 508 518 516
rect 526 508 528 516
rect 536 508 538 516
rect 546 508 548 516
rect 556 508 558 516
rect 566 508 568 516
rect 576 508 578 516
rect 586 512 600 516
rect 12 506 588 508
rect 12 14 14 506
rect 30 488 570 490
rect 30 460 32 488
rect 30 458 42 460
rect 30 450 32 458
rect 40 450 42 458
rect 50 458 62 460
rect 50 450 52 458
rect 60 450 62 458
rect 80 458 92 460
rect 80 450 82 458
rect 90 450 92 458
rect 110 458 122 460
rect 110 450 112 458
rect 120 450 122 458
rect 140 458 152 460
rect 140 450 142 458
rect 150 450 152 458
rect 170 458 182 460
rect 170 450 172 458
rect 180 450 182 458
rect 200 458 212 460
rect 200 450 202 458
rect 210 450 212 458
rect 230 458 242 460
rect 230 450 232 458
rect 240 450 242 458
rect 260 458 272 460
rect 260 450 262 458
rect 270 450 272 458
rect 290 458 302 460
rect 290 450 292 458
rect 300 450 302 458
rect 320 458 332 460
rect 320 450 322 458
rect 330 450 332 458
rect 350 458 362 460
rect 350 450 352 458
rect 360 450 362 458
rect 380 458 392 460
rect 380 450 382 458
rect 390 450 392 458
rect 410 458 422 460
rect 410 450 412 458
rect 420 450 422 458
rect 440 458 452 460
rect 440 450 442 458
rect 450 450 452 458
rect 470 458 482 460
rect 470 450 472 458
rect 480 450 482 458
rect 500 458 512 460
rect 500 450 502 458
rect 510 450 512 458
rect 530 458 542 460
rect 530 450 532 458
rect 540 450 542 458
rect 560 458 570 460
rect 560 450 562 458
rect 30 448 62 450
rect 70 448 92 450
rect 100 448 122 450
rect 130 448 152 450
rect 160 448 182 450
rect 190 448 212 450
rect 220 448 242 450
rect 250 448 272 450
rect 280 448 302 450
rect 310 448 332 450
rect 340 448 362 450
rect 370 448 392 450
rect 400 448 422 450
rect 430 448 452 450
rect 460 448 482 450
rect 490 448 512 450
rect 520 448 542 450
rect 550 448 570 450
rect 30 440 32 448
rect 40 440 42 448
rect 50 440 52 448
rect 70 440 72 448
rect 80 440 82 448
rect 100 440 102 448
rect 110 440 112 448
rect 130 440 132 448
rect 140 440 142 448
rect 160 440 162 448
rect 170 440 172 448
rect 190 440 192 448
rect 200 440 202 448
rect 220 440 222 448
rect 230 440 232 448
rect 250 440 252 448
rect 260 440 262 448
rect 280 440 282 448
rect 290 440 292 448
rect 310 440 312 448
rect 320 440 322 448
rect 340 440 342 448
rect 350 440 352 448
rect 370 440 372 448
rect 380 440 382 448
rect 400 440 402 448
rect 410 440 412 448
rect 430 440 432 448
rect 440 440 442 448
rect 460 440 462 448
rect 470 440 472 448
rect 490 440 492 448
rect 500 440 502 448
rect 520 440 522 448
rect 530 440 532 448
rect 550 440 552 448
rect 560 440 562 448
rect 30 438 62 440
rect 70 438 92 440
rect 100 438 122 440
rect 130 438 152 440
rect 160 438 182 440
rect 190 438 212 440
rect 220 438 242 440
rect 250 438 272 440
rect 280 438 302 440
rect 310 438 332 440
rect 340 438 362 440
rect 370 438 392 440
rect 400 438 422 440
rect 430 438 452 440
rect 460 438 482 440
rect 490 438 512 440
rect 520 438 542 440
rect 550 438 570 440
rect 30 430 32 438
rect 40 430 42 438
rect 50 430 52 438
rect 60 430 62 438
rect 80 430 82 438
rect 90 430 92 438
rect 110 430 112 438
rect 120 430 122 438
rect 140 430 142 438
rect 150 430 152 438
rect 170 430 172 438
rect 180 430 182 438
rect 200 430 202 438
rect 210 430 212 438
rect 230 430 232 438
rect 240 430 242 438
rect 260 430 262 438
rect 270 430 272 438
rect 290 430 292 438
rect 300 430 302 438
rect 320 430 322 438
rect 330 430 332 438
rect 350 430 352 438
rect 360 430 362 438
rect 380 430 382 438
rect 390 430 392 438
rect 410 430 412 438
rect 420 430 422 438
rect 440 430 442 438
rect 450 430 452 438
rect 470 430 472 438
rect 480 430 482 438
rect 500 430 502 438
rect 510 430 512 438
rect 530 430 532 438
rect 540 430 542 438
rect 560 430 562 438
rect 30 428 62 430
rect 70 428 92 430
rect 100 428 122 430
rect 130 428 152 430
rect 160 428 182 430
rect 190 428 212 430
rect 220 428 242 430
rect 250 428 272 430
rect 280 428 302 430
rect 310 428 332 430
rect 340 428 362 430
rect 370 428 392 430
rect 400 428 422 430
rect 430 428 452 430
rect 460 428 482 430
rect 490 428 512 430
rect 520 428 542 430
rect 550 428 570 430
rect 30 420 32 428
rect 40 420 42 428
rect 50 420 52 428
rect 70 420 72 428
rect 80 420 82 428
rect 100 420 102 428
rect 110 420 112 428
rect 130 420 132 428
rect 140 420 142 428
rect 160 420 162 428
rect 170 420 172 428
rect 190 420 192 428
rect 200 420 202 428
rect 220 420 222 428
rect 230 420 232 428
rect 250 420 252 428
rect 260 420 262 428
rect 280 420 282 428
rect 290 420 292 428
rect 310 420 312 428
rect 320 420 322 428
rect 340 420 342 428
rect 350 420 352 428
rect 370 420 372 428
rect 380 420 382 428
rect 400 420 402 428
rect 410 420 412 428
rect 430 420 432 428
rect 440 420 442 428
rect 460 420 462 428
rect 470 420 472 428
rect 490 420 492 428
rect 500 420 502 428
rect 520 420 522 428
rect 530 420 532 428
rect 550 420 552 428
rect 560 420 562 428
rect 30 418 62 420
rect 70 418 92 420
rect 100 418 122 420
rect 130 418 152 420
rect 160 418 182 420
rect 190 418 212 420
rect 220 418 242 420
rect 250 418 272 420
rect 280 418 302 420
rect 310 418 332 420
rect 340 418 362 420
rect 370 418 392 420
rect 400 418 422 420
rect 430 418 452 420
rect 460 418 482 420
rect 490 418 512 420
rect 520 418 542 420
rect 550 418 570 420
rect 30 410 32 418
rect 40 410 42 418
rect 50 410 52 418
rect 60 410 62 418
rect 80 410 82 418
rect 90 410 92 418
rect 110 410 112 418
rect 120 410 122 418
rect 140 410 142 418
rect 150 410 152 418
rect 170 410 172 418
rect 180 410 182 418
rect 200 410 202 418
rect 210 410 212 418
rect 230 410 232 418
rect 240 410 242 418
rect 260 410 262 418
rect 270 410 272 418
rect 290 410 292 418
rect 300 410 302 418
rect 320 410 322 418
rect 330 410 332 418
rect 350 410 352 418
rect 360 410 362 418
rect 380 410 382 418
rect 390 410 392 418
rect 410 410 412 418
rect 420 410 422 418
rect 440 410 442 418
rect 450 410 452 418
rect 470 410 472 418
rect 480 410 482 418
rect 500 410 502 418
rect 510 410 512 418
rect 530 410 532 418
rect 540 410 542 418
rect 560 410 562 418
rect 30 408 62 410
rect 70 408 92 410
rect 100 408 122 410
rect 130 408 152 410
rect 160 408 182 410
rect 190 408 212 410
rect 220 408 242 410
rect 250 408 272 410
rect 280 408 302 410
rect 310 408 332 410
rect 340 408 362 410
rect 370 408 392 410
rect 400 408 422 410
rect 430 408 452 410
rect 460 408 482 410
rect 490 408 512 410
rect 520 408 542 410
rect 550 408 570 410
rect 30 400 32 408
rect 40 400 42 408
rect 50 400 52 408
rect 70 400 72 408
rect 80 400 82 408
rect 100 400 102 408
rect 110 400 112 408
rect 130 400 132 408
rect 140 400 142 408
rect 160 400 162 408
rect 170 400 172 408
rect 190 400 192 408
rect 200 400 202 408
rect 220 400 222 408
rect 230 400 232 408
rect 250 400 252 408
rect 260 400 262 408
rect 280 400 282 408
rect 290 400 292 408
rect 310 400 312 408
rect 320 400 322 408
rect 340 400 342 408
rect 350 400 352 408
rect 370 400 372 408
rect 380 400 382 408
rect 400 400 402 408
rect 410 400 412 408
rect 430 400 432 408
rect 440 400 442 408
rect 460 400 462 408
rect 470 400 472 408
rect 490 400 492 408
rect 500 400 502 408
rect 520 400 522 408
rect 530 400 532 408
rect 550 400 552 408
rect 560 400 562 408
rect 30 398 62 400
rect 70 398 92 400
rect 100 398 122 400
rect 130 398 152 400
rect 160 398 182 400
rect 190 398 212 400
rect 220 398 242 400
rect 250 398 272 400
rect 280 398 302 400
rect 310 398 332 400
rect 340 398 362 400
rect 370 398 392 400
rect 400 398 422 400
rect 430 398 452 400
rect 460 398 482 400
rect 490 398 512 400
rect 520 398 542 400
rect 550 398 570 400
rect 30 370 32 398
rect 40 370 42 398
rect 50 370 52 398
rect 60 370 62 398
rect 80 370 82 398
rect 90 370 92 398
rect 110 390 112 398
rect 120 390 122 398
rect 140 390 142 398
rect 150 390 152 398
rect 170 390 172 398
rect 180 390 182 398
rect 200 390 202 398
rect 210 390 212 398
rect 230 390 232 398
rect 240 390 242 398
rect 260 390 262 398
rect 270 390 272 398
rect 290 390 292 398
rect 300 390 302 398
rect 320 390 322 398
rect 330 390 332 398
rect 350 390 352 398
rect 360 390 362 398
rect 380 390 382 398
rect 390 390 392 398
rect 410 390 412 398
rect 420 390 422 398
rect 440 390 442 398
rect 450 390 452 398
rect 470 390 472 398
rect 480 390 482 398
rect 500 380 502 398
rect 100 378 502 380
rect 110 370 112 378
rect 120 370 122 378
rect 140 370 142 378
rect 150 370 152 378
rect 170 370 172 378
rect 180 370 182 378
rect 200 370 202 378
rect 210 370 212 378
rect 230 370 232 378
rect 240 370 242 378
rect 260 370 262 378
rect 270 370 272 378
rect 290 370 292 378
rect 300 370 302 378
rect 320 370 322 378
rect 330 370 332 378
rect 350 370 352 378
rect 360 370 362 378
rect 380 370 382 378
rect 390 370 392 378
rect 410 370 412 378
rect 420 370 422 378
rect 440 370 442 378
rect 450 370 452 378
rect 470 370 472 378
rect 480 370 482 378
rect 500 370 502 378
rect 510 370 512 398
rect 530 390 532 398
rect 540 390 542 398
rect 560 390 562 398
rect 520 388 542 390
rect 550 388 570 390
rect 520 380 522 388
rect 530 380 532 388
rect 550 380 552 388
rect 560 380 562 388
rect 520 378 542 380
rect 550 378 570 380
rect 530 370 532 378
rect 540 370 542 378
rect 560 370 562 378
rect 30 368 62 370
rect 70 368 92 370
rect 100 368 122 370
rect 130 368 152 370
rect 160 368 182 370
rect 190 368 212 370
rect 220 368 242 370
rect 250 368 272 370
rect 280 368 302 370
rect 310 368 332 370
rect 340 368 362 370
rect 370 368 392 370
rect 400 368 422 370
rect 430 368 452 370
rect 460 368 482 370
rect 490 368 512 370
rect 520 368 542 370
rect 550 368 570 370
rect 30 360 32 368
rect 40 360 42 368
rect 50 360 52 368
rect 70 360 72 368
rect 80 360 82 368
rect 100 360 102 368
rect 110 360 112 368
rect 130 360 132 368
rect 140 360 142 368
rect 160 360 162 368
rect 170 360 172 368
rect 190 360 192 368
rect 200 360 202 368
rect 220 360 222 368
rect 230 360 232 368
rect 250 360 252 368
rect 260 360 262 368
rect 280 360 282 368
rect 290 360 292 368
rect 310 360 312 368
rect 320 360 322 368
rect 340 360 342 368
rect 350 360 352 368
rect 370 360 372 368
rect 380 360 382 368
rect 400 360 402 368
rect 410 360 412 368
rect 430 360 432 368
rect 440 360 442 368
rect 460 360 462 368
rect 470 360 472 368
rect 490 360 492 368
rect 500 360 502 368
rect 520 360 522 368
rect 530 360 532 368
rect 550 360 552 368
rect 560 360 562 368
rect 30 358 62 360
rect 70 358 92 360
rect 100 358 122 360
rect 130 358 152 360
rect 160 358 182 360
rect 190 358 212 360
rect 220 358 242 360
rect 250 358 272 360
rect 280 358 302 360
rect 310 358 332 360
rect 340 358 362 360
rect 370 358 392 360
rect 400 358 422 360
rect 430 358 452 360
rect 460 358 482 360
rect 490 358 512 360
rect 520 358 542 360
rect 550 358 570 360
rect 30 350 32 358
rect 40 350 42 358
rect 50 350 52 358
rect 60 350 62 358
rect 80 350 82 358
rect 90 350 92 358
rect 110 350 112 358
rect 120 350 122 358
rect 140 350 142 358
rect 150 350 152 358
rect 170 350 172 358
rect 180 350 182 358
rect 200 350 202 358
rect 210 350 212 358
rect 230 350 232 358
rect 240 350 242 358
rect 260 350 262 358
rect 270 350 272 358
rect 290 350 292 358
rect 300 350 302 358
rect 320 350 322 358
rect 330 350 332 358
rect 350 350 352 358
rect 360 350 362 358
rect 380 350 382 358
rect 390 350 392 358
rect 410 350 412 358
rect 420 350 422 358
rect 440 350 442 358
rect 450 350 452 358
rect 470 350 472 358
rect 480 350 482 358
rect 500 350 502 358
rect 510 350 512 358
rect 530 350 532 358
rect 540 350 542 358
rect 560 350 562 358
rect 30 348 62 350
rect 70 348 92 350
rect 100 348 122 350
rect 130 348 152 350
rect 160 348 182 350
rect 190 348 212 350
rect 220 348 242 350
rect 250 348 272 350
rect 280 348 302 350
rect 310 348 332 350
rect 340 348 362 350
rect 370 348 392 350
rect 400 348 422 350
rect 430 348 452 350
rect 460 348 482 350
rect 490 348 512 350
rect 520 348 542 350
rect 550 348 570 350
rect 30 340 32 348
rect 40 340 42 348
rect 50 340 52 348
rect 70 340 72 348
rect 80 340 82 348
rect 100 340 102 348
rect 110 340 112 348
rect 130 340 132 348
rect 140 340 142 348
rect 160 340 162 348
rect 170 340 172 348
rect 190 340 192 348
rect 200 340 202 348
rect 220 340 222 348
rect 230 340 232 348
rect 250 340 252 348
rect 260 340 262 348
rect 280 340 282 348
rect 290 340 292 348
rect 310 340 312 348
rect 320 340 322 348
rect 340 340 342 348
rect 350 340 352 348
rect 370 340 372 348
rect 380 340 382 348
rect 400 340 402 348
rect 410 340 412 348
rect 430 340 432 348
rect 440 340 442 348
rect 460 340 462 348
rect 470 340 472 348
rect 490 340 492 348
rect 500 340 502 348
rect 520 340 522 348
rect 530 340 532 348
rect 550 340 552 348
rect 560 340 562 348
rect 30 338 62 340
rect 70 338 92 340
rect 100 338 122 340
rect 130 338 152 340
rect 160 338 182 340
rect 190 338 212 340
rect 220 338 242 340
rect 250 338 272 340
rect 280 338 302 340
rect 310 338 332 340
rect 340 338 362 340
rect 370 338 392 340
rect 400 338 422 340
rect 430 338 452 340
rect 460 338 482 340
rect 490 338 512 340
rect 520 338 542 340
rect 550 338 570 340
rect 30 330 32 338
rect 40 330 42 338
rect 50 330 52 338
rect 60 330 62 338
rect 80 330 82 338
rect 90 330 92 338
rect 110 330 112 338
rect 120 330 122 338
rect 140 330 142 338
rect 150 330 152 338
rect 170 330 172 338
rect 180 330 182 338
rect 200 330 202 338
rect 210 330 212 338
rect 230 330 232 338
rect 240 330 242 338
rect 260 330 262 338
rect 270 330 272 338
rect 290 330 292 338
rect 300 330 302 338
rect 320 330 322 338
rect 330 330 332 338
rect 350 330 352 338
rect 360 330 362 338
rect 380 330 382 338
rect 390 330 392 338
rect 410 330 412 338
rect 420 330 422 338
rect 440 330 442 338
rect 450 330 452 338
rect 470 330 472 338
rect 480 330 482 338
rect 500 330 502 338
rect 510 330 512 338
rect 530 330 532 338
rect 540 330 542 338
rect 560 330 562 338
rect 30 328 62 330
rect 70 328 92 330
rect 100 328 122 330
rect 130 328 152 330
rect 160 328 182 330
rect 190 328 212 330
rect 220 328 242 330
rect 250 328 272 330
rect 280 328 302 330
rect 310 328 332 330
rect 340 328 362 330
rect 370 328 392 330
rect 400 328 422 330
rect 430 328 452 330
rect 460 328 482 330
rect 490 328 512 330
rect 520 328 542 330
rect 550 328 570 330
rect 30 320 32 328
rect 40 320 42 328
rect 50 320 52 328
rect 70 320 72 328
rect 80 320 82 328
rect 100 320 102 328
rect 110 320 112 328
rect 130 320 132 328
rect 140 320 142 328
rect 160 320 162 328
rect 170 320 172 328
rect 190 320 192 328
rect 200 320 202 328
rect 220 320 222 328
rect 230 320 232 328
rect 250 320 252 328
rect 260 320 262 328
rect 280 320 282 328
rect 290 320 292 328
rect 310 320 312 328
rect 320 320 322 328
rect 340 320 342 328
rect 350 320 352 328
rect 370 320 372 328
rect 380 320 382 328
rect 400 320 402 328
rect 410 320 412 328
rect 430 320 432 328
rect 440 320 442 328
rect 460 320 462 328
rect 470 320 472 328
rect 490 320 492 328
rect 500 320 502 328
rect 520 320 522 328
rect 530 320 532 328
rect 550 320 552 328
rect 560 320 562 328
rect 30 318 62 320
rect 70 318 92 320
rect 100 318 122 320
rect 130 318 152 320
rect 160 318 182 320
rect 190 318 212 320
rect 220 318 242 320
rect 250 318 272 320
rect 280 318 302 320
rect 310 318 332 320
rect 340 318 362 320
rect 370 318 392 320
rect 400 318 422 320
rect 430 318 452 320
rect 460 318 482 320
rect 490 318 512 320
rect 520 318 542 320
rect 550 318 570 320
rect 30 310 32 318
rect 40 310 42 318
rect 50 310 52 318
rect 60 310 62 318
rect 80 310 82 318
rect 90 310 92 318
rect 110 310 112 318
rect 120 310 122 318
rect 140 310 142 318
rect 150 310 152 318
rect 170 310 172 318
rect 180 310 182 318
rect 200 310 202 318
rect 210 310 212 318
rect 230 310 232 318
rect 240 310 242 318
rect 260 310 262 318
rect 270 310 272 318
rect 290 310 292 318
rect 300 310 302 318
rect 320 310 322 318
rect 330 310 332 318
rect 350 310 352 318
rect 360 310 362 318
rect 380 310 382 318
rect 390 310 392 318
rect 410 310 412 318
rect 420 310 422 318
rect 440 310 442 318
rect 450 310 452 318
rect 470 310 472 318
rect 480 310 482 318
rect 500 310 502 318
rect 510 310 512 318
rect 530 310 532 318
rect 540 310 542 318
rect 560 310 562 318
rect 30 308 62 310
rect 70 308 512 310
rect 520 308 542 310
rect 550 308 570 310
rect 30 300 32 308
rect 40 300 42 308
rect 50 300 52 308
rect 70 300 72 308
rect 80 300 82 308
rect 90 300 92 308
rect 100 300 502 308
rect 520 300 522 308
rect 530 300 532 308
rect 550 300 552 308
rect 560 300 562 308
rect 30 298 62 300
rect 70 298 512 300
rect 520 298 542 300
rect 550 298 570 300
rect 30 290 32 298
rect 40 290 42 298
rect 50 290 52 298
rect 60 290 62 298
rect 80 290 82 298
rect 90 290 92 298
rect 110 290 112 298
rect 120 290 122 298
rect 140 290 142 298
rect 150 290 152 298
rect 170 290 172 298
rect 180 290 182 298
rect 200 290 202 298
rect 210 290 212 298
rect 230 290 232 298
rect 240 290 242 298
rect 260 290 262 298
rect 270 290 272 298
rect 290 290 292 298
rect 300 290 302 298
rect 320 290 322 298
rect 330 290 332 298
rect 350 290 352 298
rect 360 290 362 298
rect 380 290 382 298
rect 390 290 392 298
rect 410 290 412 298
rect 420 290 422 298
rect 440 290 442 298
rect 450 290 452 298
rect 470 290 472 298
rect 480 290 482 298
rect 500 290 502 298
rect 510 290 512 298
rect 530 290 532 298
rect 540 290 542 298
rect 560 290 562 298
rect 30 288 62 290
rect 70 288 92 290
rect 100 288 122 290
rect 130 288 152 290
rect 160 288 182 290
rect 190 288 212 290
rect 220 288 242 290
rect 250 288 272 290
rect 280 288 302 290
rect 310 288 332 290
rect 340 288 362 290
rect 370 288 392 290
rect 400 288 422 290
rect 430 288 452 290
rect 460 288 482 290
rect 490 288 512 290
rect 520 288 542 290
rect 550 288 570 290
rect 30 280 32 288
rect 40 280 42 288
rect 50 280 52 288
rect 70 280 72 288
rect 80 280 82 288
rect 100 280 102 288
rect 110 280 112 288
rect 130 280 132 288
rect 140 280 142 288
rect 160 280 162 288
rect 170 280 172 288
rect 190 280 192 288
rect 200 280 202 288
rect 220 280 222 288
rect 230 280 232 288
rect 250 280 252 288
rect 260 280 262 288
rect 280 280 282 288
rect 290 280 292 288
rect 310 280 312 288
rect 320 280 322 288
rect 340 280 342 288
rect 350 280 352 288
rect 370 280 372 288
rect 380 280 382 288
rect 400 280 402 288
rect 410 280 412 288
rect 430 280 432 288
rect 440 280 442 288
rect 460 280 462 288
rect 470 280 472 288
rect 490 280 492 288
rect 500 280 502 288
rect 520 280 522 288
rect 530 280 532 288
rect 550 280 552 288
rect 560 280 562 288
rect 30 278 62 280
rect 70 278 92 280
rect 100 278 122 280
rect 130 278 152 280
rect 160 278 182 280
rect 190 278 212 280
rect 220 278 242 280
rect 250 278 272 280
rect 280 278 302 280
rect 310 278 332 280
rect 340 278 362 280
rect 370 278 392 280
rect 400 278 422 280
rect 430 278 452 280
rect 460 278 482 280
rect 490 278 512 280
rect 520 278 542 280
rect 550 278 570 280
rect 30 270 32 278
rect 40 270 42 278
rect 50 270 52 278
rect 60 270 62 278
rect 80 270 82 278
rect 90 270 92 278
rect 110 270 112 278
rect 120 270 122 278
rect 140 270 142 278
rect 150 270 152 278
rect 170 270 172 278
rect 180 270 182 278
rect 200 270 202 278
rect 210 270 212 278
rect 230 270 232 278
rect 240 270 242 278
rect 260 270 262 278
rect 270 270 272 278
rect 290 270 292 278
rect 300 270 302 278
rect 320 270 322 278
rect 330 270 332 278
rect 350 270 352 278
rect 360 270 362 278
rect 380 270 382 278
rect 390 270 392 278
rect 410 270 412 278
rect 420 270 422 278
rect 440 270 442 278
rect 450 270 452 278
rect 470 270 472 278
rect 480 270 482 278
rect 500 270 502 278
rect 510 270 512 278
rect 530 270 532 278
rect 540 270 542 278
rect 560 270 562 278
rect 30 268 62 270
rect 70 268 92 270
rect 100 268 122 270
rect 130 268 152 270
rect 160 268 182 270
rect 190 268 212 270
rect 220 268 242 270
rect 250 268 272 270
rect 280 268 302 270
rect 310 268 332 270
rect 340 268 362 270
rect 370 268 392 270
rect 400 268 422 270
rect 430 268 452 270
rect 460 268 482 270
rect 490 268 512 270
rect 520 268 542 270
rect 550 268 570 270
rect 30 260 32 268
rect 40 260 42 268
rect 50 260 52 268
rect 70 260 72 268
rect 80 260 82 268
rect 100 260 102 268
rect 110 260 112 268
rect 130 260 132 268
rect 140 260 142 268
rect 160 260 162 268
rect 170 260 172 268
rect 190 260 192 268
rect 200 260 202 268
rect 220 260 222 268
rect 230 260 232 268
rect 250 260 252 268
rect 260 260 262 268
rect 280 260 282 268
rect 290 260 292 268
rect 310 260 312 268
rect 320 260 322 268
rect 340 260 342 268
rect 350 260 352 268
rect 370 260 372 268
rect 380 260 382 268
rect 400 260 402 268
rect 410 260 412 268
rect 430 260 432 268
rect 440 260 442 268
rect 460 260 462 268
rect 470 260 472 268
rect 490 260 492 268
rect 500 260 502 268
rect 520 260 522 268
rect 530 260 532 268
rect 550 260 552 268
rect 560 260 562 268
rect 30 258 62 260
rect 70 258 92 260
rect 100 258 122 260
rect 130 258 152 260
rect 160 258 182 260
rect 190 258 212 260
rect 220 258 242 260
rect 250 258 272 260
rect 280 258 302 260
rect 310 258 332 260
rect 340 258 362 260
rect 370 258 392 260
rect 400 258 422 260
rect 430 258 452 260
rect 460 258 482 260
rect 490 258 512 260
rect 520 258 542 260
rect 550 258 570 260
rect 30 250 32 258
rect 40 250 42 258
rect 50 250 52 258
rect 60 250 62 258
rect 80 250 82 258
rect 90 250 92 258
rect 110 250 112 258
rect 120 250 122 258
rect 140 250 142 258
rect 150 250 152 258
rect 170 250 172 258
rect 180 250 182 258
rect 200 250 202 258
rect 210 250 212 258
rect 230 250 232 258
rect 240 250 242 258
rect 260 250 262 258
rect 270 250 272 258
rect 290 250 292 258
rect 300 250 302 258
rect 320 250 322 258
rect 330 250 332 258
rect 350 250 352 258
rect 360 250 362 258
rect 380 250 382 258
rect 390 250 392 258
rect 410 250 412 258
rect 420 250 422 258
rect 440 250 442 258
rect 450 250 452 258
rect 470 250 472 258
rect 480 250 482 258
rect 500 250 502 258
rect 510 250 512 258
rect 530 250 532 258
rect 540 250 542 258
rect 560 250 562 258
rect 30 248 62 250
rect 70 248 92 250
rect 100 248 122 250
rect 130 248 152 250
rect 160 248 182 250
rect 190 248 212 250
rect 220 248 242 250
rect 250 248 272 250
rect 280 248 302 250
rect 310 248 332 250
rect 340 248 362 250
rect 370 248 392 250
rect 400 248 422 250
rect 430 248 452 250
rect 460 248 482 250
rect 490 248 512 250
rect 520 248 542 250
rect 550 248 570 250
rect 30 240 32 248
rect 40 240 42 248
rect 50 240 52 248
rect 30 238 62 240
rect 30 230 32 238
rect 40 230 42 238
rect 50 230 52 238
rect 60 230 62 238
rect 30 228 62 230
rect 30 220 32 228
rect 40 220 42 228
rect 50 220 52 228
rect 70 220 72 248
rect 80 220 82 248
rect 100 240 102 248
rect 110 240 112 248
rect 130 240 132 248
rect 140 240 142 248
rect 160 240 162 248
rect 170 240 172 248
rect 190 240 192 248
rect 200 240 202 248
rect 220 240 222 248
rect 230 240 232 248
rect 250 240 252 248
rect 260 240 262 248
rect 280 240 282 248
rect 290 240 292 248
rect 310 240 312 248
rect 320 240 322 248
rect 340 240 342 248
rect 350 240 352 248
rect 370 240 372 248
rect 380 240 382 248
rect 400 240 402 248
rect 410 240 412 248
rect 430 240 432 248
rect 440 240 442 248
rect 460 240 462 248
rect 470 240 472 248
rect 490 240 492 248
rect 90 230 100 240
rect 500 230 502 248
rect 520 240 522 248
rect 530 240 532 248
rect 550 240 552 248
rect 560 240 562 248
rect 90 228 502 230
rect 510 238 542 240
rect 550 238 570 240
rect 510 230 512 238
rect 520 230 522 238
rect 530 230 532 238
rect 540 230 542 238
rect 560 230 562 238
rect 510 228 542 230
rect 550 228 570 230
rect 100 220 102 228
rect 110 220 112 228
rect 130 220 132 228
rect 140 220 142 228
rect 160 220 162 228
rect 170 220 172 228
rect 190 220 192 228
rect 200 220 202 228
rect 220 220 222 228
rect 230 220 232 228
rect 250 220 252 228
rect 260 220 262 228
rect 280 220 282 228
rect 290 220 292 228
rect 310 220 312 228
rect 320 220 322 228
rect 340 220 342 228
rect 350 220 352 228
rect 370 220 372 228
rect 380 220 382 228
rect 400 220 402 228
rect 410 220 412 228
rect 430 220 432 228
rect 440 220 442 228
rect 460 220 462 228
rect 470 220 472 228
rect 490 220 492 228
rect 500 220 502 228
rect 520 220 522 228
rect 530 220 532 228
rect 550 220 552 228
rect 560 220 562 228
rect 30 218 62 220
rect 70 218 92 220
rect 100 218 122 220
rect 130 218 152 220
rect 160 218 182 220
rect 190 218 212 220
rect 220 218 242 220
rect 250 218 272 220
rect 280 218 302 220
rect 310 218 332 220
rect 340 218 362 220
rect 370 218 392 220
rect 400 218 422 220
rect 430 218 452 220
rect 460 218 482 220
rect 490 218 512 220
rect 520 218 542 220
rect 550 218 570 220
rect 30 210 32 218
rect 40 210 42 218
rect 50 210 52 218
rect 60 210 62 218
rect 80 210 82 218
rect 90 210 92 218
rect 110 210 112 218
rect 120 210 122 218
rect 140 210 142 218
rect 150 210 152 218
rect 170 210 172 218
rect 180 210 182 218
rect 200 210 202 218
rect 210 210 212 218
rect 230 210 232 218
rect 240 210 242 218
rect 260 210 262 218
rect 270 210 272 218
rect 290 210 292 218
rect 300 210 302 218
rect 320 210 322 218
rect 330 210 332 218
rect 350 210 352 218
rect 360 210 362 218
rect 380 210 382 218
rect 390 210 392 218
rect 410 210 412 218
rect 420 210 422 218
rect 440 210 442 218
rect 450 210 452 218
rect 470 210 472 218
rect 480 210 482 218
rect 500 210 502 218
rect 510 210 512 218
rect 530 210 532 218
rect 540 210 542 218
rect 560 210 562 218
rect 30 208 62 210
rect 70 208 92 210
rect 100 208 122 210
rect 130 208 152 210
rect 160 208 182 210
rect 190 208 212 210
rect 220 208 242 210
rect 250 208 272 210
rect 280 208 302 210
rect 310 208 332 210
rect 340 208 362 210
rect 370 208 392 210
rect 400 208 422 210
rect 430 208 452 210
rect 460 208 482 210
rect 490 208 512 210
rect 520 208 542 210
rect 550 208 570 210
rect 30 200 32 208
rect 40 200 42 208
rect 50 200 52 208
rect 70 200 72 208
rect 80 200 82 208
rect 100 200 102 208
rect 110 200 112 208
rect 130 200 132 208
rect 140 200 142 208
rect 160 200 162 208
rect 170 200 172 208
rect 190 200 192 208
rect 200 200 202 208
rect 220 200 222 208
rect 230 200 232 208
rect 250 200 252 208
rect 260 200 262 208
rect 280 200 282 208
rect 290 200 292 208
rect 310 200 312 208
rect 320 200 322 208
rect 340 200 342 208
rect 350 200 352 208
rect 370 200 372 208
rect 380 200 382 208
rect 400 200 402 208
rect 410 200 412 208
rect 430 200 432 208
rect 440 200 442 208
rect 460 200 462 208
rect 470 200 472 208
rect 490 200 492 208
rect 500 200 502 208
rect 520 200 522 208
rect 530 200 532 208
rect 550 200 552 208
rect 560 200 562 208
rect 30 198 62 200
rect 70 198 92 200
rect 100 198 122 200
rect 130 198 152 200
rect 160 198 182 200
rect 190 198 212 200
rect 220 198 242 200
rect 250 198 272 200
rect 280 198 302 200
rect 310 198 332 200
rect 340 198 362 200
rect 370 198 392 200
rect 400 198 422 200
rect 430 198 452 200
rect 460 198 482 200
rect 490 198 512 200
rect 520 198 542 200
rect 550 198 570 200
rect 30 190 32 198
rect 40 190 42 198
rect 50 190 52 198
rect 60 190 62 198
rect 80 190 82 198
rect 90 190 92 198
rect 110 190 112 198
rect 120 190 122 198
rect 140 190 142 198
rect 150 190 152 198
rect 170 190 172 198
rect 180 190 182 198
rect 200 190 202 198
rect 210 190 212 198
rect 230 190 232 198
rect 240 190 242 198
rect 260 190 262 198
rect 270 190 272 198
rect 290 190 292 198
rect 300 190 302 198
rect 320 190 322 198
rect 330 190 332 198
rect 350 190 352 198
rect 360 190 362 198
rect 380 190 382 198
rect 390 190 392 198
rect 410 190 412 198
rect 420 190 422 198
rect 440 190 442 198
rect 450 190 452 198
rect 470 190 472 198
rect 480 190 482 198
rect 500 190 502 198
rect 510 190 512 198
rect 530 190 532 198
rect 540 190 542 198
rect 560 190 562 198
rect 30 188 62 190
rect 70 188 92 190
rect 100 188 122 190
rect 130 188 152 190
rect 160 188 182 190
rect 190 188 212 190
rect 220 188 242 190
rect 250 188 272 190
rect 280 188 302 190
rect 310 188 332 190
rect 340 188 362 190
rect 370 188 392 190
rect 400 188 422 190
rect 430 188 452 190
rect 460 188 482 190
rect 490 188 512 190
rect 520 188 542 190
rect 550 188 570 190
rect 30 180 32 188
rect 40 180 42 188
rect 50 180 52 188
rect 70 180 72 188
rect 80 180 82 188
rect 100 180 102 188
rect 110 180 112 188
rect 130 180 132 188
rect 140 180 142 188
rect 160 180 162 188
rect 170 180 172 188
rect 190 180 192 188
rect 200 180 202 188
rect 220 180 222 188
rect 230 180 232 188
rect 250 180 252 188
rect 260 180 262 188
rect 280 180 282 188
rect 290 180 292 188
rect 310 180 312 188
rect 320 180 322 188
rect 340 180 342 188
rect 350 180 352 188
rect 370 180 372 188
rect 380 180 382 188
rect 400 180 402 188
rect 410 180 412 188
rect 430 180 432 188
rect 440 180 442 188
rect 460 180 462 188
rect 470 180 472 188
rect 490 180 492 188
rect 500 180 502 188
rect 520 180 522 188
rect 530 180 532 188
rect 550 180 552 188
rect 560 180 562 188
rect 30 178 62 180
rect 70 178 92 180
rect 100 178 122 180
rect 130 178 152 180
rect 160 178 182 180
rect 190 178 212 180
rect 220 178 242 180
rect 250 178 272 180
rect 280 178 302 180
rect 310 178 332 180
rect 340 178 362 180
rect 370 178 392 180
rect 400 178 422 180
rect 430 178 452 180
rect 460 178 482 180
rect 490 178 512 180
rect 520 178 542 180
rect 550 178 570 180
rect 30 170 32 178
rect 40 170 42 178
rect 50 170 52 178
rect 60 170 62 178
rect 80 170 82 178
rect 90 170 92 178
rect 110 170 112 178
rect 120 170 122 178
rect 140 170 142 178
rect 150 170 152 178
rect 170 170 172 178
rect 180 170 182 178
rect 200 170 202 178
rect 210 170 212 178
rect 230 170 232 178
rect 240 170 242 178
rect 260 170 262 178
rect 270 170 272 178
rect 290 170 292 178
rect 300 170 302 178
rect 320 170 322 178
rect 330 170 332 178
rect 350 170 352 178
rect 360 170 362 178
rect 380 170 382 178
rect 390 170 392 178
rect 410 170 412 178
rect 420 170 422 178
rect 440 170 442 178
rect 450 170 452 178
rect 470 170 472 178
rect 480 170 482 178
rect 500 170 502 178
rect 510 170 512 178
rect 530 170 532 178
rect 540 170 542 178
rect 560 170 562 178
rect 30 168 62 170
rect 70 168 92 170
rect 100 168 122 170
rect 130 168 152 170
rect 160 168 182 170
rect 190 168 212 170
rect 220 168 242 170
rect 250 168 272 170
rect 280 168 302 170
rect 310 168 332 170
rect 340 168 362 170
rect 370 168 392 170
rect 400 168 422 170
rect 430 168 452 170
rect 460 168 482 170
rect 490 168 512 170
rect 520 168 542 170
rect 550 168 570 170
rect 30 160 32 168
rect 40 160 42 168
rect 50 160 52 168
rect 70 160 72 168
rect 80 160 82 168
rect 100 160 102 168
rect 110 160 112 168
rect 130 160 132 168
rect 140 160 142 168
rect 160 160 162 168
rect 170 160 172 168
rect 190 160 192 168
rect 200 160 202 168
rect 220 160 222 168
rect 230 160 232 168
rect 250 160 252 168
rect 260 160 262 168
rect 280 160 282 168
rect 290 160 292 168
rect 310 160 312 168
rect 320 160 322 168
rect 340 160 342 168
rect 350 160 352 168
rect 370 160 372 168
rect 380 160 382 168
rect 400 160 402 168
rect 410 160 412 168
rect 430 160 432 168
rect 440 160 442 168
rect 460 160 462 168
rect 470 160 472 168
rect 490 160 492 168
rect 500 160 502 168
rect 520 160 522 168
rect 530 160 532 168
rect 550 160 552 168
rect 560 160 562 168
rect 30 158 62 160
rect 70 158 92 160
rect 30 150 32 158
rect 40 150 42 158
rect 50 150 52 158
rect 60 150 62 158
rect 80 150 82 158
rect 90 150 92 158
rect 30 148 62 150
rect 70 148 92 150
rect 100 148 502 160
rect 510 158 542 160
rect 550 158 570 160
rect 510 150 512 158
rect 520 150 522 158
rect 530 150 532 158
rect 540 150 542 158
rect 560 150 562 158
rect 510 148 542 150
rect 550 148 570 150
rect 30 140 32 148
rect 40 140 42 148
rect 50 140 52 148
rect 70 140 72 148
rect 80 140 82 148
rect 100 140 102 148
rect 110 140 112 148
rect 130 140 132 148
rect 140 140 142 148
rect 160 140 162 148
rect 170 140 172 148
rect 190 140 192 148
rect 200 140 202 148
rect 220 140 222 148
rect 230 140 232 148
rect 250 140 252 148
rect 260 140 262 148
rect 280 140 282 148
rect 290 140 292 148
rect 310 140 312 148
rect 320 140 322 148
rect 340 140 342 148
rect 350 140 352 148
rect 370 140 372 148
rect 380 140 382 148
rect 400 140 402 148
rect 410 140 412 148
rect 430 140 432 148
rect 440 140 442 148
rect 460 140 462 148
rect 470 140 472 148
rect 490 140 492 148
rect 500 140 502 148
rect 520 140 522 148
rect 530 140 532 148
rect 550 140 552 148
rect 560 140 562 148
rect 30 138 62 140
rect 70 138 92 140
rect 100 138 122 140
rect 130 138 152 140
rect 160 138 182 140
rect 190 138 212 140
rect 220 138 242 140
rect 250 138 272 140
rect 280 138 302 140
rect 310 138 332 140
rect 340 138 362 140
rect 370 138 392 140
rect 400 138 422 140
rect 430 138 452 140
rect 460 138 482 140
rect 490 138 512 140
rect 520 138 542 140
rect 550 138 570 140
rect 30 130 32 138
rect 40 130 42 138
rect 50 130 52 138
rect 60 130 62 138
rect 80 130 82 138
rect 90 130 92 138
rect 110 130 112 138
rect 120 130 122 138
rect 140 130 142 138
rect 150 130 152 138
rect 170 130 172 138
rect 180 130 182 138
rect 200 130 202 138
rect 210 130 212 138
rect 230 130 232 138
rect 240 130 242 138
rect 260 130 262 138
rect 270 130 272 138
rect 290 130 292 138
rect 300 130 302 138
rect 320 130 322 138
rect 330 130 332 138
rect 350 130 352 138
rect 360 130 362 138
rect 380 130 382 138
rect 390 130 392 138
rect 410 130 412 138
rect 420 130 422 138
rect 440 130 442 138
rect 450 130 452 138
rect 470 130 472 138
rect 480 130 482 138
rect 500 130 502 138
rect 510 130 512 138
rect 530 130 532 138
rect 540 130 542 138
rect 560 130 562 138
rect 30 128 62 130
rect 70 128 92 130
rect 100 128 122 130
rect 130 128 152 130
rect 160 128 182 130
rect 190 128 212 130
rect 220 128 242 130
rect 250 128 272 130
rect 280 128 302 130
rect 310 128 332 130
rect 340 128 362 130
rect 370 128 392 130
rect 400 128 422 130
rect 430 128 452 130
rect 460 128 482 130
rect 490 128 512 130
rect 520 128 542 130
rect 550 128 570 130
rect 30 120 32 128
rect 40 120 42 128
rect 50 120 52 128
rect 70 120 72 128
rect 80 120 82 128
rect 100 120 102 128
rect 110 120 112 128
rect 130 120 132 128
rect 140 120 142 128
rect 160 120 162 128
rect 170 120 172 128
rect 190 120 192 128
rect 200 120 202 128
rect 220 120 222 128
rect 230 120 232 128
rect 250 120 252 128
rect 260 120 262 128
rect 280 120 282 128
rect 290 120 292 128
rect 310 120 312 128
rect 320 120 322 128
rect 340 120 342 128
rect 350 120 352 128
rect 370 120 372 128
rect 380 120 382 128
rect 400 120 402 128
rect 410 120 412 128
rect 430 120 432 128
rect 440 120 442 128
rect 460 120 462 128
rect 470 120 472 128
rect 490 120 492 128
rect 500 120 502 128
rect 520 120 522 128
rect 530 120 532 128
rect 550 120 552 128
rect 560 120 562 128
rect 30 118 62 120
rect 70 118 92 120
rect 100 118 122 120
rect 130 118 152 120
rect 160 118 182 120
rect 190 118 212 120
rect 220 118 242 120
rect 250 118 272 120
rect 280 118 302 120
rect 310 118 332 120
rect 340 118 362 120
rect 370 118 392 120
rect 400 118 422 120
rect 430 118 452 120
rect 460 118 482 120
rect 490 118 512 120
rect 520 118 542 120
rect 550 118 570 120
rect 30 110 32 118
rect 40 110 42 118
rect 50 110 52 118
rect 60 110 62 118
rect 80 110 82 118
rect 90 110 92 118
rect 110 110 112 118
rect 120 110 122 118
rect 140 110 142 118
rect 150 110 152 118
rect 170 110 172 118
rect 180 110 182 118
rect 200 110 202 118
rect 210 110 212 118
rect 230 110 232 118
rect 240 110 242 118
rect 260 110 262 118
rect 270 110 272 118
rect 290 110 292 118
rect 300 110 302 118
rect 320 110 322 118
rect 330 110 332 118
rect 350 110 352 118
rect 360 110 362 118
rect 380 110 382 118
rect 390 110 392 118
rect 410 110 412 118
rect 420 110 422 118
rect 440 110 442 118
rect 450 110 452 118
rect 470 110 472 118
rect 480 110 482 118
rect 500 110 502 118
rect 510 110 512 118
rect 530 110 532 118
rect 540 110 542 118
rect 560 110 562 118
rect 30 108 62 110
rect 70 108 92 110
rect 100 108 122 110
rect 130 108 152 110
rect 160 108 182 110
rect 190 108 212 110
rect 220 108 242 110
rect 250 108 272 110
rect 280 108 302 110
rect 310 108 332 110
rect 340 108 362 110
rect 370 108 392 110
rect 400 108 422 110
rect 430 108 452 110
rect 460 108 482 110
rect 490 108 512 110
rect 520 108 542 110
rect 550 108 570 110
rect 30 100 32 108
rect 40 100 42 108
rect 50 100 52 108
rect 70 100 72 108
rect 80 100 82 108
rect 100 100 102 108
rect 110 100 112 108
rect 130 100 132 108
rect 140 100 142 108
rect 160 100 162 108
rect 170 100 172 108
rect 190 100 192 108
rect 200 100 202 108
rect 220 100 222 108
rect 230 100 232 108
rect 250 100 252 108
rect 260 100 262 108
rect 280 100 282 108
rect 290 100 292 108
rect 310 100 312 108
rect 320 100 322 108
rect 340 100 342 108
rect 350 100 352 108
rect 370 100 372 108
rect 380 100 382 108
rect 400 100 402 108
rect 410 100 412 108
rect 430 100 432 108
rect 440 100 442 108
rect 460 100 462 108
rect 470 100 472 108
rect 490 100 492 108
rect 500 100 502 108
rect 520 100 522 108
rect 530 100 532 108
rect 550 100 552 108
rect 560 100 562 108
rect 30 98 62 100
rect 70 98 92 100
rect 100 98 122 100
rect 130 98 152 100
rect 160 98 182 100
rect 190 98 212 100
rect 220 98 242 100
rect 250 98 272 100
rect 280 98 302 100
rect 310 98 332 100
rect 340 98 362 100
rect 370 98 392 100
rect 400 98 422 100
rect 430 98 452 100
rect 460 98 482 100
rect 490 98 512 100
rect 520 98 542 100
rect 550 98 570 100
rect 30 90 32 98
rect 40 90 42 98
rect 50 90 52 98
rect 60 90 62 98
rect 80 90 82 98
rect 90 90 92 98
rect 110 90 112 98
rect 120 90 122 98
rect 140 90 142 98
rect 150 90 152 98
rect 170 90 172 98
rect 180 90 182 98
rect 200 90 202 98
rect 210 90 212 98
rect 230 90 232 98
rect 240 90 242 98
rect 260 90 262 98
rect 270 90 272 98
rect 290 90 292 98
rect 300 90 302 98
rect 320 90 322 98
rect 330 90 332 98
rect 350 90 352 98
rect 360 90 362 98
rect 380 90 382 98
rect 390 90 392 98
rect 410 90 412 98
rect 420 90 422 98
rect 440 90 442 98
rect 450 90 452 98
rect 470 90 472 98
rect 480 90 482 98
rect 500 90 502 98
rect 510 90 512 98
rect 530 90 532 98
rect 540 90 542 98
rect 560 90 562 98
rect 30 88 62 90
rect 70 88 92 90
rect 100 88 122 90
rect 130 88 152 90
rect 160 88 182 90
rect 190 88 212 90
rect 220 88 242 90
rect 250 88 272 90
rect 280 88 302 90
rect 310 88 332 90
rect 340 88 362 90
rect 370 88 392 90
rect 400 88 422 90
rect 430 88 452 90
rect 460 88 482 90
rect 490 88 512 90
rect 520 88 542 90
rect 550 88 570 90
rect 30 80 32 88
rect 40 80 42 88
rect 50 80 52 88
rect 70 80 72 88
rect 80 80 82 88
rect 100 80 102 88
rect 110 80 112 88
rect 130 80 132 88
rect 140 80 142 88
rect 160 80 162 88
rect 170 80 172 88
rect 190 80 192 88
rect 200 80 202 88
rect 220 80 222 88
rect 230 80 232 88
rect 250 80 252 88
rect 260 80 262 88
rect 280 80 282 88
rect 290 80 292 88
rect 310 80 312 88
rect 320 80 322 88
rect 340 80 342 88
rect 350 80 352 88
rect 370 80 372 88
rect 380 80 382 88
rect 400 80 402 88
rect 410 80 412 88
rect 430 80 432 88
rect 440 80 442 88
rect 460 80 462 88
rect 470 80 472 88
rect 490 80 492 88
rect 500 80 502 88
rect 520 80 522 88
rect 530 80 532 88
rect 550 80 552 88
rect 560 80 562 88
rect 30 78 62 80
rect 70 78 92 80
rect 100 78 122 80
rect 130 78 152 80
rect 160 78 182 80
rect 190 78 212 80
rect 220 78 242 80
rect 250 78 272 80
rect 280 78 302 80
rect 310 78 332 80
rect 340 78 362 80
rect 370 78 392 80
rect 400 78 422 80
rect 430 78 452 80
rect 460 78 482 80
rect 490 78 512 80
rect 520 78 542 80
rect 550 78 570 80
rect 30 70 32 78
rect 40 70 42 78
rect 50 70 52 78
rect 60 70 62 78
rect 80 70 82 78
rect 90 70 92 78
rect 110 70 112 78
rect 120 70 122 78
rect 140 70 142 78
rect 150 70 152 78
rect 170 70 172 78
rect 180 70 182 78
rect 200 70 202 78
rect 210 70 212 78
rect 230 70 232 78
rect 240 70 242 78
rect 260 70 262 78
rect 270 70 272 78
rect 290 70 292 78
rect 300 70 302 78
rect 320 70 322 78
rect 330 70 332 78
rect 350 70 352 78
rect 360 70 362 78
rect 380 70 382 78
rect 390 70 392 78
rect 410 70 412 78
rect 420 70 422 78
rect 440 70 442 78
rect 450 70 452 78
rect 470 70 472 78
rect 480 70 482 78
rect 500 70 502 78
rect 510 70 512 78
rect 530 70 532 78
rect 540 70 542 78
rect 560 70 562 78
rect 30 68 62 70
rect 70 68 92 70
rect 100 68 122 70
rect 130 68 152 70
rect 160 68 182 70
rect 190 68 212 70
rect 220 68 242 70
rect 250 68 272 70
rect 280 68 302 70
rect 310 68 332 70
rect 340 68 362 70
rect 370 68 392 70
rect 400 68 422 70
rect 430 68 452 70
rect 460 68 482 70
rect 490 68 512 70
rect 520 68 542 70
rect 550 68 570 70
rect 30 60 32 68
rect 40 60 42 68
rect 50 60 52 68
rect 70 60 72 68
rect 80 60 82 68
rect 100 60 102 68
rect 110 60 112 68
rect 130 60 132 68
rect 140 60 142 68
rect 160 60 162 68
rect 170 60 172 68
rect 190 60 192 68
rect 200 60 202 68
rect 220 60 222 68
rect 230 60 232 68
rect 250 60 252 68
rect 260 60 262 68
rect 280 60 282 68
rect 290 60 292 68
rect 310 60 312 68
rect 320 60 322 68
rect 340 60 342 68
rect 350 60 352 68
rect 370 60 372 68
rect 380 60 382 68
rect 400 60 402 68
rect 410 60 412 68
rect 430 60 432 68
rect 440 60 442 68
rect 460 60 462 68
rect 470 60 472 68
rect 490 60 492 68
rect 500 60 502 68
rect 520 60 522 68
rect 530 60 532 68
rect 550 60 552 68
rect 560 60 562 68
rect 30 58 62 60
rect 70 58 92 60
rect 100 58 122 60
rect 130 58 152 60
rect 160 58 182 60
rect 190 58 212 60
rect 220 58 242 60
rect 250 58 272 60
rect 280 58 302 60
rect 310 58 332 60
rect 340 58 362 60
rect 370 58 392 60
rect 400 58 422 60
rect 430 58 452 60
rect 460 58 482 60
rect 490 58 512 60
rect 520 58 542 60
rect 550 58 570 60
rect 30 50 32 58
rect 40 50 42 58
rect 50 50 52 58
rect 60 50 62 58
rect 80 50 82 58
rect 90 50 92 58
rect 110 50 112 58
rect 120 50 122 58
rect 140 50 142 58
rect 150 50 152 58
rect 170 50 172 58
rect 180 50 182 58
rect 200 50 202 58
rect 210 50 212 58
rect 230 50 232 58
rect 240 50 242 58
rect 260 50 262 58
rect 270 50 272 58
rect 290 50 292 58
rect 300 50 302 58
rect 320 50 322 58
rect 330 50 332 58
rect 350 50 352 58
rect 360 50 362 58
rect 380 50 382 58
rect 390 50 392 58
rect 410 50 412 58
rect 420 50 422 58
rect 440 50 442 58
rect 450 50 452 58
rect 470 50 472 58
rect 480 50 482 58
rect 500 50 502 58
rect 510 50 512 58
rect 530 50 532 58
rect 540 50 542 58
rect 560 50 562 58
rect 30 48 62 50
rect 70 48 92 50
rect 100 48 122 50
rect 130 48 152 50
rect 160 48 182 50
rect 190 48 212 50
rect 220 48 242 50
rect 250 48 272 50
rect 280 48 302 50
rect 310 48 332 50
rect 340 48 362 50
rect 370 48 392 50
rect 400 48 422 50
rect 430 48 452 50
rect 460 48 482 50
rect 490 48 512 50
rect 520 48 542 50
rect 550 48 570 50
rect 30 40 32 48
rect 40 40 42 48
rect 50 40 52 48
rect 70 40 72 48
rect 80 40 82 48
rect 100 40 102 48
rect 110 40 112 48
rect 130 40 132 48
rect 140 40 142 48
rect 160 40 162 48
rect 170 40 172 48
rect 190 40 192 48
rect 200 40 202 48
rect 220 40 222 48
rect 230 40 232 48
rect 250 40 252 48
rect 260 40 262 48
rect 280 40 282 48
rect 290 40 292 48
rect 310 40 312 48
rect 320 40 322 48
rect 340 40 342 48
rect 350 40 352 48
rect 370 40 372 48
rect 380 40 382 48
rect 400 40 402 48
rect 410 40 412 48
rect 430 40 432 48
rect 440 40 442 48
rect 460 40 462 48
rect 470 40 472 48
rect 490 40 492 48
rect 500 40 502 48
rect 520 40 522 48
rect 530 40 532 48
rect 550 40 552 48
rect 560 40 562 48
rect 30 38 62 40
rect 70 38 92 40
rect 100 38 122 40
rect 130 38 152 40
rect 160 38 182 40
rect 190 38 212 40
rect 220 38 242 40
rect 250 38 272 40
rect 280 38 302 40
rect 310 38 332 40
rect 340 38 362 40
rect 370 38 392 40
rect 400 38 422 40
rect 430 38 452 40
rect 460 38 482 40
rect 490 38 512 40
rect 520 38 542 40
rect 550 38 570 40
rect 30 30 32 38
rect 40 30 42 38
rect 50 30 52 38
rect 60 30 62 38
rect 80 30 82 38
rect 90 30 92 38
rect 110 30 112 38
rect 120 30 122 38
rect 140 30 142 38
rect 150 30 152 38
rect 170 30 172 38
rect 180 30 182 38
rect 200 30 202 38
rect 210 30 212 38
rect 230 30 232 38
rect 240 30 242 38
rect 260 30 262 38
rect 270 30 272 38
rect 290 30 292 38
rect 300 30 302 38
rect 320 30 322 38
rect 330 30 332 38
rect 350 30 352 38
rect 360 30 362 38
rect 380 30 382 38
rect 390 30 392 38
rect 410 30 412 38
rect 420 30 422 38
rect 440 30 442 38
rect 450 30 452 38
rect 470 30 472 38
rect 480 30 482 38
rect 500 30 502 38
rect 510 30 512 38
rect 530 30 532 38
rect 540 30 542 38
rect 560 30 562 38
rect 586 14 588 506
rect 12 12 588 14
rect 12 4 16 12
rect 584 4 588 12
rect 596 4 600 512
rect 0 2 600 4
<< m2contact >>
rect 56 1290 64 1298
rect 86 1290 94 1298
rect 116 1290 124 1298
rect 146 1290 154 1298
rect 176 1290 184 1298
rect 206 1290 214 1298
rect 236 1290 244 1298
rect 266 1290 274 1298
rect 296 1290 304 1298
rect 326 1290 334 1298
rect 356 1290 364 1298
rect 386 1290 394 1298
rect 416 1290 424 1298
rect 446 1290 454 1298
rect 476 1290 484 1298
rect 506 1290 514 1298
rect 536 1290 544 1298
rect 46 1280 54 1288
rect 66 1280 74 1288
rect 96 1280 104 1288
rect 126 1280 134 1288
rect 156 1280 164 1288
rect 186 1280 194 1288
rect 216 1280 224 1288
rect 246 1280 254 1288
rect 276 1280 284 1288
rect 306 1280 314 1288
rect 336 1280 344 1288
rect 366 1280 374 1288
rect 396 1280 404 1288
rect 426 1280 434 1288
rect 456 1280 464 1288
rect 486 1280 494 1288
rect 516 1280 524 1288
rect 546 1280 554 1288
rect 56 1270 64 1278
rect 86 1270 94 1278
rect 116 1270 124 1278
rect 146 1270 154 1278
rect 176 1270 184 1278
rect 206 1270 214 1278
rect 236 1270 244 1278
rect 266 1270 274 1278
rect 296 1270 304 1278
rect 326 1270 334 1278
rect 356 1270 364 1278
rect 386 1270 394 1278
rect 416 1270 424 1278
rect 446 1270 454 1278
rect 476 1270 484 1278
rect 506 1270 514 1278
rect 536 1270 544 1278
rect 46 1260 54 1268
rect 66 1260 74 1268
rect 96 1260 104 1268
rect 126 1260 134 1268
rect 156 1260 164 1268
rect 186 1260 194 1268
rect 216 1260 224 1268
rect 246 1260 254 1268
rect 276 1260 284 1268
rect 306 1260 314 1268
rect 336 1260 344 1268
rect 366 1260 374 1268
rect 396 1260 404 1268
rect 426 1260 434 1268
rect 456 1260 464 1268
rect 486 1260 494 1268
rect 516 1260 524 1268
rect 546 1260 554 1268
rect 56 1250 64 1258
rect 86 1250 94 1258
rect 116 1250 124 1258
rect 146 1250 154 1258
rect 176 1250 184 1258
rect 206 1250 214 1258
rect 236 1250 244 1258
rect 266 1250 274 1258
rect 296 1250 304 1258
rect 326 1250 334 1258
rect 356 1250 364 1258
rect 386 1250 394 1258
rect 416 1250 424 1258
rect 446 1250 454 1258
rect 476 1250 484 1258
rect 506 1250 514 1258
rect 536 1250 544 1258
rect 46 1240 54 1248
rect 66 1240 74 1248
rect 96 1240 104 1248
rect 126 1240 134 1248
rect 156 1240 164 1248
rect 186 1240 194 1248
rect 216 1240 224 1248
rect 246 1240 254 1248
rect 276 1240 284 1248
rect 306 1240 314 1248
rect 336 1240 344 1248
rect 366 1240 374 1248
rect 396 1240 404 1248
rect 426 1240 434 1248
rect 456 1240 464 1248
rect 486 1240 494 1248
rect 516 1240 524 1248
rect 546 1240 554 1248
rect 56 1230 64 1238
rect 86 1230 94 1238
rect 116 1230 124 1238
rect 146 1230 154 1238
rect 176 1230 184 1238
rect 206 1230 214 1238
rect 236 1230 244 1238
rect 266 1230 274 1238
rect 296 1230 304 1238
rect 326 1230 334 1238
rect 356 1230 364 1238
rect 386 1230 394 1238
rect 416 1230 424 1238
rect 446 1230 454 1238
rect 476 1230 484 1238
rect 506 1230 514 1238
rect 536 1230 544 1238
rect 46 1220 54 1228
rect 66 1220 74 1228
rect 96 1220 104 1228
rect 126 1220 134 1228
rect 156 1220 164 1228
rect 186 1220 194 1228
rect 216 1220 224 1228
rect 246 1220 254 1228
rect 276 1220 284 1228
rect 306 1220 314 1228
rect 336 1220 344 1228
rect 366 1220 374 1228
rect 396 1220 404 1228
rect 426 1220 434 1228
rect 456 1220 464 1228
rect 486 1220 494 1228
rect 516 1220 524 1228
rect 546 1220 554 1228
rect 56 1210 64 1218
rect 86 1210 94 1218
rect 116 1210 124 1218
rect 146 1210 154 1218
rect 176 1210 184 1218
rect 206 1210 214 1218
rect 236 1210 244 1218
rect 266 1210 274 1218
rect 296 1210 304 1218
rect 326 1210 334 1218
rect 356 1210 364 1218
rect 386 1210 394 1218
rect 416 1210 424 1218
rect 446 1210 454 1218
rect 476 1210 484 1218
rect 506 1210 514 1218
rect 536 1210 544 1218
rect 46 1200 54 1208
rect 66 1200 74 1208
rect 96 1200 104 1208
rect 126 1200 134 1208
rect 156 1200 164 1208
rect 186 1200 194 1208
rect 216 1200 224 1208
rect 246 1200 254 1208
rect 276 1200 284 1208
rect 306 1200 314 1208
rect 336 1200 344 1208
rect 366 1200 374 1208
rect 396 1200 404 1208
rect 426 1200 434 1208
rect 456 1200 464 1208
rect 486 1200 494 1208
rect 516 1200 524 1208
rect 546 1200 554 1208
rect 56 1190 64 1198
rect 86 1190 94 1198
rect 116 1190 124 1198
rect 146 1190 154 1198
rect 176 1190 184 1198
rect 206 1190 214 1198
rect 236 1190 244 1198
rect 266 1190 274 1198
rect 296 1190 304 1198
rect 326 1190 334 1198
rect 356 1190 364 1198
rect 386 1190 394 1198
rect 416 1190 424 1198
rect 446 1190 454 1198
rect 476 1190 484 1198
rect 506 1190 514 1198
rect 536 1190 544 1198
rect 46 1180 54 1188
rect 66 1180 74 1188
rect 516 1180 524 1188
rect 546 1180 554 1188
rect 56 1170 64 1178
rect 86 1170 94 1178
rect 116 1170 124 1178
rect 146 1170 154 1178
rect 176 1170 184 1178
rect 206 1170 214 1178
rect 236 1170 244 1178
rect 266 1170 274 1178
rect 296 1170 304 1178
rect 326 1170 334 1178
rect 356 1170 364 1178
rect 386 1170 394 1178
rect 416 1170 424 1178
rect 446 1170 454 1178
rect 476 1170 484 1178
rect 506 1170 514 1178
rect 536 1170 544 1178
rect 46 1160 54 1168
rect 66 1160 74 1168
rect 96 1160 104 1168
rect 126 1160 134 1168
rect 156 1160 164 1168
rect 186 1160 194 1168
rect 216 1160 224 1168
rect 246 1160 254 1168
rect 276 1160 284 1168
rect 306 1160 314 1168
rect 336 1160 344 1168
rect 366 1160 374 1168
rect 396 1160 404 1168
rect 426 1160 434 1168
rect 456 1160 464 1168
rect 486 1160 494 1168
rect 516 1160 524 1168
rect 546 1160 554 1168
rect 56 1150 64 1158
rect 86 1150 94 1158
rect 116 1150 124 1158
rect 146 1150 154 1158
rect 176 1150 184 1158
rect 206 1150 214 1158
rect 236 1150 244 1158
rect 266 1150 274 1158
rect 296 1150 304 1158
rect 326 1150 334 1158
rect 356 1150 364 1158
rect 386 1150 394 1158
rect 416 1150 424 1158
rect 446 1150 454 1158
rect 476 1150 484 1158
rect 506 1150 514 1158
rect 536 1150 544 1158
rect 46 1140 54 1148
rect 66 1140 74 1148
rect 96 1140 104 1148
rect 126 1140 134 1148
rect 156 1140 164 1148
rect 186 1140 194 1148
rect 216 1140 224 1148
rect 246 1140 254 1148
rect 276 1140 284 1148
rect 306 1140 314 1148
rect 336 1140 344 1148
rect 366 1140 374 1148
rect 396 1140 404 1148
rect 426 1140 434 1148
rect 456 1140 464 1148
rect 486 1140 494 1148
rect 516 1140 524 1148
rect 546 1140 554 1148
rect 56 1130 64 1138
rect 86 1130 94 1138
rect 116 1130 124 1138
rect 146 1130 154 1138
rect 176 1130 184 1138
rect 206 1130 214 1138
rect 236 1130 244 1138
rect 266 1130 274 1138
rect 296 1130 304 1138
rect 326 1130 334 1138
rect 356 1130 364 1138
rect 386 1130 394 1138
rect 416 1130 424 1138
rect 446 1130 454 1138
rect 476 1130 484 1138
rect 506 1130 514 1138
rect 536 1130 544 1138
rect 46 1120 54 1128
rect 66 1120 74 1128
rect 96 1120 104 1128
rect 126 1120 134 1128
rect 156 1120 164 1128
rect 186 1120 194 1128
rect 216 1120 224 1128
rect 246 1120 254 1128
rect 276 1120 284 1128
rect 306 1120 314 1128
rect 336 1120 344 1128
rect 366 1120 374 1128
rect 396 1120 404 1128
rect 426 1120 434 1128
rect 456 1120 464 1128
rect 486 1120 494 1128
rect 56 1110 64 1118
rect 76 1110 84 1118
rect 46 1100 54 1108
rect 66 1100 74 1108
rect 96 1100 104 1108
rect 126 1100 134 1108
rect 156 1100 164 1108
rect 186 1100 194 1108
rect 216 1100 224 1108
rect 246 1100 254 1108
rect 276 1100 284 1108
rect 306 1100 314 1108
rect 336 1100 344 1108
rect 366 1100 374 1108
rect 396 1100 404 1108
rect 426 1100 434 1108
rect 456 1100 464 1108
rect 486 1100 494 1108
rect 516 1100 524 1128
rect 546 1120 554 1128
rect 536 1110 544 1118
rect 546 1100 554 1108
rect 56 1090 64 1098
rect 86 1090 94 1098
rect 116 1090 124 1098
rect 146 1090 154 1098
rect 176 1090 184 1098
rect 206 1090 214 1098
rect 236 1090 244 1098
rect 266 1090 274 1098
rect 296 1090 304 1098
rect 326 1090 334 1098
rect 356 1090 364 1098
rect 386 1090 394 1098
rect 416 1090 424 1098
rect 446 1090 454 1098
rect 476 1090 484 1098
rect 506 1090 514 1098
rect 536 1090 544 1098
rect 46 1080 54 1088
rect 66 1080 74 1088
rect 96 1080 104 1088
rect 126 1080 134 1088
rect 156 1080 164 1088
rect 186 1080 194 1088
rect 216 1080 224 1088
rect 246 1080 254 1088
rect 276 1080 284 1088
rect 306 1080 314 1088
rect 336 1080 344 1088
rect 366 1080 374 1088
rect 396 1080 404 1088
rect 426 1080 434 1088
rect 456 1080 464 1088
rect 486 1080 494 1088
rect 516 1080 524 1088
rect 546 1080 554 1088
rect 56 1070 64 1078
rect 86 1070 94 1078
rect 116 1070 124 1078
rect 146 1070 154 1078
rect 176 1070 184 1078
rect 206 1070 214 1078
rect 236 1070 244 1078
rect 266 1070 274 1078
rect 296 1070 304 1078
rect 326 1070 334 1078
rect 356 1070 364 1078
rect 386 1070 394 1078
rect 416 1070 424 1078
rect 446 1070 454 1078
rect 476 1070 484 1078
rect 506 1070 514 1078
rect 536 1070 544 1078
rect 46 1060 54 1068
rect 66 1060 74 1068
rect 96 1060 104 1068
rect 126 1060 134 1068
rect 156 1060 164 1068
rect 186 1060 194 1068
rect 216 1060 224 1068
rect 246 1060 254 1068
rect 276 1060 284 1068
rect 306 1060 314 1068
rect 336 1060 344 1068
rect 366 1060 374 1068
rect 396 1060 404 1068
rect 426 1060 434 1068
rect 456 1060 464 1068
rect 486 1060 494 1068
rect 516 1060 524 1068
rect 546 1060 554 1068
rect 56 1050 64 1058
rect 86 1050 94 1058
rect 116 1050 124 1058
rect 146 1050 154 1058
rect 176 1050 184 1058
rect 206 1050 214 1058
rect 236 1050 244 1058
rect 266 1050 274 1058
rect 296 1050 304 1058
rect 326 1050 334 1058
rect 356 1050 364 1058
rect 386 1050 394 1058
rect 416 1050 424 1058
rect 446 1050 454 1058
rect 476 1050 484 1058
rect 506 1050 514 1058
rect 536 1050 544 1058
rect 46 1040 54 1048
rect 66 1040 74 1048
rect 96 1040 104 1048
rect 126 1040 134 1048
rect 156 1040 164 1048
rect 186 1040 194 1048
rect 216 1040 224 1048
rect 246 1040 254 1048
rect 276 1040 284 1048
rect 306 1040 314 1048
rect 336 1040 344 1048
rect 366 1040 374 1048
rect 396 1040 404 1048
rect 426 1040 434 1048
rect 456 1040 464 1048
rect 486 1040 494 1048
rect 56 1030 64 1038
rect 86 1030 94 1038
rect 46 1020 54 1028
rect 66 1020 74 1028
rect 96 1020 104 1028
rect 126 1020 134 1028
rect 156 1020 164 1028
rect 186 1020 194 1028
rect 216 1020 224 1028
rect 246 1020 254 1028
rect 276 1020 284 1028
rect 306 1020 314 1028
rect 336 1020 344 1028
rect 366 1020 374 1028
rect 396 1020 404 1028
rect 426 1020 434 1028
rect 456 1020 464 1028
rect 486 1020 494 1028
rect 516 1020 524 1048
rect 546 1040 554 1048
rect 536 1030 544 1038
rect 546 1020 554 1028
rect 56 1010 64 1018
rect 86 1010 94 1018
rect 116 1010 124 1018
rect 146 1010 154 1018
rect 176 1010 184 1018
rect 206 1010 214 1018
rect 236 1010 244 1018
rect 266 1010 274 1018
rect 296 1010 304 1018
rect 326 1010 334 1018
rect 356 1010 364 1018
rect 386 1010 394 1018
rect 416 1010 424 1018
rect 446 1010 454 1018
rect 476 1010 484 1018
rect 506 1010 514 1018
rect 536 1010 544 1018
rect 46 1000 54 1008
rect 66 1000 74 1008
rect 96 1000 104 1008
rect 126 1000 134 1008
rect 156 1000 164 1008
rect 186 1000 194 1008
rect 216 1000 224 1008
rect 246 1000 254 1008
rect 276 1000 284 1008
rect 306 1000 314 1008
rect 336 1000 344 1008
rect 366 1000 374 1008
rect 396 1000 404 1008
rect 426 1000 434 1008
rect 456 1000 464 1008
rect 486 1000 494 1008
rect 516 1000 524 1008
rect 546 1000 554 1008
rect 56 990 64 998
rect 86 990 94 998
rect 116 990 124 998
rect 146 990 154 998
rect 176 990 184 998
rect 206 990 214 998
rect 236 990 244 998
rect 266 990 274 998
rect 296 990 304 998
rect 326 990 334 998
rect 356 990 364 998
rect 386 990 394 998
rect 416 990 424 998
rect 446 990 454 998
rect 476 990 484 998
rect 506 990 514 998
rect 536 990 544 998
rect 46 980 54 988
rect 66 980 74 988
rect 96 980 104 988
rect 126 980 134 988
rect 156 980 164 988
rect 186 980 194 988
rect 216 980 224 988
rect 246 980 254 988
rect 276 980 284 988
rect 306 980 314 988
rect 336 980 344 988
rect 366 980 374 988
rect 396 980 404 988
rect 426 980 434 988
rect 456 980 464 988
rect 486 980 494 988
rect 516 980 524 988
rect 546 980 554 988
rect 56 970 64 978
rect 86 970 94 978
rect 116 970 124 978
rect 146 970 154 978
rect 176 970 184 978
rect 206 970 214 978
rect 236 970 244 978
rect 266 970 274 978
rect 296 970 304 978
rect 326 970 334 978
rect 356 970 364 978
rect 386 970 394 978
rect 416 970 424 978
rect 446 970 454 978
rect 476 970 484 978
rect 506 970 514 978
rect 536 970 544 978
rect 46 960 54 968
rect 546 960 554 968
rect 56 950 64 958
rect 86 950 94 958
rect 116 950 124 958
rect 146 950 154 958
rect 176 950 184 958
rect 206 950 214 958
rect 236 950 244 958
rect 266 950 274 958
rect 296 950 304 958
rect 326 950 334 958
rect 356 950 364 958
rect 386 950 394 958
rect 416 950 424 958
rect 446 950 454 958
rect 476 950 484 958
rect 506 950 514 958
rect 536 950 544 958
rect 46 940 54 948
rect 66 940 74 948
rect 96 940 104 948
rect 126 940 134 948
rect 156 940 164 948
rect 186 940 194 948
rect 216 940 224 948
rect 246 940 254 948
rect 276 940 284 948
rect 306 940 314 948
rect 336 940 344 948
rect 366 940 374 948
rect 396 940 404 948
rect 426 940 434 948
rect 456 940 464 948
rect 486 940 494 948
rect 516 940 524 948
rect 546 940 554 948
rect 56 930 64 938
rect 86 930 94 938
rect 116 930 124 938
rect 146 930 154 938
rect 176 930 184 938
rect 206 930 214 938
rect 236 930 244 938
rect 266 930 274 938
rect 296 930 304 938
rect 326 930 334 938
rect 356 930 364 938
rect 386 930 394 938
rect 416 930 424 938
rect 446 930 454 938
rect 476 930 484 938
rect 506 930 514 938
rect 536 930 544 938
rect 46 920 54 928
rect 66 920 74 928
rect 96 920 104 928
rect 126 920 134 928
rect 156 920 164 928
rect 186 920 194 928
rect 216 920 224 928
rect 246 920 254 928
rect 276 920 284 928
rect 306 920 314 928
rect 336 920 344 928
rect 366 920 374 928
rect 396 920 404 928
rect 426 920 434 928
rect 456 920 464 928
rect 486 920 494 928
rect 516 920 524 928
rect 546 920 554 928
rect 56 910 64 918
rect 86 910 94 918
rect 116 910 124 918
rect 146 910 154 918
rect 176 910 184 918
rect 206 910 214 918
rect 236 910 244 918
rect 266 910 274 918
rect 296 910 304 918
rect 326 910 334 918
rect 356 910 364 918
rect 386 910 394 918
rect 416 910 424 918
rect 446 910 454 918
rect 476 910 484 918
rect 506 910 514 918
rect 536 910 544 918
rect 46 900 54 908
rect 66 900 74 908
rect 96 900 104 908
rect 126 900 134 908
rect 156 900 164 908
rect 186 900 194 908
rect 216 900 224 908
rect 246 900 254 908
rect 276 900 284 908
rect 306 900 314 908
rect 336 900 344 908
rect 366 900 374 908
rect 396 900 404 908
rect 426 900 434 908
rect 456 900 464 908
rect 486 900 494 908
rect 516 900 524 908
rect 546 900 554 908
rect 56 890 64 898
rect 86 890 94 898
rect 116 890 124 898
rect 146 890 154 898
rect 176 890 184 898
rect 206 890 214 898
rect 236 890 244 898
rect 266 890 274 898
rect 296 890 304 898
rect 326 890 334 898
rect 356 890 364 898
rect 386 890 394 898
rect 416 890 424 898
rect 446 890 454 898
rect 476 890 484 898
rect 506 890 514 898
rect 536 890 544 898
rect 46 880 54 888
rect 66 880 74 888
rect 96 880 104 888
rect 126 880 134 888
rect 156 880 164 888
rect 186 880 194 888
rect 216 880 224 888
rect 246 880 254 888
rect 276 880 284 888
rect 306 880 314 888
rect 336 880 344 888
rect 366 880 374 888
rect 396 880 404 888
rect 426 880 434 888
rect 456 880 464 888
rect 486 880 494 888
rect 516 880 524 888
rect 546 880 554 888
rect 14 828 22 836
rect 44 828 52 836
rect 74 828 82 836
rect 104 828 112 836
rect 134 828 142 836
rect 164 828 172 836
rect 194 828 202 836
rect 224 828 232 836
rect 244 828 252 836
rect 266 828 274 836
rect 296 828 304 836
rect 326 828 334 836
rect 348 828 356 836
rect 368 828 376 836
rect 398 828 406 836
rect 428 828 436 836
rect 458 828 466 836
rect 488 828 496 836
rect 518 828 526 836
rect 548 828 556 836
rect 578 828 586 836
rect 4 818 12 826
rect 24 818 32 826
rect 54 818 62 826
rect 84 818 92 826
rect 114 818 122 826
rect 144 818 152 826
rect 174 818 182 826
rect 204 818 212 826
rect 234 818 242 826
rect 256 818 264 826
rect 276 818 284 826
rect 306 818 314 826
rect 336 818 344 826
rect 358 818 366 826
rect 388 818 396 826
rect 418 818 426 826
rect 448 818 456 826
rect 478 818 486 826
rect 508 818 516 826
rect 538 818 546 826
rect 568 818 576 826
rect 588 818 596 826
rect 14 808 22 816
rect 44 808 52 816
rect 74 808 82 816
rect 104 808 112 816
rect 134 808 142 816
rect 164 808 172 816
rect 194 808 202 816
rect 224 808 232 816
rect 244 808 252 816
rect 266 808 274 816
rect 296 808 304 816
rect 326 808 334 816
rect 348 808 356 816
rect 368 808 376 816
rect 398 808 406 816
rect 428 808 436 816
rect 458 808 466 816
rect 488 808 496 816
rect 518 808 526 816
rect 548 808 556 816
rect 578 808 586 816
rect 4 798 12 806
rect 24 798 32 806
rect 54 798 62 806
rect 84 798 92 806
rect 114 798 122 806
rect 144 798 152 806
rect 174 798 182 806
rect 204 798 212 806
rect 234 798 242 806
rect 256 798 264 806
rect 276 798 284 806
rect 306 798 314 806
rect 336 798 344 806
rect 358 798 366 806
rect 388 798 396 806
rect 418 798 426 806
rect 448 798 456 806
rect 478 798 486 806
rect 508 798 516 806
rect 538 798 546 806
rect 568 798 576 806
rect 588 798 596 806
rect 14 788 22 796
rect 44 788 52 796
rect 74 788 82 796
rect 104 788 112 796
rect 134 788 142 796
rect 164 788 172 796
rect 194 788 202 796
rect 224 788 232 796
rect 244 788 252 796
rect 266 788 274 796
rect 296 788 304 796
rect 326 788 334 796
rect 348 788 356 796
rect 368 788 376 796
rect 398 788 406 796
rect 428 788 436 796
rect 458 788 466 796
rect 488 788 496 796
rect 518 788 526 796
rect 548 788 556 796
rect 578 788 586 796
rect 4 778 12 786
rect 24 778 32 786
rect 54 778 62 786
rect 84 778 92 786
rect 114 778 122 786
rect 144 778 152 786
rect 174 778 182 786
rect 204 778 212 786
rect 234 778 242 786
rect 256 778 264 786
rect 276 778 284 786
rect 306 778 314 786
rect 336 778 344 786
rect 358 778 366 786
rect 388 778 396 786
rect 418 778 426 786
rect 448 778 456 786
rect 478 778 486 786
rect 508 778 516 786
rect 538 778 546 786
rect 568 778 576 786
rect 588 778 596 786
rect 14 768 22 776
rect 44 768 52 776
rect 74 768 82 776
rect 518 768 526 776
rect 548 768 556 776
rect 578 768 586 776
rect 4 758 12 766
rect 24 758 32 766
rect 54 758 62 766
rect 84 758 92 766
rect 114 758 122 766
rect 144 758 152 766
rect 174 758 182 766
rect 204 758 212 766
rect 234 758 242 766
rect 256 758 264 766
rect 276 758 284 766
rect 306 758 314 766
rect 336 758 344 766
rect 358 758 366 766
rect 388 758 396 766
rect 418 758 426 766
rect 448 758 456 766
rect 478 758 486 766
rect 508 758 516 766
rect 538 758 546 766
rect 568 758 576 766
rect 588 758 596 766
rect 14 748 22 756
rect 44 748 52 756
rect 74 748 82 756
rect 104 748 112 756
rect 134 748 142 756
rect 164 748 172 756
rect 194 748 202 756
rect 224 748 232 756
rect 244 748 252 756
rect 266 748 274 756
rect 296 748 304 756
rect 326 748 334 756
rect 348 748 356 756
rect 368 748 376 756
rect 398 748 406 756
rect 428 748 436 756
rect 458 748 466 756
rect 488 748 496 756
rect 518 748 526 756
rect 548 748 556 756
rect 578 748 586 756
rect 4 738 12 746
rect 24 738 32 746
rect 54 738 62 746
rect 84 738 92 746
rect 114 738 122 746
rect 144 738 152 746
rect 174 738 182 746
rect 204 738 212 746
rect 234 738 242 746
rect 256 738 264 746
rect 276 738 284 746
rect 306 738 314 746
rect 336 738 344 746
rect 358 738 366 746
rect 388 738 396 746
rect 418 738 426 746
rect 448 738 456 746
rect 478 738 486 746
rect 508 738 516 746
rect 538 738 546 746
rect 568 738 576 746
rect 588 738 596 746
rect 14 728 22 736
rect 224 728 232 736
rect 244 728 252 736
rect 266 728 274 736
rect 296 728 304 736
rect 326 728 334 736
rect 348 728 356 736
rect 368 728 376 736
rect 578 728 586 736
rect 4 718 12 726
rect 24 718 32 726
rect 54 718 62 726
rect 84 718 92 726
rect 114 718 122 726
rect 144 718 152 726
rect 174 718 182 726
rect 204 718 212 726
rect 234 718 242 726
rect 256 718 264 726
rect 276 718 284 726
rect 306 718 314 726
rect 336 718 344 726
rect 358 718 366 726
rect 388 718 396 726
rect 418 718 426 726
rect 448 718 456 726
rect 478 718 486 726
rect 508 718 516 726
rect 538 718 546 726
rect 568 718 576 726
rect 588 718 596 726
rect 14 708 22 716
rect 44 708 52 716
rect 74 708 82 716
rect 104 708 112 716
rect 134 708 142 716
rect 164 708 172 716
rect 194 708 202 716
rect 224 708 232 716
rect 244 708 252 716
rect 266 708 274 716
rect 296 708 304 716
rect 326 708 334 716
rect 348 708 356 716
rect 368 708 376 716
rect 398 708 406 716
rect 428 708 436 716
rect 458 708 466 716
rect 488 708 496 716
rect 518 708 526 716
rect 548 708 556 716
rect 578 708 586 716
rect 4 698 12 706
rect 24 698 32 706
rect 54 698 62 706
rect 84 698 92 706
rect 114 698 122 706
rect 144 698 152 706
rect 174 698 182 706
rect 204 698 212 706
rect 234 698 242 706
rect 256 698 264 706
rect 276 698 284 706
rect 306 698 314 706
rect 336 698 344 706
rect 358 698 366 706
rect 388 698 396 706
rect 418 698 426 706
rect 448 698 456 706
rect 478 698 486 706
rect 508 698 516 706
rect 538 698 546 706
rect 568 698 576 706
rect 588 698 596 706
rect 14 688 22 696
rect 44 688 52 696
rect 74 688 82 696
rect 104 688 112 696
rect 134 688 142 696
rect 164 688 172 696
rect 194 688 202 696
rect 224 688 232 696
rect 244 688 252 696
rect 266 688 274 696
rect 296 688 304 696
rect 326 688 334 696
rect 348 688 356 696
rect 368 688 376 696
rect 398 688 406 696
rect 428 688 436 696
rect 458 688 466 696
rect 488 688 496 696
rect 518 688 526 696
rect 548 688 556 696
rect 578 688 586 696
rect 14 644 22 652
rect 44 644 52 652
rect 74 644 82 652
rect 104 644 112 652
rect 134 644 142 652
rect 164 644 172 652
rect 194 644 202 652
rect 224 644 232 652
rect 244 644 252 652
rect 266 644 274 652
rect 296 644 304 652
rect 326 644 334 652
rect 348 644 356 652
rect 368 644 376 652
rect 398 644 406 652
rect 428 644 436 652
rect 458 644 466 652
rect 488 644 496 652
rect 518 644 526 652
rect 548 644 556 652
rect 578 644 586 652
rect 4 634 12 642
rect 24 634 32 642
rect 54 634 62 642
rect 84 634 92 642
rect 114 634 122 642
rect 144 634 152 642
rect 174 634 182 642
rect 204 634 212 642
rect 234 634 242 642
rect 256 634 264 642
rect 276 634 284 642
rect 306 634 314 642
rect 336 634 344 642
rect 358 634 366 642
rect 388 634 396 642
rect 418 634 426 642
rect 448 634 456 642
rect 478 634 486 642
rect 508 634 516 642
rect 538 634 546 642
rect 568 634 576 642
rect 588 634 596 642
rect 14 624 22 632
rect 44 624 52 632
rect 74 624 82 632
rect 104 624 112 632
rect 134 624 142 632
rect 164 624 172 632
rect 194 624 202 632
rect 224 624 232 632
rect 244 624 252 632
rect 266 624 274 632
rect 296 624 304 632
rect 326 624 334 632
rect 348 624 356 632
rect 368 624 376 632
rect 398 624 406 632
rect 428 624 436 632
rect 458 624 466 632
rect 488 624 496 632
rect 518 624 526 632
rect 548 624 556 632
rect 578 624 586 632
rect 4 614 12 622
rect 24 614 32 622
rect 54 614 62 622
rect 84 614 92 622
rect 114 614 122 622
rect 144 614 152 622
rect 174 614 182 622
rect 204 614 212 622
rect 234 614 242 622
rect 256 614 264 622
rect 276 614 284 622
rect 306 614 314 622
rect 336 614 344 622
rect 358 614 366 622
rect 388 614 396 622
rect 418 614 426 622
rect 448 614 456 622
rect 478 614 486 622
rect 508 614 516 622
rect 538 614 546 622
rect 568 614 576 622
rect 588 614 596 622
rect 14 604 22 612
rect 224 604 232 612
rect 244 604 252 612
rect 266 604 274 612
rect 296 604 304 612
rect 326 604 334 612
rect 348 604 356 612
rect 368 604 376 612
rect 578 604 586 612
rect 4 594 12 602
rect 24 594 32 602
rect 54 594 62 602
rect 84 594 92 602
rect 114 594 122 602
rect 144 594 152 602
rect 174 594 182 602
rect 204 594 212 602
rect 234 594 242 602
rect 256 594 264 602
rect 276 594 284 602
rect 306 594 314 602
rect 336 594 344 602
rect 358 594 366 602
rect 388 594 396 602
rect 418 594 426 602
rect 448 594 456 602
rect 478 594 486 602
rect 508 594 516 602
rect 538 594 546 602
rect 568 594 576 602
rect 588 594 596 602
rect 14 584 22 592
rect 44 584 52 592
rect 74 584 82 592
rect 104 584 112 592
rect 134 584 142 592
rect 164 584 172 592
rect 194 584 202 592
rect 224 584 232 592
rect 244 584 252 592
rect 4 574 12 582
rect 24 574 32 582
rect 54 574 62 582
rect 84 574 92 582
rect 348 584 356 592
rect 368 584 376 592
rect 398 584 406 592
rect 428 584 436 592
rect 458 584 466 592
rect 488 584 496 592
rect 518 584 526 592
rect 548 584 556 592
rect 578 584 586 592
rect 508 574 516 582
rect 538 574 546 582
rect 568 574 576 582
rect 588 574 596 582
rect 14 564 22 572
rect 44 564 52 572
rect 74 564 82 572
rect 104 564 112 572
rect 134 564 142 572
rect 164 564 172 572
rect 194 564 202 572
rect 224 564 232 572
rect 244 564 252 572
rect 266 564 274 572
rect 296 564 304 572
rect 326 564 334 572
rect 348 564 356 572
rect 368 564 376 572
rect 398 564 406 572
rect 428 564 436 572
rect 458 564 466 572
rect 488 564 496 572
rect 518 564 526 572
rect 548 564 556 572
rect 578 564 586 572
rect 4 554 12 562
rect 24 554 32 562
rect 54 554 62 562
rect 84 554 92 562
rect 114 554 122 562
rect 144 554 152 562
rect 174 554 182 562
rect 204 554 212 562
rect 234 554 242 562
rect 256 554 264 562
rect 276 554 284 562
rect 306 554 314 562
rect 336 554 344 562
rect 358 554 366 562
rect 388 554 396 562
rect 418 554 426 562
rect 448 554 456 562
rect 478 554 486 562
rect 508 554 516 562
rect 538 554 546 562
rect 568 554 576 562
rect 588 554 596 562
rect 14 544 22 552
rect 44 544 52 552
rect 74 544 82 552
rect 104 544 112 552
rect 134 544 142 552
rect 164 544 172 552
rect 194 544 202 552
rect 224 544 232 552
rect 244 544 252 552
rect 266 544 274 552
rect 296 544 304 552
rect 326 544 334 552
rect 348 544 356 552
rect 368 544 376 552
rect 398 544 406 552
rect 428 544 436 552
rect 458 544 466 552
rect 488 544 496 552
rect 518 544 526 552
rect 548 544 556 552
rect 578 544 586 552
rect 4 534 12 542
rect 24 534 32 542
rect 54 534 62 542
rect 84 534 92 542
rect 114 534 122 542
rect 144 534 152 542
rect 174 534 182 542
rect 204 534 212 542
rect 234 534 242 542
rect 256 534 264 542
rect 276 534 284 542
rect 306 534 314 542
rect 336 534 344 542
rect 358 534 366 542
rect 388 534 396 542
rect 418 534 426 542
rect 448 534 456 542
rect 478 534 486 542
rect 508 534 516 542
rect 538 534 546 542
rect 568 534 576 542
rect 588 534 596 542
rect 14 524 22 532
rect 44 524 52 532
rect 74 524 82 532
rect 104 524 112 532
rect 134 524 142 532
rect 164 524 172 532
rect 194 524 202 532
rect 224 524 232 532
rect 244 524 252 532
rect 266 524 274 532
rect 296 524 304 532
rect 326 524 334 532
rect 348 524 356 532
rect 368 524 376 532
rect 398 524 406 532
rect 428 524 436 532
rect 458 524 466 532
rect 488 524 496 532
rect 518 524 526 532
rect 548 524 556 532
rect 578 524 586 532
rect 14 508 22 516
rect 34 508 42 516
rect 54 508 62 516
rect 74 508 82 516
rect 94 508 102 516
rect 114 508 122 516
rect 134 508 142 516
rect 154 508 162 516
rect 174 508 182 516
rect 194 508 202 516
rect 214 508 222 516
rect 234 508 242 516
rect 254 508 262 516
rect 274 508 282 516
rect 294 508 302 516
rect 308 508 316 516
rect 328 508 336 516
rect 348 508 356 516
rect 368 508 376 516
rect 388 508 396 516
rect 408 508 416 516
rect 428 508 436 516
rect 448 508 456 516
rect 468 508 476 516
rect 488 508 496 516
rect 508 508 516 516
rect 528 508 536 516
rect 548 508 556 516
rect 568 508 576 516
rect 32 450 40 458
rect 52 450 60 458
rect 82 450 90 458
rect 112 450 120 458
rect 142 450 150 458
rect 172 450 180 458
rect 202 450 210 458
rect 232 450 240 458
rect 262 450 270 458
rect 292 450 300 458
rect 322 450 330 458
rect 352 450 360 458
rect 382 450 390 458
rect 412 450 420 458
rect 442 450 450 458
rect 472 450 480 458
rect 502 450 510 458
rect 532 450 540 458
rect 562 450 570 458
rect 42 440 50 448
rect 72 440 80 448
rect 102 440 110 448
rect 132 440 140 448
rect 162 440 170 448
rect 192 440 200 448
rect 222 440 230 448
rect 252 440 260 448
rect 282 440 290 448
rect 312 440 320 448
rect 342 440 350 448
rect 372 440 380 448
rect 402 440 410 448
rect 432 440 440 448
rect 462 440 470 448
rect 492 440 500 448
rect 522 440 530 448
rect 552 440 560 448
rect 32 430 40 438
rect 52 430 60 438
rect 82 430 90 438
rect 112 430 120 438
rect 142 430 150 438
rect 172 430 180 438
rect 202 430 210 438
rect 232 430 240 438
rect 262 430 270 438
rect 292 430 300 438
rect 322 430 330 438
rect 352 430 360 438
rect 382 430 390 438
rect 412 430 420 438
rect 442 430 450 438
rect 472 430 480 438
rect 502 430 510 438
rect 532 430 540 438
rect 562 430 570 438
rect 42 420 50 428
rect 72 420 80 428
rect 102 420 110 428
rect 132 420 140 428
rect 162 420 170 428
rect 192 420 200 428
rect 222 420 230 428
rect 252 420 260 428
rect 282 420 290 428
rect 312 420 320 428
rect 342 420 350 428
rect 372 420 380 428
rect 402 420 410 428
rect 432 420 440 428
rect 462 420 470 428
rect 492 420 500 428
rect 522 420 530 428
rect 552 420 560 428
rect 32 410 40 418
rect 52 410 60 418
rect 82 410 90 418
rect 112 410 120 418
rect 142 410 150 418
rect 172 410 180 418
rect 202 410 210 418
rect 232 410 240 418
rect 262 410 270 418
rect 292 410 300 418
rect 322 410 330 418
rect 352 410 360 418
rect 382 410 390 418
rect 412 410 420 418
rect 442 410 450 418
rect 472 410 480 418
rect 502 410 510 418
rect 532 410 540 418
rect 562 410 570 418
rect 42 400 50 408
rect 72 400 80 408
rect 102 400 110 408
rect 132 400 140 408
rect 162 400 170 408
rect 192 400 200 408
rect 222 400 230 408
rect 252 400 260 408
rect 282 400 290 408
rect 312 400 320 408
rect 342 400 350 408
rect 372 400 380 408
rect 402 400 410 408
rect 432 400 440 408
rect 462 400 470 408
rect 492 400 500 408
rect 522 400 530 408
rect 552 400 560 408
rect 32 370 40 398
rect 52 370 60 398
rect 82 370 90 398
rect 112 390 120 398
rect 142 390 150 398
rect 172 390 180 398
rect 202 390 210 398
rect 232 390 240 398
rect 262 390 270 398
rect 292 390 300 398
rect 322 390 330 398
rect 352 390 360 398
rect 382 390 390 398
rect 412 390 420 398
rect 442 390 450 398
rect 472 390 480 398
rect 112 370 120 378
rect 142 370 150 378
rect 172 370 180 378
rect 202 370 210 378
rect 232 370 240 378
rect 262 370 270 378
rect 292 370 300 378
rect 322 370 330 378
rect 352 370 360 378
rect 382 370 390 378
rect 412 370 420 378
rect 442 370 450 378
rect 472 370 480 378
rect 502 370 510 398
rect 532 390 540 398
rect 562 390 570 398
rect 522 380 530 388
rect 552 380 560 388
rect 532 370 540 378
rect 562 370 570 378
rect 42 360 50 368
rect 72 360 80 368
rect 102 360 110 368
rect 132 360 140 368
rect 162 360 170 368
rect 192 360 200 368
rect 222 360 230 368
rect 252 360 260 368
rect 282 360 290 368
rect 312 360 320 368
rect 342 360 350 368
rect 372 360 380 368
rect 402 360 410 368
rect 432 360 440 368
rect 462 360 470 368
rect 492 360 500 368
rect 522 360 530 368
rect 552 360 560 368
rect 32 350 40 358
rect 52 350 60 358
rect 82 350 90 358
rect 112 350 120 358
rect 142 350 150 358
rect 172 350 180 358
rect 202 350 210 358
rect 232 350 240 358
rect 262 350 270 358
rect 292 350 300 358
rect 322 350 330 358
rect 352 350 360 358
rect 382 350 390 358
rect 412 350 420 358
rect 442 350 450 358
rect 472 350 480 358
rect 502 350 510 358
rect 532 350 540 358
rect 562 350 570 358
rect 42 340 50 348
rect 72 340 80 348
rect 102 340 110 348
rect 132 340 140 348
rect 162 340 170 348
rect 192 340 200 348
rect 222 340 230 348
rect 252 340 260 348
rect 282 340 290 348
rect 312 340 320 348
rect 342 340 350 348
rect 372 340 380 348
rect 402 340 410 348
rect 432 340 440 348
rect 462 340 470 348
rect 492 340 500 348
rect 522 340 530 348
rect 552 340 560 348
rect 32 330 40 338
rect 52 330 60 338
rect 82 330 90 338
rect 112 330 120 338
rect 142 330 150 338
rect 172 330 180 338
rect 202 330 210 338
rect 232 330 240 338
rect 262 330 270 338
rect 292 330 300 338
rect 322 330 330 338
rect 352 330 360 338
rect 382 330 390 338
rect 412 330 420 338
rect 442 330 450 338
rect 472 330 480 338
rect 502 330 510 338
rect 532 330 540 338
rect 562 330 570 338
rect 42 320 50 328
rect 72 320 80 328
rect 102 320 110 328
rect 132 320 140 328
rect 162 320 170 328
rect 192 320 200 328
rect 222 320 230 328
rect 252 320 260 328
rect 282 320 290 328
rect 312 320 320 328
rect 342 320 350 328
rect 372 320 380 328
rect 402 320 410 328
rect 432 320 440 328
rect 462 320 470 328
rect 492 320 500 328
rect 522 320 530 328
rect 552 320 560 328
rect 32 310 40 318
rect 52 310 60 318
rect 82 310 90 318
rect 112 310 120 318
rect 142 310 150 318
rect 172 310 180 318
rect 202 310 210 318
rect 232 310 240 318
rect 262 310 270 318
rect 292 310 300 318
rect 322 310 330 318
rect 352 310 360 318
rect 382 310 390 318
rect 412 310 420 318
rect 442 310 450 318
rect 472 310 480 318
rect 502 310 510 318
rect 532 310 540 318
rect 562 310 570 318
rect 42 300 50 308
rect 72 300 80 308
rect 92 300 100 308
rect 522 300 530 308
rect 552 300 560 308
rect 32 290 40 298
rect 52 290 60 298
rect 82 290 90 298
rect 112 290 120 298
rect 142 290 150 298
rect 172 290 180 298
rect 202 290 210 298
rect 232 290 240 298
rect 262 290 270 298
rect 292 290 300 298
rect 322 290 330 298
rect 352 290 360 298
rect 382 290 390 298
rect 412 290 420 298
rect 442 290 450 298
rect 472 290 480 298
rect 502 290 510 298
rect 532 290 540 298
rect 562 290 570 298
rect 42 280 50 288
rect 72 280 80 288
rect 102 280 110 288
rect 132 280 140 288
rect 162 280 170 288
rect 192 280 200 288
rect 222 280 230 288
rect 252 280 260 288
rect 282 280 290 288
rect 312 280 320 288
rect 342 280 350 288
rect 372 280 380 288
rect 402 280 410 288
rect 432 280 440 288
rect 462 280 470 288
rect 492 280 500 288
rect 522 280 530 288
rect 552 280 560 288
rect 32 270 40 278
rect 52 270 60 278
rect 82 270 90 278
rect 112 270 120 278
rect 142 270 150 278
rect 172 270 180 278
rect 202 270 210 278
rect 232 270 240 278
rect 262 270 270 278
rect 292 270 300 278
rect 322 270 330 278
rect 352 270 360 278
rect 382 270 390 278
rect 412 270 420 278
rect 442 270 450 278
rect 472 270 480 278
rect 502 270 510 278
rect 532 270 540 278
rect 562 270 570 278
rect 42 260 50 268
rect 72 260 80 268
rect 102 260 110 268
rect 132 260 140 268
rect 162 260 170 268
rect 192 260 200 268
rect 222 260 230 268
rect 252 260 260 268
rect 282 260 290 268
rect 312 260 320 268
rect 342 260 350 268
rect 372 260 380 268
rect 402 260 410 268
rect 432 260 440 268
rect 462 260 470 268
rect 492 260 500 268
rect 522 260 530 268
rect 552 260 560 268
rect 32 250 40 258
rect 52 250 60 258
rect 82 250 90 258
rect 112 250 120 258
rect 142 250 150 258
rect 172 250 180 258
rect 202 250 210 258
rect 232 250 240 258
rect 262 250 270 258
rect 292 250 300 258
rect 322 250 330 258
rect 352 250 360 258
rect 382 250 390 258
rect 412 250 420 258
rect 442 250 450 258
rect 472 250 480 258
rect 502 250 510 258
rect 532 250 540 258
rect 562 250 570 258
rect 42 240 50 248
rect 32 230 40 238
rect 52 230 60 238
rect 42 220 50 228
rect 72 220 80 248
rect 102 240 110 248
rect 132 240 140 248
rect 162 240 170 248
rect 192 240 200 248
rect 222 240 230 248
rect 252 240 260 248
rect 282 240 290 248
rect 312 240 320 248
rect 342 240 350 248
rect 372 240 380 248
rect 402 240 410 248
rect 432 240 440 248
rect 462 240 470 248
rect 492 240 500 248
rect 522 240 530 248
rect 552 240 560 248
rect 512 230 520 238
rect 532 230 540 238
rect 562 230 570 238
rect 102 220 110 228
rect 132 220 140 228
rect 162 220 170 228
rect 192 220 200 228
rect 222 220 230 228
rect 252 220 260 228
rect 282 220 290 228
rect 312 220 320 228
rect 342 220 350 228
rect 372 220 380 228
rect 402 220 410 228
rect 432 220 440 228
rect 462 220 470 228
rect 492 220 500 228
rect 522 220 530 228
rect 552 220 560 228
rect 32 210 40 218
rect 52 210 60 218
rect 82 210 90 218
rect 112 210 120 218
rect 142 210 150 218
rect 172 210 180 218
rect 202 210 210 218
rect 232 210 240 218
rect 262 210 270 218
rect 292 210 300 218
rect 322 210 330 218
rect 352 210 360 218
rect 382 210 390 218
rect 412 210 420 218
rect 442 210 450 218
rect 472 210 480 218
rect 502 210 510 218
rect 532 210 540 218
rect 562 210 570 218
rect 42 200 50 208
rect 72 200 80 208
rect 102 200 110 208
rect 132 200 140 208
rect 162 200 170 208
rect 192 200 200 208
rect 222 200 230 208
rect 252 200 260 208
rect 282 200 290 208
rect 312 200 320 208
rect 342 200 350 208
rect 372 200 380 208
rect 402 200 410 208
rect 432 200 440 208
rect 462 200 470 208
rect 492 200 500 208
rect 522 200 530 208
rect 552 200 560 208
rect 32 190 40 198
rect 52 190 60 198
rect 82 190 90 198
rect 112 190 120 198
rect 142 190 150 198
rect 172 190 180 198
rect 202 190 210 198
rect 232 190 240 198
rect 262 190 270 198
rect 292 190 300 198
rect 322 190 330 198
rect 352 190 360 198
rect 382 190 390 198
rect 412 190 420 198
rect 442 190 450 198
rect 472 190 480 198
rect 502 190 510 198
rect 532 190 540 198
rect 562 190 570 198
rect 42 180 50 188
rect 72 180 80 188
rect 102 180 110 188
rect 132 180 140 188
rect 162 180 170 188
rect 192 180 200 188
rect 222 180 230 188
rect 252 180 260 188
rect 282 180 290 188
rect 312 180 320 188
rect 342 180 350 188
rect 372 180 380 188
rect 402 180 410 188
rect 432 180 440 188
rect 462 180 470 188
rect 492 180 500 188
rect 522 180 530 188
rect 552 180 560 188
rect 32 170 40 178
rect 52 170 60 178
rect 82 170 90 178
rect 112 170 120 178
rect 142 170 150 178
rect 172 170 180 178
rect 202 170 210 178
rect 232 170 240 178
rect 262 170 270 178
rect 292 170 300 178
rect 322 170 330 178
rect 352 170 360 178
rect 382 170 390 178
rect 412 170 420 178
rect 442 170 450 178
rect 472 170 480 178
rect 502 170 510 178
rect 532 170 540 178
rect 562 170 570 178
rect 42 160 50 168
rect 72 160 80 168
rect 102 160 110 168
rect 132 160 140 168
rect 162 160 170 168
rect 192 160 200 168
rect 222 160 230 168
rect 252 160 260 168
rect 282 160 290 168
rect 312 160 320 168
rect 342 160 350 168
rect 372 160 380 168
rect 402 160 410 168
rect 432 160 440 168
rect 462 160 470 168
rect 492 160 500 168
rect 522 160 530 168
rect 552 160 560 168
rect 32 150 40 158
rect 52 150 60 158
rect 82 150 90 158
rect 512 150 520 158
rect 532 150 540 158
rect 562 150 570 158
rect 42 140 50 148
rect 72 140 80 148
rect 102 140 110 148
rect 132 140 140 148
rect 162 140 170 148
rect 192 140 200 148
rect 222 140 230 148
rect 252 140 260 148
rect 282 140 290 148
rect 312 140 320 148
rect 342 140 350 148
rect 372 140 380 148
rect 402 140 410 148
rect 432 140 440 148
rect 462 140 470 148
rect 492 140 500 148
rect 522 140 530 148
rect 552 140 560 148
rect 32 130 40 138
rect 52 130 60 138
rect 82 130 90 138
rect 112 130 120 138
rect 142 130 150 138
rect 172 130 180 138
rect 202 130 210 138
rect 232 130 240 138
rect 262 130 270 138
rect 292 130 300 138
rect 322 130 330 138
rect 352 130 360 138
rect 382 130 390 138
rect 412 130 420 138
rect 442 130 450 138
rect 472 130 480 138
rect 502 130 510 138
rect 532 130 540 138
rect 562 130 570 138
rect 42 120 50 128
rect 72 120 80 128
rect 102 120 110 128
rect 132 120 140 128
rect 162 120 170 128
rect 192 120 200 128
rect 222 120 230 128
rect 252 120 260 128
rect 282 120 290 128
rect 312 120 320 128
rect 342 120 350 128
rect 372 120 380 128
rect 402 120 410 128
rect 432 120 440 128
rect 462 120 470 128
rect 492 120 500 128
rect 522 120 530 128
rect 552 120 560 128
rect 32 110 40 118
rect 52 110 60 118
rect 82 110 90 118
rect 112 110 120 118
rect 142 110 150 118
rect 172 110 180 118
rect 202 110 210 118
rect 232 110 240 118
rect 262 110 270 118
rect 292 110 300 118
rect 322 110 330 118
rect 352 110 360 118
rect 382 110 390 118
rect 412 110 420 118
rect 442 110 450 118
rect 472 110 480 118
rect 502 110 510 118
rect 532 110 540 118
rect 562 110 570 118
rect 42 100 50 108
rect 72 100 80 108
rect 102 100 110 108
rect 132 100 140 108
rect 162 100 170 108
rect 192 100 200 108
rect 222 100 230 108
rect 252 100 260 108
rect 282 100 290 108
rect 312 100 320 108
rect 342 100 350 108
rect 372 100 380 108
rect 402 100 410 108
rect 432 100 440 108
rect 462 100 470 108
rect 492 100 500 108
rect 522 100 530 108
rect 552 100 560 108
rect 32 90 40 98
rect 52 90 60 98
rect 82 90 90 98
rect 112 90 120 98
rect 142 90 150 98
rect 172 90 180 98
rect 202 90 210 98
rect 232 90 240 98
rect 262 90 270 98
rect 292 90 300 98
rect 322 90 330 98
rect 352 90 360 98
rect 382 90 390 98
rect 412 90 420 98
rect 442 90 450 98
rect 472 90 480 98
rect 502 90 510 98
rect 532 90 540 98
rect 562 90 570 98
rect 42 80 50 88
rect 72 80 80 88
rect 102 80 110 88
rect 132 80 140 88
rect 162 80 170 88
rect 192 80 200 88
rect 222 80 230 88
rect 252 80 260 88
rect 282 80 290 88
rect 312 80 320 88
rect 342 80 350 88
rect 372 80 380 88
rect 402 80 410 88
rect 432 80 440 88
rect 462 80 470 88
rect 492 80 500 88
rect 522 80 530 88
rect 552 80 560 88
rect 32 70 40 78
rect 52 70 60 78
rect 82 70 90 78
rect 112 70 120 78
rect 142 70 150 78
rect 172 70 180 78
rect 202 70 210 78
rect 232 70 240 78
rect 262 70 270 78
rect 292 70 300 78
rect 322 70 330 78
rect 352 70 360 78
rect 382 70 390 78
rect 412 70 420 78
rect 442 70 450 78
rect 472 70 480 78
rect 502 70 510 78
rect 532 70 540 78
rect 562 70 570 78
rect 42 60 50 68
rect 72 60 80 68
rect 102 60 110 68
rect 132 60 140 68
rect 162 60 170 68
rect 192 60 200 68
rect 222 60 230 68
rect 252 60 260 68
rect 282 60 290 68
rect 312 60 320 68
rect 342 60 350 68
rect 372 60 380 68
rect 402 60 410 68
rect 432 60 440 68
rect 462 60 470 68
rect 492 60 500 68
rect 522 60 530 68
rect 552 60 560 68
rect 32 50 40 58
rect 52 50 60 58
rect 82 50 90 58
rect 112 50 120 58
rect 142 50 150 58
rect 172 50 180 58
rect 202 50 210 58
rect 232 50 240 58
rect 262 50 270 58
rect 292 50 300 58
rect 322 50 330 58
rect 352 50 360 58
rect 382 50 390 58
rect 412 50 420 58
rect 442 50 450 58
rect 472 50 480 58
rect 502 50 510 58
rect 532 50 540 58
rect 562 50 570 58
rect 42 40 50 48
rect 72 40 80 48
rect 102 40 110 48
rect 132 40 140 48
rect 162 40 170 48
rect 192 40 200 48
rect 222 40 230 48
rect 252 40 260 48
rect 282 40 290 48
rect 312 40 320 48
rect 342 40 350 48
rect 372 40 380 48
rect 402 40 410 48
rect 432 40 440 48
rect 462 40 470 48
rect 492 40 500 48
rect 522 40 530 48
rect 552 40 560 48
rect 32 30 40 38
rect 52 30 60 38
rect 82 30 90 38
rect 112 30 120 38
rect 142 30 150 38
rect 172 30 180 38
rect 202 30 210 38
rect 232 30 240 38
rect 262 30 270 38
rect 292 30 300 38
rect 322 30 330 38
rect 352 30 360 38
rect 382 30 390 38
rect 412 30 420 38
rect 442 30 450 38
rect 472 30 480 38
rect 502 30 510 38
rect 532 30 540 38
rect 562 30 570 38
<< metal2 >>
rect 0 1298 600 1340
rect 0 1290 56 1298
rect 64 1290 86 1298
rect 94 1290 116 1298
rect 124 1290 146 1298
rect 154 1290 176 1298
rect 184 1290 206 1298
rect 214 1290 236 1298
rect 244 1290 266 1298
rect 274 1290 296 1298
rect 304 1290 326 1298
rect 334 1290 356 1298
rect 364 1290 386 1298
rect 394 1290 416 1298
rect 424 1290 446 1298
rect 454 1290 476 1298
rect 484 1290 506 1298
rect 514 1290 536 1298
rect 544 1290 600 1298
rect 0 1288 600 1290
rect 0 1280 46 1288
rect 54 1280 66 1288
rect 74 1280 96 1288
rect 104 1280 126 1288
rect 134 1280 156 1288
rect 164 1280 186 1288
rect 194 1280 216 1288
rect 224 1280 246 1288
rect 254 1280 276 1288
rect 284 1280 306 1288
rect 314 1280 336 1288
rect 344 1280 366 1288
rect 374 1280 396 1288
rect 404 1280 426 1288
rect 434 1280 456 1288
rect 464 1280 486 1288
rect 494 1280 516 1288
rect 524 1280 546 1288
rect 554 1280 600 1288
rect 0 1278 600 1280
rect 0 1270 56 1278
rect 64 1270 86 1278
rect 94 1270 116 1278
rect 124 1270 146 1278
rect 154 1270 176 1278
rect 184 1270 206 1278
rect 214 1270 236 1278
rect 244 1270 266 1278
rect 274 1270 296 1278
rect 304 1270 326 1278
rect 334 1270 356 1278
rect 364 1270 386 1278
rect 394 1270 416 1278
rect 424 1270 446 1278
rect 454 1270 476 1278
rect 484 1270 506 1278
rect 514 1270 536 1278
rect 544 1270 600 1278
rect 0 1268 600 1270
rect 0 1260 46 1268
rect 54 1260 66 1268
rect 74 1260 96 1268
rect 104 1260 126 1268
rect 134 1260 156 1268
rect 164 1260 186 1268
rect 194 1260 216 1268
rect 224 1260 246 1268
rect 254 1260 276 1268
rect 284 1260 306 1268
rect 314 1260 336 1268
rect 344 1260 366 1268
rect 374 1260 396 1268
rect 404 1260 426 1268
rect 434 1260 456 1268
rect 464 1260 486 1268
rect 494 1260 516 1268
rect 524 1260 546 1268
rect 554 1260 600 1268
rect 0 1258 600 1260
rect 0 1250 56 1258
rect 64 1250 86 1258
rect 94 1250 116 1258
rect 124 1250 146 1258
rect 154 1250 176 1258
rect 184 1250 206 1258
rect 214 1250 236 1258
rect 244 1250 266 1258
rect 274 1250 296 1258
rect 304 1250 326 1258
rect 334 1250 356 1258
rect 364 1250 386 1258
rect 394 1250 416 1258
rect 424 1250 446 1258
rect 454 1250 476 1258
rect 484 1250 506 1258
rect 514 1250 536 1258
rect 544 1250 600 1258
rect 0 1248 600 1250
rect 0 1240 46 1248
rect 54 1240 66 1248
rect 74 1240 96 1248
rect 104 1240 126 1248
rect 134 1240 156 1248
rect 164 1240 186 1248
rect 194 1240 216 1248
rect 224 1240 246 1248
rect 254 1240 276 1248
rect 284 1240 306 1248
rect 314 1240 336 1248
rect 344 1240 366 1248
rect 374 1240 396 1248
rect 404 1240 426 1248
rect 434 1240 456 1248
rect 464 1240 486 1248
rect 494 1240 516 1248
rect 524 1240 546 1248
rect 554 1240 600 1248
rect 0 1238 600 1240
rect 0 1230 56 1238
rect 64 1230 86 1238
rect 94 1230 116 1238
rect 124 1230 146 1238
rect 154 1230 176 1238
rect 184 1230 206 1238
rect 214 1230 236 1238
rect 244 1230 266 1238
rect 274 1230 296 1238
rect 304 1230 326 1238
rect 334 1230 356 1238
rect 364 1230 386 1238
rect 394 1230 416 1238
rect 424 1230 446 1238
rect 454 1230 476 1238
rect 484 1230 506 1238
rect 514 1230 536 1238
rect 544 1230 600 1238
rect 0 1228 600 1230
rect 0 1220 46 1228
rect 54 1220 66 1228
rect 74 1220 96 1228
rect 104 1220 126 1228
rect 134 1220 156 1228
rect 164 1220 186 1228
rect 194 1220 216 1228
rect 224 1220 246 1228
rect 254 1220 276 1228
rect 284 1220 306 1228
rect 314 1220 336 1228
rect 344 1220 366 1228
rect 374 1220 396 1228
rect 404 1220 426 1228
rect 434 1220 456 1228
rect 464 1220 486 1228
rect 494 1220 516 1228
rect 524 1220 546 1228
rect 554 1220 600 1228
rect 0 1218 600 1220
rect 0 1210 56 1218
rect 64 1210 86 1218
rect 94 1210 116 1218
rect 124 1210 146 1218
rect 154 1210 176 1218
rect 184 1210 206 1218
rect 214 1210 236 1218
rect 244 1210 266 1218
rect 274 1210 296 1218
rect 304 1210 326 1218
rect 334 1210 356 1218
rect 364 1210 386 1218
rect 394 1210 416 1218
rect 424 1210 446 1218
rect 454 1210 476 1218
rect 484 1210 506 1218
rect 514 1210 536 1218
rect 544 1210 600 1218
rect 0 1208 600 1210
rect 0 1200 46 1208
rect 54 1200 66 1208
rect 74 1200 96 1208
rect 104 1200 126 1208
rect 134 1200 156 1208
rect 164 1200 186 1208
rect 194 1200 216 1208
rect 224 1200 246 1208
rect 254 1200 276 1208
rect 284 1200 306 1208
rect 314 1200 336 1208
rect 344 1200 366 1208
rect 374 1200 396 1208
rect 404 1200 426 1208
rect 434 1200 456 1208
rect 464 1200 486 1208
rect 494 1200 516 1208
rect 524 1200 546 1208
rect 554 1200 600 1208
rect 0 1198 600 1200
rect 0 1190 56 1198
rect 64 1190 86 1198
rect 94 1190 116 1198
rect 124 1190 146 1198
rect 154 1190 176 1198
rect 184 1190 206 1198
rect 214 1190 236 1198
rect 244 1190 266 1198
rect 274 1190 296 1198
rect 304 1190 326 1198
rect 334 1190 356 1198
rect 364 1190 386 1198
rect 394 1190 416 1198
rect 424 1190 446 1198
rect 454 1190 476 1198
rect 484 1190 506 1198
rect 514 1190 536 1198
rect 544 1190 600 1198
rect 0 1188 100 1190
rect 0 1180 46 1188
rect 54 1180 66 1188
rect 74 1180 100 1188
rect 500 1188 600 1190
rect 500 1180 516 1188
rect 524 1180 546 1188
rect 554 1180 600 1188
rect 0 1178 600 1180
rect 0 1170 56 1178
rect 64 1170 86 1178
rect 94 1170 116 1178
rect 124 1170 146 1178
rect 154 1170 176 1178
rect 184 1170 206 1178
rect 214 1170 236 1178
rect 244 1170 266 1178
rect 274 1170 296 1178
rect 304 1170 326 1178
rect 334 1170 356 1178
rect 364 1170 386 1178
rect 394 1170 416 1178
rect 424 1170 446 1178
rect 454 1170 476 1178
rect 484 1170 506 1178
rect 514 1170 536 1178
rect 544 1170 600 1178
rect 0 1168 600 1170
rect 0 1160 46 1168
rect 54 1160 66 1168
rect 74 1160 96 1168
rect 104 1160 126 1168
rect 134 1160 156 1168
rect 164 1160 186 1168
rect 194 1160 216 1168
rect 224 1160 246 1168
rect 254 1160 276 1168
rect 284 1160 306 1168
rect 314 1160 336 1168
rect 344 1160 366 1168
rect 374 1160 396 1168
rect 404 1160 426 1168
rect 434 1160 456 1168
rect 464 1160 486 1168
rect 494 1160 516 1168
rect 524 1160 546 1168
rect 554 1160 600 1168
rect 0 1158 600 1160
rect 0 1150 56 1158
rect 64 1150 86 1158
rect 94 1150 116 1158
rect 124 1150 146 1158
rect 154 1150 176 1158
rect 184 1150 206 1158
rect 214 1150 236 1158
rect 244 1150 266 1158
rect 274 1150 296 1158
rect 304 1150 326 1158
rect 334 1150 356 1158
rect 364 1150 386 1158
rect 394 1150 416 1158
rect 424 1150 446 1158
rect 454 1150 476 1158
rect 484 1150 506 1158
rect 514 1150 536 1158
rect 544 1150 600 1158
rect 0 1148 600 1150
rect 0 1140 46 1148
rect 54 1140 66 1148
rect 74 1140 96 1148
rect 104 1140 126 1148
rect 134 1140 156 1148
rect 164 1140 186 1148
rect 194 1140 216 1148
rect 224 1140 246 1148
rect 254 1140 276 1148
rect 284 1140 306 1148
rect 314 1140 336 1148
rect 344 1140 366 1148
rect 374 1140 396 1148
rect 404 1140 426 1148
rect 434 1140 456 1148
rect 464 1140 486 1148
rect 494 1140 516 1148
rect 524 1140 546 1148
rect 554 1140 600 1148
rect 0 1138 600 1140
rect 0 1130 56 1138
rect 64 1130 86 1138
rect 94 1130 116 1138
rect 124 1130 146 1138
rect 154 1130 176 1138
rect 184 1130 206 1138
rect 214 1130 236 1138
rect 244 1130 266 1138
rect 274 1130 296 1138
rect 304 1130 326 1138
rect 334 1130 356 1138
rect 364 1130 386 1138
rect 394 1130 416 1138
rect 424 1130 446 1138
rect 454 1130 476 1138
rect 484 1130 506 1138
rect 514 1130 536 1138
rect 544 1130 600 1138
rect 0 1128 600 1130
rect 0 1120 46 1128
rect 54 1120 66 1128
rect 74 1120 96 1128
rect 104 1120 126 1128
rect 134 1120 156 1128
rect 164 1120 186 1128
rect 194 1120 216 1128
rect 224 1120 246 1128
rect 254 1120 276 1128
rect 284 1120 306 1128
rect 314 1120 336 1128
rect 344 1120 366 1128
rect 374 1120 396 1128
rect 404 1120 426 1128
rect 434 1120 456 1128
rect 464 1120 486 1128
rect 494 1120 516 1128
rect 0 1118 516 1120
rect 0 1110 56 1118
rect 64 1110 76 1118
rect 84 1110 516 1118
rect 0 1108 516 1110
rect 0 1100 46 1108
rect 54 1100 66 1108
rect 74 1100 96 1108
rect 104 1100 126 1108
rect 134 1100 156 1108
rect 164 1100 186 1108
rect 194 1100 216 1108
rect 224 1100 246 1108
rect 254 1100 276 1108
rect 284 1100 306 1108
rect 314 1100 336 1108
rect 344 1100 366 1108
rect 374 1100 396 1108
rect 404 1100 426 1108
rect 434 1100 456 1108
rect 464 1100 486 1108
rect 494 1100 516 1108
rect 524 1120 546 1128
rect 554 1120 600 1128
rect 524 1118 600 1120
rect 524 1110 536 1118
rect 544 1110 600 1118
rect 524 1108 600 1110
rect 524 1100 546 1108
rect 554 1100 600 1108
rect 0 1098 600 1100
rect 0 1090 56 1098
rect 64 1090 86 1098
rect 94 1090 116 1098
rect 124 1090 146 1098
rect 154 1090 176 1098
rect 184 1090 206 1098
rect 214 1090 236 1098
rect 244 1090 266 1098
rect 274 1090 296 1098
rect 304 1090 326 1098
rect 334 1090 356 1098
rect 364 1090 386 1098
rect 394 1090 416 1098
rect 424 1090 446 1098
rect 454 1090 476 1098
rect 484 1090 506 1098
rect 514 1090 536 1098
rect 544 1090 600 1098
rect 0 1088 600 1090
rect 0 1080 46 1088
rect 54 1080 66 1088
rect 74 1080 96 1088
rect 104 1080 126 1088
rect 134 1080 156 1088
rect 164 1080 186 1088
rect 194 1080 216 1088
rect 224 1080 246 1088
rect 254 1080 276 1088
rect 284 1080 306 1088
rect 314 1080 336 1088
rect 344 1080 366 1088
rect 374 1080 396 1088
rect 404 1080 426 1088
rect 434 1080 456 1088
rect 464 1080 486 1088
rect 494 1080 516 1088
rect 524 1080 546 1088
rect 554 1080 600 1088
rect 0 1078 600 1080
rect 0 1070 56 1078
rect 64 1070 86 1078
rect 94 1070 116 1078
rect 124 1070 146 1078
rect 154 1070 176 1078
rect 184 1070 206 1078
rect 214 1070 236 1078
rect 244 1070 266 1078
rect 274 1070 296 1078
rect 304 1070 326 1078
rect 334 1070 356 1078
rect 364 1070 386 1078
rect 394 1070 416 1078
rect 424 1070 446 1078
rect 454 1070 476 1078
rect 484 1070 506 1078
rect 514 1070 536 1078
rect 544 1070 600 1078
rect 0 1068 600 1070
rect 0 1060 46 1068
rect 54 1060 66 1068
rect 74 1060 96 1068
rect 104 1060 126 1068
rect 134 1060 156 1068
rect 164 1060 186 1068
rect 194 1060 216 1068
rect 224 1060 246 1068
rect 254 1060 276 1068
rect 284 1060 306 1068
rect 314 1060 336 1068
rect 344 1060 366 1068
rect 374 1060 396 1068
rect 404 1060 426 1068
rect 434 1060 456 1068
rect 464 1060 486 1068
rect 494 1060 516 1068
rect 524 1060 546 1068
rect 554 1060 600 1068
rect 0 1058 600 1060
rect 0 1050 56 1058
rect 64 1050 86 1058
rect 94 1050 116 1058
rect 124 1050 146 1058
rect 154 1050 176 1058
rect 184 1050 206 1058
rect 214 1050 236 1058
rect 244 1050 266 1058
rect 274 1050 296 1058
rect 304 1050 326 1058
rect 334 1050 356 1058
rect 364 1050 386 1058
rect 394 1050 416 1058
rect 424 1050 446 1058
rect 454 1050 476 1058
rect 484 1050 506 1058
rect 514 1050 536 1058
rect 544 1050 600 1058
rect 0 1048 600 1050
rect 0 1040 46 1048
rect 54 1040 66 1048
rect 74 1040 96 1048
rect 104 1040 126 1048
rect 134 1040 156 1048
rect 164 1040 186 1048
rect 194 1040 216 1048
rect 224 1040 246 1048
rect 254 1040 276 1048
rect 284 1040 306 1048
rect 314 1040 336 1048
rect 344 1040 366 1048
rect 374 1040 396 1048
rect 404 1040 426 1048
rect 434 1040 456 1048
rect 464 1040 486 1048
rect 494 1040 516 1048
rect 0 1038 100 1040
rect 0 1030 56 1038
rect 64 1030 86 1038
rect 94 1030 100 1038
rect 500 1030 516 1040
rect 0 1028 516 1030
rect 0 1020 46 1028
rect 54 1020 66 1028
rect 74 1020 96 1028
rect 104 1020 126 1028
rect 134 1020 156 1028
rect 164 1020 186 1028
rect 194 1020 216 1028
rect 224 1020 246 1028
rect 254 1020 276 1028
rect 284 1020 306 1028
rect 314 1020 336 1028
rect 344 1020 366 1028
rect 374 1020 396 1028
rect 404 1020 426 1028
rect 434 1020 456 1028
rect 464 1020 486 1028
rect 494 1020 516 1028
rect 524 1040 546 1048
rect 554 1040 600 1048
rect 524 1038 600 1040
rect 524 1030 536 1038
rect 544 1030 600 1038
rect 524 1028 600 1030
rect 524 1020 546 1028
rect 554 1020 600 1028
rect 0 1018 600 1020
rect 0 1010 56 1018
rect 64 1010 86 1018
rect 94 1010 116 1018
rect 124 1010 146 1018
rect 154 1010 176 1018
rect 184 1010 206 1018
rect 214 1010 236 1018
rect 244 1010 266 1018
rect 274 1010 296 1018
rect 304 1010 326 1018
rect 334 1010 356 1018
rect 364 1010 386 1018
rect 394 1010 416 1018
rect 424 1010 446 1018
rect 454 1010 476 1018
rect 484 1010 506 1018
rect 514 1010 536 1018
rect 544 1010 600 1018
rect 0 1008 600 1010
rect 0 1000 46 1008
rect 54 1000 66 1008
rect 74 1000 96 1008
rect 104 1000 126 1008
rect 134 1000 156 1008
rect 164 1000 186 1008
rect 194 1000 216 1008
rect 224 1000 246 1008
rect 254 1000 276 1008
rect 284 1000 306 1008
rect 314 1000 336 1008
rect 344 1000 366 1008
rect 374 1000 396 1008
rect 404 1000 426 1008
rect 434 1000 456 1008
rect 464 1000 486 1008
rect 494 1000 516 1008
rect 524 1000 546 1008
rect 554 1000 600 1008
rect 0 998 600 1000
rect 0 990 56 998
rect 64 990 86 998
rect 94 990 116 998
rect 124 990 146 998
rect 154 990 176 998
rect 184 990 206 998
rect 214 990 236 998
rect 244 990 266 998
rect 274 990 296 998
rect 304 990 326 998
rect 334 990 356 998
rect 364 990 386 998
rect 394 990 416 998
rect 424 990 446 998
rect 454 990 476 998
rect 484 990 506 998
rect 514 990 536 998
rect 544 990 600 998
rect 0 988 600 990
rect 0 980 46 988
rect 54 980 66 988
rect 74 980 96 988
rect 104 980 126 988
rect 134 980 156 988
rect 164 980 186 988
rect 194 980 216 988
rect 224 980 246 988
rect 254 980 276 988
rect 284 980 306 988
rect 314 980 336 988
rect 344 980 366 988
rect 374 980 396 988
rect 404 980 426 988
rect 434 980 456 988
rect 464 980 486 988
rect 494 980 516 988
rect 524 980 546 988
rect 554 980 600 988
rect 0 978 600 980
rect 0 970 56 978
rect 64 970 86 978
rect 94 970 116 978
rect 124 970 146 978
rect 154 970 176 978
rect 184 970 206 978
rect 214 970 236 978
rect 244 970 266 978
rect 274 970 296 978
rect 304 970 326 978
rect 334 970 356 978
rect 364 970 386 978
rect 394 970 416 978
rect 424 970 446 978
rect 454 970 476 978
rect 484 970 506 978
rect 514 970 536 978
rect 544 970 600 978
rect 0 968 600 970
rect 0 960 46 968
rect 54 960 546 968
rect 554 960 600 968
rect 0 958 600 960
rect 0 950 56 958
rect 64 950 86 958
rect 94 950 116 958
rect 124 950 146 958
rect 154 950 176 958
rect 184 950 206 958
rect 214 950 236 958
rect 244 950 266 958
rect 274 950 296 958
rect 304 950 326 958
rect 334 950 356 958
rect 364 950 386 958
rect 394 950 416 958
rect 424 950 446 958
rect 454 950 476 958
rect 484 950 506 958
rect 514 950 536 958
rect 544 950 600 958
rect 0 948 600 950
rect 0 940 46 948
rect 54 940 66 948
rect 74 940 96 948
rect 104 940 126 948
rect 134 940 156 948
rect 164 940 186 948
rect 194 940 216 948
rect 224 940 246 948
rect 254 940 276 948
rect 284 940 306 948
rect 314 940 336 948
rect 344 940 366 948
rect 374 940 396 948
rect 404 940 426 948
rect 434 940 456 948
rect 464 940 486 948
rect 494 940 516 948
rect 524 940 546 948
rect 554 940 600 948
rect 0 938 600 940
rect 0 930 56 938
rect 64 930 86 938
rect 94 930 116 938
rect 124 930 146 938
rect 154 930 176 938
rect 184 930 206 938
rect 214 930 236 938
rect 244 930 266 938
rect 274 930 296 938
rect 304 930 326 938
rect 334 930 356 938
rect 364 930 386 938
rect 394 930 416 938
rect 424 930 446 938
rect 454 930 476 938
rect 484 930 506 938
rect 514 930 536 938
rect 544 930 600 938
rect 0 928 600 930
rect 0 920 46 928
rect 54 920 66 928
rect 74 920 96 928
rect 104 920 126 928
rect 134 920 156 928
rect 164 920 186 928
rect 194 920 216 928
rect 224 920 246 928
rect 254 920 276 928
rect 284 920 306 928
rect 314 920 336 928
rect 344 920 366 928
rect 374 920 396 928
rect 404 920 426 928
rect 434 920 456 928
rect 464 920 486 928
rect 494 920 516 928
rect 524 920 546 928
rect 554 920 600 928
rect 0 918 600 920
rect 0 910 56 918
rect 64 910 86 918
rect 94 910 116 918
rect 124 910 146 918
rect 154 910 176 918
rect 184 910 206 918
rect 214 910 236 918
rect 244 910 266 918
rect 274 910 296 918
rect 304 910 326 918
rect 334 910 356 918
rect 364 910 386 918
rect 394 910 416 918
rect 424 910 446 918
rect 454 910 476 918
rect 484 910 506 918
rect 514 910 536 918
rect 544 910 600 918
rect 0 908 600 910
rect 0 900 46 908
rect 54 900 66 908
rect 74 900 96 908
rect 104 900 126 908
rect 134 900 156 908
rect 164 900 186 908
rect 194 900 216 908
rect 224 900 246 908
rect 254 900 276 908
rect 284 900 306 908
rect 314 900 336 908
rect 344 900 366 908
rect 374 900 396 908
rect 404 900 426 908
rect 434 900 456 908
rect 464 900 486 908
rect 494 900 516 908
rect 524 900 546 908
rect 554 900 600 908
rect 0 898 600 900
rect 0 890 56 898
rect 64 890 86 898
rect 94 890 116 898
rect 124 890 146 898
rect 154 890 176 898
rect 184 890 206 898
rect 214 890 236 898
rect 244 890 266 898
rect 274 890 296 898
rect 304 890 326 898
rect 334 890 356 898
rect 364 890 386 898
rect 394 890 416 898
rect 424 890 446 898
rect 454 890 476 898
rect 484 890 506 898
rect 514 890 536 898
rect 544 890 600 898
rect 0 888 600 890
rect 0 880 46 888
rect 54 880 66 888
rect 74 880 96 888
rect 104 880 126 888
rect 134 880 156 888
rect 164 880 186 888
rect 194 880 216 888
rect 224 880 246 888
rect 254 880 276 888
rect 284 880 306 888
rect 314 880 336 888
rect 344 880 366 888
rect 374 880 396 888
rect 404 880 426 888
rect 434 880 456 888
rect 464 880 486 888
rect 494 880 516 888
rect 524 880 546 888
rect 554 880 600 888
rect 0 836 600 848
rect 0 828 14 836
rect 22 828 44 836
rect 52 828 74 836
rect 82 828 104 836
rect 112 828 134 836
rect 142 828 164 836
rect 172 828 194 836
rect 202 828 224 836
rect 232 828 244 836
rect 252 828 266 836
rect 274 828 296 836
rect 304 828 326 836
rect 334 828 348 836
rect 356 828 368 836
rect 376 828 398 836
rect 406 828 428 836
rect 436 828 458 836
rect 466 828 488 836
rect 496 828 518 836
rect 526 828 548 836
rect 556 828 578 836
rect 586 828 600 836
rect 0 826 600 828
rect 0 818 4 826
rect 12 818 24 826
rect 32 818 54 826
rect 62 818 84 826
rect 92 818 114 826
rect 122 818 144 826
rect 152 818 174 826
rect 182 818 204 826
rect 212 818 234 826
rect 242 818 256 826
rect 264 818 276 826
rect 284 818 306 826
rect 314 818 336 826
rect 344 818 358 826
rect 366 818 388 826
rect 396 818 418 826
rect 426 818 448 826
rect 456 818 478 826
rect 486 818 508 826
rect 516 818 538 826
rect 546 818 568 826
rect 576 818 588 826
rect 596 818 600 826
rect 0 816 600 818
rect 0 808 14 816
rect 22 808 44 816
rect 52 808 74 816
rect 82 808 104 816
rect 112 808 134 816
rect 142 808 164 816
rect 172 808 194 816
rect 202 808 224 816
rect 232 808 244 816
rect 252 808 266 816
rect 274 808 296 816
rect 304 808 326 816
rect 334 808 348 816
rect 356 808 368 816
rect 376 808 398 816
rect 406 808 428 816
rect 436 808 458 816
rect 466 808 488 816
rect 496 808 518 816
rect 526 808 548 816
rect 556 808 578 816
rect 586 808 600 816
rect 0 806 600 808
rect 0 798 4 806
rect 12 798 24 806
rect 32 798 54 806
rect 62 798 84 806
rect 92 798 114 806
rect 122 798 144 806
rect 152 798 174 806
rect 182 798 204 806
rect 212 798 234 806
rect 242 798 256 806
rect 264 798 276 806
rect 284 798 306 806
rect 314 798 336 806
rect 344 798 358 806
rect 366 798 388 806
rect 396 798 418 806
rect 426 798 448 806
rect 456 798 478 806
rect 486 798 508 806
rect 516 798 538 806
rect 546 798 568 806
rect 576 798 588 806
rect 596 798 600 806
rect 0 796 600 798
rect 0 788 14 796
rect 22 788 44 796
rect 52 788 74 796
rect 82 788 104 796
rect 112 788 134 796
rect 142 788 164 796
rect 172 788 194 796
rect 202 788 224 796
rect 232 788 244 796
rect 252 788 266 796
rect 274 788 296 796
rect 304 788 326 796
rect 334 788 348 796
rect 356 788 368 796
rect 376 788 398 796
rect 406 788 428 796
rect 436 788 458 796
rect 466 788 488 796
rect 496 788 518 796
rect 526 788 548 796
rect 556 788 578 796
rect 586 788 600 796
rect 0 786 600 788
rect 0 778 4 786
rect 12 778 24 786
rect 32 778 54 786
rect 62 778 84 786
rect 92 778 114 786
rect 122 778 144 786
rect 152 778 174 786
rect 182 778 204 786
rect 212 778 234 786
rect 242 778 256 786
rect 264 778 276 786
rect 284 778 306 786
rect 314 778 336 786
rect 344 778 358 786
rect 366 778 388 786
rect 396 778 418 786
rect 426 778 448 786
rect 456 778 478 786
rect 486 778 508 786
rect 516 778 538 786
rect 546 778 568 786
rect 576 778 588 786
rect 596 778 600 786
rect 0 776 100 778
rect 0 768 14 776
rect 22 768 44 776
rect 52 768 74 776
rect 82 768 100 776
rect 500 776 600 778
rect 500 768 518 776
rect 526 768 548 776
rect 556 768 578 776
rect 586 768 600 776
rect 0 766 600 768
rect 0 758 4 766
rect 12 758 24 766
rect 32 758 54 766
rect 62 758 84 766
rect 92 758 114 766
rect 122 758 144 766
rect 152 758 174 766
rect 182 758 204 766
rect 212 758 234 766
rect 242 758 256 766
rect 264 758 276 766
rect 284 758 306 766
rect 314 758 336 766
rect 344 758 358 766
rect 366 758 388 766
rect 396 758 418 766
rect 426 758 448 766
rect 456 758 478 766
rect 486 758 508 766
rect 516 758 538 766
rect 546 758 568 766
rect 576 758 588 766
rect 596 758 600 766
rect 0 756 600 758
rect 0 748 14 756
rect 22 748 44 756
rect 52 748 74 756
rect 82 748 104 756
rect 112 748 134 756
rect 142 748 164 756
rect 172 748 194 756
rect 202 748 224 756
rect 232 748 244 756
rect 252 748 266 756
rect 274 748 296 756
rect 304 748 326 756
rect 334 748 348 756
rect 356 748 368 756
rect 376 748 398 756
rect 406 748 428 756
rect 436 748 458 756
rect 466 748 488 756
rect 496 748 518 756
rect 526 748 548 756
rect 556 748 578 756
rect 586 748 600 756
rect 0 746 600 748
rect 0 738 4 746
rect 12 738 24 746
rect 32 738 54 746
rect 62 738 84 746
rect 92 738 114 746
rect 122 738 144 746
rect 152 738 174 746
rect 182 738 204 746
rect 212 738 234 746
rect 242 738 256 746
rect 264 738 276 746
rect 284 738 306 746
rect 314 738 336 746
rect 344 738 358 746
rect 366 738 388 746
rect 396 738 418 746
rect 426 738 448 746
rect 456 738 478 746
rect 486 738 508 746
rect 516 738 538 746
rect 546 738 568 746
rect 576 738 588 746
rect 596 738 600 746
rect 0 736 600 738
rect 0 728 14 736
rect 22 728 224 736
rect 232 728 244 736
rect 252 728 266 736
rect 274 728 296 736
rect 304 728 326 736
rect 334 728 348 736
rect 356 728 368 736
rect 376 728 578 736
rect 586 728 600 736
rect 0 726 600 728
rect 0 718 4 726
rect 12 718 24 726
rect 32 718 54 726
rect 62 718 84 726
rect 92 718 114 726
rect 122 718 144 726
rect 152 718 174 726
rect 182 718 204 726
rect 212 718 234 726
rect 242 718 256 726
rect 264 718 276 726
rect 284 718 306 726
rect 314 718 336 726
rect 344 718 358 726
rect 366 718 388 726
rect 396 718 418 726
rect 426 718 448 726
rect 456 718 478 726
rect 486 718 508 726
rect 516 718 538 726
rect 546 718 568 726
rect 576 718 588 726
rect 596 718 600 726
rect 0 716 600 718
rect 0 708 14 716
rect 22 708 44 716
rect 52 708 74 716
rect 82 708 104 716
rect 112 708 134 716
rect 142 708 164 716
rect 172 708 194 716
rect 202 708 224 716
rect 232 708 244 716
rect 252 708 266 716
rect 274 708 296 716
rect 304 708 326 716
rect 334 708 348 716
rect 356 708 368 716
rect 376 708 398 716
rect 406 708 428 716
rect 436 708 458 716
rect 466 708 488 716
rect 496 708 518 716
rect 526 708 548 716
rect 556 708 578 716
rect 586 708 600 716
rect 0 706 600 708
rect 0 698 4 706
rect 12 698 24 706
rect 32 698 54 706
rect 62 698 84 706
rect 92 698 114 706
rect 122 698 144 706
rect 152 698 174 706
rect 182 698 204 706
rect 212 698 234 706
rect 242 698 256 706
rect 264 698 276 706
rect 284 698 306 706
rect 314 698 336 706
rect 344 698 358 706
rect 366 698 388 706
rect 396 698 418 706
rect 426 698 448 706
rect 456 698 478 706
rect 486 698 508 706
rect 516 698 538 706
rect 546 698 568 706
rect 576 698 588 706
rect 596 698 600 706
rect 0 696 600 698
rect 0 688 14 696
rect 22 688 44 696
rect 52 688 74 696
rect 82 688 104 696
rect 112 688 134 696
rect 142 688 164 696
rect 172 688 194 696
rect 202 688 224 696
rect 232 688 244 696
rect 252 688 266 696
rect 274 688 296 696
rect 304 688 326 696
rect 334 688 348 696
rect 356 688 368 696
rect 376 688 398 696
rect 406 688 428 696
rect 436 688 458 696
rect 466 688 488 696
rect 496 688 518 696
rect 526 688 548 696
rect 556 688 578 696
rect 586 688 600 696
rect 0 644 14 652
rect 22 644 44 652
rect 52 644 74 652
rect 82 644 104 652
rect 112 644 134 652
rect 142 644 164 652
rect 172 644 194 652
rect 202 644 224 652
rect 232 644 244 652
rect 252 644 266 652
rect 274 644 296 652
rect 304 644 326 652
rect 334 644 348 652
rect 356 644 368 652
rect 376 644 398 652
rect 406 644 428 652
rect 436 644 458 652
rect 466 644 488 652
rect 496 644 518 652
rect 526 644 548 652
rect 556 644 578 652
rect 586 644 600 652
rect 0 642 600 644
rect 0 634 4 642
rect 12 634 24 642
rect 32 634 54 642
rect 62 634 84 642
rect 92 634 114 642
rect 122 634 144 642
rect 152 634 174 642
rect 182 634 204 642
rect 212 634 234 642
rect 242 634 256 642
rect 264 634 276 642
rect 284 634 306 642
rect 314 634 336 642
rect 344 634 358 642
rect 366 634 388 642
rect 396 634 418 642
rect 426 634 448 642
rect 456 634 478 642
rect 486 634 508 642
rect 516 634 538 642
rect 546 634 568 642
rect 576 634 588 642
rect 596 634 600 642
rect 0 632 600 634
rect 0 624 14 632
rect 22 624 44 632
rect 52 624 74 632
rect 82 624 104 632
rect 112 624 134 632
rect 142 624 164 632
rect 172 624 194 632
rect 202 624 224 632
rect 232 624 244 632
rect 252 624 266 632
rect 274 624 296 632
rect 304 624 326 632
rect 334 624 348 632
rect 356 624 368 632
rect 376 624 398 632
rect 406 624 428 632
rect 436 624 458 632
rect 466 624 488 632
rect 496 624 518 632
rect 526 624 548 632
rect 556 624 578 632
rect 586 624 600 632
rect 0 622 600 624
rect 0 614 4 622
rect 12 614 24 622
rect 32 614 54 622
rect 62 614 84 622
rect 92 614 114 622
rect 122 614 144 622
rect 152 614 174 622
rect 182 614 204 622
rect 212 614 234 622
rect 242 614 256 622
rect 264 614 276 622
rect 284 614 306 622
rect 314 614 336 622
rect 344 614 358 622
rect 366 614 388 622
rect 396 614 418 622
rect 426 614 448 622
rect 456 614 478 622
rect 486 614 508 622
rect 516 614 538 622
rect 546 614 568 622
rect 576 614 588 622
rect 596 614 600 622
rect 0 612 600 614
rect 0 604 14 612
rect 22 604 224 612
rect 232 604 244 612
rect 252 604 266 612
rect 274 604 296 612
rect 304 604 326 612
rect 334 604 348 612
rect 356 604 368 612
rect 376 604 578 612
rect 586 604 600 612
rect 0 602 600 604
rect 0 594 4 602
rect 12 594 24 602
rect 32 594 54 602
rect 62 594 84 602
rect 92 594 114 602
rect 122 594 144 602
rect 152 594 174 602
rect 182 594 204 602
rect 212 594 234 602
rect 242 594 256 602
rect 264 594 276 602
rect 284 594 306 602
rect 314 594 336 602
rect 344 594 358 602
rect 366 594 388 602
rect 396 594 418 602
rect 426 594 448 602
rect 456 594 478 602
rect 486 594 508 602
rect 516 594 538 602
rect 546 594 568 602
rect 576 594 588 602
rect 596 594 600 602
rect 0 592 600 594
rect 0 584 14 592
rect 22 584 44 592
rect 52 584 74 592
rect 82 584 104 592
rect 112 584 134 592
rect 142 584 164 592
rect 172 584 194 592
rect 202 584 224 592
rect 232 584 244 592
rect 252 584 348 592
rect 356 584 368 592
rect 376 584 398 592
rect 406 584 428 592
rect 436 584 458 592
rect 466 584 488 592
rect 496 584 518 592
rect 526 584 548 592
rect 556 584 578 592
rect 586 584 600 592
rect 0 582 600 584
rect 0 574 4 582
rect 12 574 24 582
rect 32 574 54 582
rect 62 574 84 582
rect 92 574 100 582
rect 0 572 100 574
rect 500 574 508 582
rect 516 574 538 582
rect 546 574 568 582
rect 576 574 588 582
rect 596 574 600 582
rect 500 572 600 574
rect 0 564 14 572
rect 22 564 44 572
rect 52 564 74 572
rect 82 564 104 572
rect 112 564 134 572
rect 142 564 164 572
rect 172 564 194 572
rect 202 564 224 572
rect 232 564 244 572
rect 252 564 266 572
rect 274 564 296 572
rect 304 564 326 572
rect 334 564 348 572
rect 356 564 368 572
rect 376 564 398 572
rect 406 564 428 572
rect 436 564 458 572
rect 466 564 488 572
rect 496 564 518 572
rect 526 564 548 572
rect 556 564 578 572
rect 586 564 600 572
rect 0 562 600 564
rect 0 554 4 562
rect 12 554 24 562
rect 32 554 54 562
rect 62 554 84 562
rect 92 554 114 562
rect 122 554 144 562
rect 152 554 174 562
rect 182 554 204 562
rect 212 554 234 562
rect 242 554 256 562
rect 264 554 276 562
rect 284 554 306 562
rect 314 554 336 562
rect 344 554 358 562
rect 366 554 388 562
rect 396 554 418 562
rect 426 554 448 562
rect 456 554 478 562
rect 486 554 508 562
rect 516 554 538 562
rect 546 554 568 562
rect 576 554 588 562
rect 596 554 600 562
rect 0 552 600 554
rect 0 544 14 552
rect 22 544 44 552
rect 52 544 74 552
rect 82 544 104 552
rect 112 544 134 552
rect 142 544 164 552
rect 172 544 194 552
rect 202 544 224 552
rect 232 544 244 552
rect 252 544 266 552
rect 274 544 296 552
rect 304 544 326 552
rect 334 544 348 552
rect 356 544 368 552
rect 376 544 398 552
rect 406 544 428 552
rect 436 544 458 552
rect 466 544 488 552
rect 496 544 518 552
rect 526 544 548 552
rect 556 544 578 552
rect 586 544 600 552
rect 0 542 600 544
rect 0 534 4 542
rect 12 534 24 542
rect 32 534 54 542
rect 62 534 84 542
rect 92 534 114 542
rect 122 534 144 542
rect 152 534 174 542
rect 182 534 204 542
rect 212 534 234 542
rect 242 534 256 542
rect 264 534 276 542
rect 284 534 306 542
rect 314 534 336 542
rect 344 534 358 542
rect 366 534 388 542
rect 396 534 418 542
rect 426 534 448 542
rect 456 534 478 542
rect 486 534 508 542
rect 516 534 538 542
rect 546 534 568 542
rect 576 534 588 542
rect 596 534 600 542
rect 0 532 600 534
rect 0 524 14 532
rect 22 524 44 532
rect 52 524 74 532
rect 82 524 104 532
rect 112 524 134 532
rect 142 524 164 532
rect 172 524 194 532
rect 202 524 224 532
rect 232 524 244 532
rect 252 524 266 532
rect 274 524 296 532
rect 304 524 326 532
rect 334 524 348 532
rect 356 524 368 532
rect 376 524 398 532
rect 406 524 428 532
rect 436 524 458 532
rect 466 524 488 532
rect 496 524 518 532
rect 526 524 548 532
rect 556 524 578 532
rect 586 524 600 532
rect 0 516 600 524
rect 0 508 14 516
rect 22 508 34 516
rect 42 508 54 516
rect 62 508 74 516
rect 82 508 94 516
rect 102 508 114 516
rect 122 508 134 516
rect 142 508 154 516
rect 162 508 174 516
rect 182 508 194 516
rect 202 508 214 516
rect 222 508 234 516
rect 242 508 254 516
rect 262 508 274 516
rect 282 508 294 516
rect 302 508 308 516
rect 316 508 328 516
rect 336 508 348 516
rect 356 508 368 516
rect 376 508 388 516
rect 396 508 408 516
rect 416 508 428 516
rect 436 508 448 516
rect 456 508 468 516
rect 476 508 488 516
rect 496 508 508 516
rect 516 508 528 516
rect 536 508 548 516
rect 556 508 568 516
rect 576 508 600 516
rect 0 492 600 508
rect 0 458 600 460
rect 0 450 32 458
rect 40 450 52 458
rect 60 450 82 458
rect 90 450 112 458
rect 120 450 142 458
rect 150 450 172 458
rect 180 450 202 458
rect 210 450 232 458
rect 240 450 262 458
rect 270 450 292 458
rect 300 450 322 458
rect 330 450 352 458
rect 360 450 382 458
rect 390 450 412 458
rect 420 450 442 458
rect 450 450 472 458
rect 480 450 502 458
rect 510 450 532 458
rect 540 450 562 458
rect 570 450 600 458
rect 0 448 600 450
rect 0 440 42 448
rect 50 440 72 448
rect 80 440 102 448
rect 110 440 132 448
rect 140 440 162 448
rect 170 440 192 448
rect 200 440 222 448
rect 230 440 252 448
rect 260 440 282 448
rect 290 440 312 448
rect 320 440 342 448
rect 350 440 372 448
rect 380 440 402 448
rect 410 440 432 448
rect 440 440 462 448
rect 470 440 492 448
rect 500 440 522 448
rect 530 440 552 448
rect 560 440 600 448
rect 0 438 600 440
rect 0 430 32 438
rect 40 430 52 438
rect 60 430 82 438
rect 90 430 112 438
rect 120 430 142 438
rect 150 430 172 438
rect 180 430 202 438
rect 210 430 232 438
rect 240 430 262 438
rect 270 430 292 438
rect 300 430 322 438
rect 330 430 352 438
rect 360 430 382 438
rect 390 430 412 438
rect 420 430 442 438
rect 450 430 472 438
rect 480 430 502 438
rect 510 430 532 438
rect 540 430 562 438
rect 570 430 600 438
rect 0 428 600 430
rect 0 420 42 428
rect 50 420 72 428
rect 80 420 102 428
rect 110 420 132 428
rect 140 420 162 428
rect 170 420 192 428
rect 200 420 222 428
rect 230 420 252 428
rect 260 420 282 428
rect 290 420 312 428
rect 320 420 342 428
rect 350 420 372 428
rect 380 420 402 428
rect 410 420 432 428
rect 440 420 462 428
rect 470 420 492 428
rect 500 420 522 428
rect 530 420 552 428
rect 560 420 600 428
rect 0 418 600 420
rect 0 410 32 418
rect 40 410 52 418
rect 60 410 82 418
rect 90 410 112 418
rect 120 410 142 418
rect 150 410 172 418
rect 180 410 202 418
rect 210 410 232 418
rect 240 410 262 418
rect 270 410 292 418
rect 300 410 322 418
rect 330 410 352 418
rect 360 410 382 418
rect 390 410 412 418
rect 420 410 442 418
rect 450 410 472 418
rect 480 410 502 418
rect 510 410 532 418
rect 540 410 562 418
rect 570 410 600 418
rect 0 408 600 410
rect 0 400 42 408
rect 50 400 72 408
rect 80 400 102 408
rect 110 400 132 408
rect 140 400 162 408
rect 170 400 192 408
rect 200 400 222 408
rect 230 400 252 408
rect 260 400 282 408
rect 290 400 312 408
rect 320 400 342 408
rect 350 400 372 408
rect 380 400 402 408
rect 410 400 432 408
rect 440 400 462 408
rect 470 400 492 408
rect 500 400 522 408
rect 530 400 552 408
rect 560 400 600 408
rect 0 398 600 400
rect 0 370 32 398
rect 40 370 52 398
rect 60 370 82 398
rect 90 390 112 398
rect 120 390 142 398
rect 150 390 172 398
rect 180 390 202 398
rect 210 390 232 398
rect 240 390 262 398
rect 270 390 292 398
rect 300 390 322 398
rect 330 390 352 398
rect 360 390 382 398
rect 390 390 412 398
rect 420 390 442 398
rect 450 390 472 398
rect 480 390 502 398
rect 90 378 502 390
rect 90 370 112 378
rect 120 370 142 378
rect 150 370 172 378
rect 180 370 202 378
rect 210 370 232 378
rect 240 370 262 378
rect 270 370 292 378
rect 300 370 322 378
rect 330 370 352 378
rect 360 370 382 378
rect 390 370 412 378
rect 420 370 442 378
rect 450 370 472 378
rect 480 370 502 378
rect 510 390 532 398
rect 540 390 562 398
rect 570 390 600 398
rect 510 388 600 390
rect 510 380 522 388
rect 530 380 552 388
rect 560 380 600 388
rect 510 378 600 380
rect 510 370 532 378
rect 540 370 562 378
rect 570 370 600 378
rect 0 368 600 370
rect 0 360 42 368
rect 50 360 72 368
rect 80 360 102 368
rect 110 360 132 368
rect 140 360 162 368
rect 170 360 192 368
rect 200 360 222 368
rect 230 360 252 368
rect 260 360 282 368
rect 290 360 312 368
rect 320 360 342 368
rect 350 360 372 368
rect 380 360 402 368
rect 410 360 432 368
rect 440 360 462 368
rect 470 360 492 368
rect 500 360 522 368
rect 530 360 552 368
rect 560 360 600 368
rect 0 358 600 360
rect 0 350 32 358
rect 40 350 52 358
rect 60 350 82 358
rect 90 350 112 358
rect 120 350 142 358
rect 150 350 172 358
rect 180 350 202 358
rect 210 350 232 358
rect 240 350 262 358
rect 270 350 292 358
rect 300 350 322 358
rect 330 350 352 358
rect 360 350 382 358
rect 390 350 412 358
rect 420 350 442 358
rect 450 350 472 358
rect 480 350 502 358
rect 510 350 532 358
rect 540 350 562 358
rect 570 350 600 358
rect 0 348 600 350
rect 0 340 42 348
rect 50 340 72 348
rect 80 340 102 348
rect 110 340 132 348
rect 140 340 162 348
rect 170 340 192 348
rect 200 340 222 348
rect 230 340 252 348
rect 260 340 282 348
rect 290 340 312 348
rect 320 340 342 348
rect 350 340 372 348
rect 380 340 402 348
rect 410 340 432 348
rect 440 340 462 348
rect 470 340 492 348
rect 500 340 522 348
rect 530 340 552 348
rect 560 340 600 348
rect 0 338 600 340
rect 0 330 32 338
rect 40 330 52 338
rect 60 330 82 338
rect 90 330 112 338
rect 120 330 142 338
rect 150 330 172 338
rect 180 330 202 338
rect 210 330 232 338
rect 240 330 262 338
rect 270 330 292 338
rect 300 330 322 338
rect 330 330 352 338
rect 360 330 382 338
rect 390 330 412 338
rect 420 330 442 338
rect 450 330 472 338
rect 480 330 502 338
rect 510 330 532 338
rect 540 330 562 338
rect 570 330 600 338
rect 0 328 600 330
rect 0 320 42 328
rect 50 320 72 328
rect 80 320 102 328
rect 110 320 132 328
rect 140 320 162 328
rect 170 320 192 328
rect 200 320 222 328
rect 230 320 252 328
rect 260 320 282 328
rect 290 320 312 328
rect 320 320 342 328
rect 350 320 372 328
rect 380 320 402 328
rect 410 320 432 328
rect 440 320 462 328
rect 470 320 492 328
rect 500 320 522 328
rect 530 320 552 328
rect 560 320 600 328
rect 0 318 600 320
rect 0 310 32 318
rect 40 310 52 318
rect 60 310 82 318
rect 90 310 112 318
rect 120 310 142 318
rect 150 310 172 318
rect 180 310 202 318
rect 210 310 232 318
rect 240 310 262 318
rect 270 310 292 318
rect 300 310 322 318
rect 330 310 352 318
rect 360 310 382 318
rect 390 310 412 318
rect 420 310 442 318
rect 450 310 472 318
rect 480 310 502 318
rect 510 310 532 318
rect 540 310 562 318
rect 570 310 600 318
rect 0 308 100 310
rect 0 300 42 308
rect 50 300 72 308
rect 80 300 92 308
rect 500 308 600 310
rect 500 300 522 308
rect 530 300 552 308
rect 560 300 600 308
rect 0 298 600 300
rect 0 290 32 298
rect 40 290 52 298
rect 60 290 82 298
rect 90 290 112 298
rect 120 290 142 298
rect 150 290 172 298
rect 180 290 202 298
rect 210 290 232 298
rect 240 290 262 298
rect 270 290 292 298
rect 300 290 322 298
rect 330 290 352 298
rect 360 290 382 298
rect 390 290 412 298
rect 420 290 442 298
rect 450 290 472 298
rect 480 290 502 298
rect 510 290 532 298
rect 540 290 562 298
rect 570 290 600 298
rect 0 288 600 290
rect 0 280 42 288
rect 50 280 72 288
rect 80 280 102 288
rect 110 280 132 288
rect 140 280 162 288
rect 170 280 192 288
rect 200 280 222 288
rect 230 280 252 288
rect 260 280 282 288
rect 290 280 312 288
rect 320 280 342 288
rect 350 280 372 288
rect 380 280 402 288
rect 410 280 432 288
rect 440 280 462 288
rect 470 280 492 288
rect 500 280 522 288
rect 530 280 552 288
rect 560 280 600 288
rect 0 278 600 280
rect 0 270 32 278
rect 40 270 52 278
rect 60 270 82 278
rect 90 270 112 278
rect 120 270 142 278
rect 150 270 172 278
rect 180 270 202 278
rect 210 270 232 278
rect 240 270 262 278
rect 270 270 292 278
rect 300 270 322 278
rect 330 270 352 278
rect 360 270 382 278
rect 390 270 412 278
rect 420 270 442 278
rect 450 270 472 278
rect 480 270 502 278
rect 510 270 532 278
rect 540 270 562 278
rect 570 270 600 278
rect 0 268 600 270
rect 0 260 42 268
rect 50 260 72 268
rect 80 260 102 268
rect 110 260 132 268
rect 140 260 162 268
rect 170 260 192 268
rect 200 260 222 268
rect 230 260 252 268
rect 260 260 282 268
rect 290 260 312 268
rect 320 260 342 268
rect 350 260 372 268
rect 380 260 402 268
rect 410 260 432 268
rect 440 260 462 268
rect 470 260 492 268
rect 500 260 522 268
rect 530 260 552 268
rect 560 260 600 268
rect 0 258 600 260
rect 0 250 32 258
rect 40 250 52 258
rect 60 250 82 258
rect 90 250 112 258
rect 120 250 142 258
rect 150 250 172 258
rect 180 250 202 258
rect 210 250 232 258
rect 240 250 262 258
rect 270 250 292 258
rect 300 250 322 258
rect 330 250 352 258
rect 360 250 382 258
rect 390 250 412 258
rect 420 250 442 258
rect 450 250 472 258
rect 480 250 502 258
rect 510 250 532 258
rect 540 250 562 258
rect 570 250 600 258
rect 0 248 600 250
rect 0 240 42 248
rect 50 240 72 248
rect 0 238 72 240
rect 0 230 32 238
rect 40 230 52 238
rect 60 230 72 238
rect 0 228 72 230
rect 0 220 42 228
rect 50 220 72 228
rect 80 240 102 248
rect 110 240 132 248
rect 140 240 162 248
rect 170 240 192 248
rect 200 240 222 248
rect 230 240 252 248
rect 260 240 282 248
rect 290 240 312 248
rect 320 240 342 248
rect 350 240 372 248
rect 380 240 402 248
rect 410 240 432 248
rect 440 240 462 248
rect 470 240 492 248
rect 500 240 522 248
rect 530 240 552 248
rect 560 240 600 248
rect 80 238 600 240
rect 80 230 512 238
rect 520 230 532 238
rect 540 230 562 238
rect 570 230 600 238
rect 80 228 600 230
rect 80 220 102 228
rect 110 220 132 228
rect 140 220 162 228
rect 170 220 192 228
rect 200 220 222 228
rect 230 220 252 228
rect 260 220 282 228
rect 290 220 312 228
rect 320 220 342 228
rect 350 220 372 228
rect 380 220 402 228
rect 410 220 432 228
rect 440 220 462 228
rect 470 220 492 228
rect 500 220 522 228
rect 530 220 552 228
rect 560 220 600 228
rect 0 218 600 220
rect 0 210 32 218
rect 40 210 52 218
rect 60 210 82 218
rect 90 210 112 218
rect 120 210 142 218
rect 150 210 172 218
rect 180 210 202 218
rect 210 210 232 218
rect 240 210 262 218
rect 270 210 292 218
rect 300 210 322 218
rect 330 210 352 218
rect 360 210 382 218
rect 390 210 412 218
rect 420 210 442 218
rect 450 210 472 218
rect 480 210 502 218
rect 510 210 532 218
rect 540 210 562 218
rect 570 210 600 218
rect 0 208 600 210
rect 0 200 42 208
rect 50 200 72 208
rect 80 200 102 208
rect 110 200 132 208
rect 140 200 162 208
rect 170 200 192 208
rect 200 200 222 208
rect 230 200 252 208
rect 260 200 282 208
rect 290 200 312 208
rect 320 200 342 208
rect 350 200 372 208
rect 380 200 402 208
rect 410 200 432 208
rect 440 200 462 208
rect 470 200 492 208
rect 500 200 522 208
rect 530 200 552 208
rect 560 200 600 208
rect 0 198 600 200
rect 0 190 32 198
rect 40 190 52 198
rect 60 190 82 198
rect 90 190 112 198
rect 120 190 142 198
rect 150 190 172 198
rect 180 190 202 198
rect 210 190 232 198
rect 240 190 262 198
rect 270 190 292 198
rect 300 190 322 198
rect 330 190 352 198
rect 360 190 382 198
rect 390 190 412 198
rect 420 190 442 198
rect 450 190 472 198
rect 480 190 502 198
rect 510 190 532 198
rect 540 190 562 198
rect 570 190 600 198
rect 0 188 600 190
rect 0 180 42 188
rect 50 180 72 188
rect 80 180 102 188
rect 110 180 132 188
rect 140 180 162 188
rect 170 180 192 188
rect 200 180 222 188
rect 230 180 252 188
rect 260 180 282 188
rect 290 180 312 188
rect 320 180 342 188
rect 350 180 372 188
rect 380 180 402 188
rect 410 180 432 188
rect 440 180 462 188
rect 470 180 492 188
rect 500 180 522 188
rect 530 180 552 188
rect 560 180 600 188
rect 0 178 600 180
rect 0 170 32 178
rect 40 170 52 178
rect 60 170 82 178
rect 90 170 112 178
rect 120 170 142 178
rect 150 170 172 178
rect 180 170 202 178
rect 210 170 232 178
rect 240 170 262 178
rect 270 170 292 178
rect 300 170 322 178
rect 330 170 352 178
rect 360 170 382 178
rect 390 170 412 178
rect 420 170 442 178
rect 450 170 472 178
rect 480 170 502 178
rect 510 170 532 178
rect 540 170 562 178
rect 570 170 600 178
rect 0 168 600 170
rect 0 160 42 168
rect 50 160 72 168
rect 80 160 102 168
rect 110 160 132 168
rect 140 160 162 168
rect 170 160 192 168
rect 200 160 222 168
rect 230 160 252 168
rect 260 160 282 168
rect 290 160 312 168
rect 320 160 342 168
rect 350 160 372 168
rect 380 160 402 168
rect 410 160 432 168
rect 440 160 462 168
rect 470 160 492 168
rect 500 160 522 168
rect 530 160 552 168
rect 560 160 600 168
rect 0 158 100 160
rect 0 150 32 158
rect 40 150 52 158
rect 60 150 82 158
rect 90 150 100 158
rect 500 158 600 160
rect 500 150 512 158
rect 520 150 532 158
rect 540 150 562 158
rect 570 150 600 158
rect 0 148 600 150
rect 0 140 42 148
rect 50 140 72 148
rect 80 140 102 148
rect 110 140 132 148
rect 140 140 162 148
rect 170 140 192 148
rect 200 140 222 148
rect 230 140 252 148
rect 260 140 282 148
rect 290 140 312 148
rect 320 140 342 148
rect 350 140 372 148
rect 380 140 402 148
rect 410 140 432 148
rect 440 140 462 148
rect 470 140 492 148
rect 500 140 522 148
rect 530 140 552 148
rect 560 140 600 148
rect 0 138 600 140
rect 0 130 32 138
rect 40 130 52 138
rect 60 130 82 138
rect 90 130 112 138
rect 120 130 142 138
rect 150 130 172 138
rect 180 130 202 138
rect 210 130 232 138
rect 240 130 262 138
rect 270 130 292 138
rect 300 130 322 138
rect 330 130 352 138
rect 360 130 382 138
rect 390 130 412 138
rect 420 130 442 138
rect 450 130 472 138
rect 480 130 502 138
rect 510 130 532 138
rect 540 130 562 138
rect 570 130 600 138
rect 0 128 600 130
rect 0 120 42 128
rect 50 120 72 128
rect 80 120 102 128
rect 110 120 132 128
rect 140 120 162 128
rect 170 120 192 128
rect 200 120 222 128
rect 230 120 252 128
rect 260 120 282 128
rect 290 120 312 128
rect 320 120 342 128
rect 350 120 372 128
rect 380 120 402 128
rect 410 120 432 128
rect 440 120 462 128
rect 470 120 492 128
rect 500 120 522 128
rect 530 120 552 128
rect 560 120 600 128
rect 0 118 600 120
rect 0 110 32 118
rect 40 110 52 118
rect 60 110 82 118
rect 90 110 112 118
rect 120 110 142 118
rect 150 110 172 118
rect 180 110 202 118
rect 210 110 232 118
rect 240 110 262 118
rect 270 110 292 118
rect 300 110 322 118
rect 330 110 352 118
rect 360 110 382 118
rect 390 110 412 118
rect 420 110 442 118
rect 450 110 472 118
rect 480 110 502 118
rect 510 110 532 118
rect 540 110 562 118
rect 570 110 600 118
rect 0 108 600 110
rect 0 100 42 108
rect 50 100 72 108
rect 80 100 102 108
rect 110 100 132 108
rect 140 100 162 108
rect 170 100 192 108
rect 200 100 222 108
rect 230 100 252 108
rect 260 100 282 108
rect 290 100 312 108
rect 320 100 342 108
rect 350 100 372 108
rect 380 100 402 108
rect 410 100 432 108
rect 440 100 462 108
rect 470 100 492 108
rect 500 100 522 108
rect 530 100 552 108
rect 560 100 600 108
rect 0 98 600 100
rect 0 90 32 98
rect 40 90 52 98
rect 60 90 82 98
rect 90 90 112 98
rect 120 90 142 98
rect 150 90 172 98
rect 180 90 202 98
rect 210 90 232 98
rect 240 90 262 98
rect 270 90 292 98
rect 300 90 322 98
rect 330 90 352 98
rect 360 90 382 98
rect 390 90 412 98
rect 420 90 442 98
rect 450 90 472 98
rect 480 90 502 98
rect 510 90 532 98
rect 540 90 562 98
rect 570 90 600 98
rect 0 88 600 90
rect 0 80 42 88
rect 50 80 72 88
rect 80 80 102 88
rect 110 80 132 88
rect 140 80 162 88
rect 170 80 192 88
rect 200 80 222 88
rect 230 80 252 88
rect 260 80 282 88
rect 290 80 312 88
rect 320 80 342 88
rect 350 80 372 88
rect 380 80 402 88
rect 410 80 432 88
rect 440 80 462 88
rect 470 80 492 88
rect 500 80 522 88
rect 530 80 552 88
rect 560 80 600 88
rect 0 78 600 80
rect 0 70 32 78
rect 40 70 52 78
rect 60 70 82 78
rect 90 70 112 78
rect 120 70 142 78
rect 150 70 172 78
rect 180 70 202 78
rect 210 70 232 78
rect 240 70 262 78
rect 270 70 292 78
rect 300 70 322 78
rect 330 70 352 78
rect 360 70 382 78
rect 390 70 412 78
rect 420 70 442 78
rect 450 70 472 78
rect 480 70 502 78
rect 510 70 532 78
rect 540 70 562 78
rect 570 70 600 78
rect 0 68 600 70
rect 0 60 42 68
rect 50 60 72 68
rect 80 60 102 68
rect 110 60 132 68
rect 140 60 162 68
rect 170 60 192 68
rect 200 60 222 68
rect 230 60 252 68
rect 260 60 282 68
rect 290 60 312 68
rect 320 60 342 68
rect 350 60 372 68
rect 380 60 402 68
rect 410 60 432 68
rect 440 60 462 68
rect 470 60 492 68
rect 500 60 522 68
rect 530 60 552 68
rect 560 60 600 68
rect 0 58 600 60
rect 0 50 32 58
rect 40 50 52 58
rect 60 50 82 58
rect 90 50 112 58
rect 120 50 142 58
rect 150 50 172 58
rect 180 50 202 58
rect 210 50 232 58
rect 240 50 262 58
rect 270 50 292 58
rect 300 50 322 58
rect 330 50 352 58
rect 360 50 382 58
rect 390 50 412 58
rect 420 50 442 58
rect 450 50 472 58
rect 480 50 502 58
rect 510 50 532 58
rect 540 50 562 58
rect 570 50 600 58
rect 0 48 600 50
rect 0 40 42 48
rect 50 40 72 48
rect 80 40 102 48
rect 110 40 132 48
rect 140 40 162 48
rect 170 40 192 48
rect 200 40 222 48
rect 230 40 252 48
rect 260 40 282 48
rect 290 40 312 48
rect 320 40 342 48
rect 350 40 372 48
rect 380 40 402 48
rect 410 40 432 48
rect 440 40 462 48
rect 470 40 492 48
rect 500 40 522 48
rect 530 40 552 48
rect 560 40 600 48
rect 0 38 600 40
rect 0 30 32 38
rect 40 30 52 38
rect 60 30 82 38
rect 90 30 112 38
rect 120 30 142 38
rect 150 30 172 38
rect 180 30 202 38
rect 210 30 232 38
rect 240 30 262 38
rect 270 30 292 38
rect 300 30 322 38
rect 330 30 352 38
rect 360 30 382 38
rect 390 30 412 38
rect 420 30 442 38
rect 450 30 472 38
rect 480 30 502 38
rect 510 30 532 38
rect 540 30 562 38
rect 570 30 600 38
rect 0 0 600 30
use PadBox  PadBox_0
timestamp 1570494029
transform 1 0 40 0 1 1480
box 0 0 520 520
<< labels >>
flabel nwell 600 -6 600 -6 6 FreeSans 16 0 0 0 VddNW
flabel nwell 0 -6 0 -6 4 FreeSans 16 0 0 0 VddNW
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 VddAct
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 VddAct
flabel psubstratepdiff 0 686 0 686 4 FreeSans 16 0 0 0 GndAct
flabel psubstratepdiff 600 686 600 686 6 FreeSans 16 0 0 0 GndAct
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 688 600 688 6 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 688 0 688 4 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 880 0 880 4 FreeSans 16 0 0 0 VddM2A
flabel metal2 600 880 600 880 6 FreeSans 16 0 0 0 VddM2A
flabel metal2 0 492 0 492 4 FreeSans 16 0 0 0 VddM2B
flabel metal2 600 492 600 492 6 FreeSans 16 0 0 0 VddM2B
<< properties >>
string path 0.000 1035.000 225.000 1035.000 225.000 337.500 1125.000 337.500 1125.000 360.000 225.000 360.000 225.000 675.000 1125.000 675.000 1125.000 697.500 225.000 697.500 225.000 1035.000 1350.000 1035.000 1350.000 0.000 0.000 0.000 0.000 1035.000 
<< end >>
