magic
tech amic5n
timestamp 1623365459
<< nwell >>
rect -130 550 3285 1495
<< ntransistor >>
rect 165 95 225 375
rect 355 95 415 375
rect 545 95 605 375
rect 695 95 755 375
rect 965 95 1025 375
rect 1115 95 1175 375
rect 1310 95 1370 375
rect 1950 95 2010 375
rect 2100 95 2160 375
rect 2370 95 2430 375
rect 2520 95 2580 375
rect 2735 95 2795 375
rect 2925 95 2985 375
<< ptransistor >>
rect 165 865 225 1345
rect 355 865 415 1345
rect 545 865 605 1345
rect 725 865 785 1345
rect 965 865 1025 1345
rect 1115 865 1175 1345
rect 1310 865 1370 1345
rect 1950 865 2010 1345
rect 2100 865 2160 1345
rect 2370 1065 2430 1345
rect 2520 1065 2580 1345
rect 2735 865 2795 1345
rect 2925 865 2985 1345
<< nselect >>
rect 1650 835 1830 1240
rect -10 165 1650 430
rect 1830 165 3160 430
rect -10 0 3160 165
<< pselect >>
rect 2570 1440 2805 1445
rect -10 1240 3160 1440
rect -10 835 1650 1240
rect 1830 835 3160 1240
rect 1650 165 1830 430
<< ndiffusion >>
rect 45 345 165 375
rect 45 295 75 345
rect 125 295 165 345
rect 45 175 165 295
rect 45 125 75 175
rect 125 125 165 175
rect 45 95 165 125
rect 225 345 355 375
rect 225 295 265 345
rect 315 295 355 345
rect 225 175 355 295
rect 225 125 265 175
rect 315 125 355 175
rect 225 95 355 125
rect 415 345 545 375
rect 415 295 455 345
rect 505 295 545 345
rect 415 175 545 295
rect 415 125 455 175
rect 505 125 545 175
rect 415 95 545 125
rect 605 95 695 375
rect 755 345 965 375
rect 755 295 850 345
rect 900 295 965 345
rect 755 200 965 295
rect 755 150 850 200
rect 900 150 965 200
rect 755 95 965 150
rect 1025 95 1115 375
rect 1175 345 1310 375
rect 1175 295 1220 345
rect 1270 295 1310 345
rect 1175 175 1310 295
rect 1175 125 1220 175
rect 1270 125 1310 175
rect 1175 95 1310 125
rect 1370 345 1490 375
rect 1370 295 1410 345
rect 1460 295 1490 345
rect 1370 175 1490 295
rect 1370 125 1410 175
rect 1460 125 1490 175
rect 1830 345 1950 375
rect 1830 295 1860 345
rect 1910 295 1950 345
rect 1830 175 1950 295
rect 1370 95 1490 125
rect 1830 125 1860 175
rect 1910 125 1950 175
rect 1830 95 1950 125
rect 2010 95 2100 375
rect 2160 345 2370 375
rect 2160 295 2240 345
rect 2290 295 2370 345
rect 2160 175 2370 295
rect 2160 125 2240 175
rect 2290 125 2370 175
rect 2160 95 2370 125
rect 2430 95 2520 375
rect 2580 345 2735 375
rect 2580 295 2635 345
rect 2685 295 2735 345
rect 2580 175 2735 295
rect 2580 125 2635 175
rect 2685 125 2735 175
rect 2580 95 2735 125
rect 2795 345 2925 375
rect 2795 295 2835 345
rect 2885 295 2925 345
rect 2795 175 2925 295
rect 2795 125 2835 175
rect 2885 125 2925 175
rect 2795 95 2925 125
rect 2985 345 3105 375
rect 2985 295 3025 345
rect 3075 295 3105 345
rect 2985 175 3105 295
rect 2985 125 3025 175
rect 3075 125 3105 175
rect 2985 95 3105 125
<< pdiffusion >>
rect 45 1315 165 1345
rect 45 1265 75 1315
rect 125 1265 165 1315
rect 45 1195 165 1265
rect 45 1145 75 1195
rect 125 1145 165 1195
rect 45 1070 165 1145
rect 45 1020 75 1070
rect 125 1020 165 1070
rect 45 945 165 1020
rect 45 895 75 945
rect 125 895 165 945
rect 45 865 165 895
rect 225 1315 355 1345
rect 225 1265 265 1315
rect 315 1265 355 1315
rect 225 1195 355 1265
rect 225 1145 265 1195
rect 315 1145 355 1195
rect 225 1070 355 1145
rect 225 1020 265 1070
rect 315 1020 355 1070
rect 225 945 355 1020
rect 225 895 265 945
rect 315 895 355 945
rect 225 865 355 895
rect 415 1315 545 1345
rect 415 1265 455 1315
rect 505 1265 545 1315
rect 415 1200 545 1265
rect 415 1150 455 1200
rect 505 1150 545 1200
rect 415 1085 545 1150
rect 415 1035 455 1085
rect 505 1035 545 1085
rect 415 975 545 1035
rect 415 925 455 975
rect 505 925 545 975
rect 415 865 545 925
rect 605 865 725 1345
rect 785 1315 965 1345
rect 785 1265 845 1315
rect 895 1265 965 1315
rect 785 1195 965 1265
rect 785 1145 845 1195
rect 895 1145 965 1195
rect 785 1080 965 1145
rect 785 1030 845 1080
rect 895 1030 965 1080
rect 785 945 965 1030
rect 785 895 845 945
rect 895 895 965 945
rect 785 865 965 895
rect 1025 865 1115 1345
rect 1175 1315 1310 1345
rect 1175 1265 1220 1315
rect 1270 1265 1310 1315
rect 1175 1200 1310 1265
rect 1175 1150 1220 1200
rect 1270 1150 1310 1200
rect 1175 1085 1310 1150
rect 1175 1035 1220 1085
rect 1270 1035 1310 1085
rect 1175 975 1310 1035
rect 1175 925 1220 975
rect 1270 925 1310 975
rect 1175 865 1310 925
rect 1370 1315 1490 1345
rect 1370 1265 1410 1315
rect 1460 1265 1490 1315
rect 1370 1195 1490 1265
rect 1830 1315 1950 1345
rect 1830 1265 1860 1315
rect 1910 1265 1950 1315
rect 1370 1145 1410 1195
rect 1460 1145 1490 1195
rect 1370 1070 1490 1145
rect 1370 1020 1410 1070
rect 1460 1020 1490 1070
rect 1370 945 1490 1020
rect 1370 895 1410 945
rect 1460 895 1490 945
rect 1370 865 1490 895
rect 1830 1200 1950 1265
rect 1830 1150 1860 1200
rect 1910 1150 1950 1200
rect 1830 1085 1950 1150
rect 1830 1035 1860 1085
rect 1910 1035 1950 1085
rect 1830 975 1950 1035
rect 1830 925 1860 975
rect 1910 925 1950 975
rect 1830 865 1950 925
rect 2010 865 2100 1345
rect 2160 1315 2370 1345
rect 2160 1265 2240 1315
rect 2290 1265 2370 1315
rect 2160 1195 2370 1265
rect 2160 1145 2240 1195
rect 2290 1145 2370 1195
rect 2160 1070 2370 1145
rect 2160 1020 2240 1070
rect 2290 1065 2370 1070
rect 2430 1065 2520 1345
rect 2580 1315 2735 1345
rect 2580 1265 2630 1315
rect 2680 1265 2735 1315
rect 2580 1145 2735 1265
rect 2580 1095 2630 1145
rect 2680 1095 2735 1145
rect 2580 1065 2735 1095
rect 2290 1020 2340 1065
rect 2160 945 2340 1020
rect 2160 895 2240 945
rect 2290 895 2340 945
rect 2160 865 2340 895
rect 2670 865 2735 1065
rect 2795 1315 2925 1345
rect 2795 1265 2835 1315
rect 2885 1265 2925 1315
rect 2795 1195 2925 1265
rect 2795 1145 2835 1195
rect 2885 1145 2925 1195
rect 2795 1070 2925 1145
rect 2795 1020 2835 1070
rect 2885 1020 2925 1070
rect 2795 945 2925 1020
rect 2795 895 2835 945
rect 2885 895 2925 945
rect 2795 865 2925 895
rect 2985 1315 3105 1345
rect 2985 1265 3025 1315
rect 3075 1265 3105 1315
rect 2985 1195 3105 1265
rect 2985 1145 3025 1195
rect 3075 1145 3105 1195
rect 2985 1070 3105 1145
rect 2985 1020 3025 1070
rect 3075 1020 3105 1070
rect 2985 945 3105 1020
rect 2985 895 3025 945
rect 3075 895 3105 945
rect 2985 865 3105 895
<< psubstratepdiff >>
rect 1720 345 1830 375
rect 1720 295 1750 345
rect 1800 295 1830 345
rect 1720 245 1830 295
rect 1720 195 1750 245
rect 1800 195 1830 245
rect 1720 165 1830 195
<< nsubstratendiff >>
rect 1710 1175 1830 1240
rect 1710 1125 1745 1175
rect 1795 1125 1830 1175
rect 1710 1075 1830 1125
rect 1710 1025 1745 1075
rect 1795 1025 1830 1075
rect 1710 975 1830 1025
rect 1710 925 1745 975
rect 1795 925 1830 975
rect 1710 865 1830 925
<< nsubstratencontact >>
rect 1745 1125 1795 1175
rect 1745 1025 1795 1075
rect 1745 925 1795 975
<< psubstratepcontact >>
rect 1750 295 1800 345
rect 1750 195 1800 245
<< ndcontact >>
rect 75 295 125 345
rect 75 125 125 175
rect 265 295 315 345
rect 265 125 315 175
rect 455 295 505 345
rect 455 125 505 175
rect 850 295 900 345
rect 850 150 900 200
rect 1220 295 1270 345
rect 1220 125 1270 175
rect 1410 295 1460 345
rect 1410 125 1460 175
rect 1860 295 1910 345
rect 1860 125 1910 175
rect 2240 295 2290 345
rect 2240 125 2290 175
rect 2635 295 2685 345
rect 2635 125 2685 175
rect 2835 295 2885 345
rect 2835 125 2885 175
rect 3025 295 3075 345
rect 3025 125 3075 175
<< pdcontact >>
rect 75 1265 125 1315
rect 75 1145 125 1195
rect 75 1020 125 1070
rect 75 895 125 945
rect 265 1265 315 1315
rect 265 1145 315 1195
rect 265 1020 315 1070
rect 265 895 315 945
rect 455 1265 505 1315
rect 455 1150 505 1200
rect 455 1035 505 1085
rect 455 925 505 975
rect 845 1265 895 1315
rect 845 1145 895 1195
rect 845 1030 895 1080
rect 845 895 895 945
rect 1220 1265 1270 1315
rect 1220 1150 1270 1200
rect 1220 1035 1270 1085
rect 1220 925 1270 975
rect 1410 1265 1460 1315
rect 1860 1265 1910 1315
rect 1410 1145 1460 1195
rect 1410 1020 1460 1070
rect 1410 895 1460 945
rect 1860 1150 1910 1200
rect 1860 1035 1910 1085
rect 1860 925 1910 975
rect 2240 1265 2290 1315
rect 2240 1145 2290 1195
rect 2240 1020 2290 1070
rect 2630 1265 2680 1315
rect 2630 1095 2680 1145
rect 2240 895 2290 945
rect 2835 1265 2885 1315
rect 2835 1145 2885 1195
rect 2835 1020 2885 1070
rect 2835 895 2885 945
rect 3025 1265 3075 1315
rect 3025 1145 3075 1195
rect 3025 1020 3075 1070
rect 3025 895 3075 945
<< polysilicon >>
rect 165 1345 225 1410
rect 355 1345 415 1410
rect 545 1345 605 1410
rect 725 1345 785 1410
rect 965 1345 1025 1410
rect 1115 1345 1175 1410
rect 1310 1345 1370 1410
rect 1950 1345 2010 1410
rect 2100 1345 2160 1410
rect 2370 1345 2430 1410
rect 2520 1345 2580 1410
rect 2735 1345 2795 1410
rect 2925 1345 2985 1410
rect 165 845 225 865
rect 355 845 415 865
rect 545 845 605 865
rect 725 845 785 865
rect 165 785 415 845
rect 515 825 605 845
rect 165 525 225 785
rect 515 775 535 825
rect 585 775 605 825
rect 515 755 605 775
rect 665 825 785 845
rect 665 775 685 825
rect 735 775 785 825
rect 665 755 785 775
rect 165 505 485 525
rect 165 455 415 505
rect 465 455 485 505
rect 165 435 485 455
rect 165 375 225 435
rect 355 375 415 435
rect 545 375 605 755
rect 965 685 1025 865
rect 950 665 1040 685
rect 950 655 970 665
rect 695 615 970 655
rect 1020 615 1040 665
rect 695 595 1040 615
rect 695 375 755 595
rect 1115 525 1175 865
rect 1310 845 1370 865
rect 1950 845 2010 865
rect 1235 825 1370 845
rect 1235 775 1255 825
rect 1305 775 1370 825
rect 1235 755 1370 775
rect 1905 825 2010 845
rect 1905 775 1925 825
rect 1975 775 2010 825
rect 1905 755 2010 775
rect 950 505 1040 525
rect 950 455 970 505
rect 1020 455 1040 505
rect 950 435 1040 455
rect 1100 505 1190 525
rect 1100 455 1120 505
rect 1170 455 1190 505
rect 1100 435 1190 455
rect 965 375 1025 435
rect 1115 375 1175 435
rect 1310 375 1370 755
rect 1950 375 2010 755
rect 2100 685 2160 865
rect 2070 665 2160 685
rect 2070 615 2090 665
rect 2140 655 2160 665
rect 2370 685 2430 1065
rect 2370 665 2460 685
rect 2140 615 2295 655
rect 2070 595 2295 615
rect 2370 615 2390 665
rect 2440 615 2460 665
rect 2370 595 2460 615
rect 2070 505 2160 525
rect 2070 455 2090 505
rect 2140 455 2160 505
rect 2070 435 2160 455
rect 2100 375 2160 435
rect 2235 455 2295 595
rect 2520 525 2580 1065
rect 2735 845 2795 865
rect 2925 845 2985 865
rect 2665 825 2985 845
rect 2665 775 2685 825
rect 2735 785 2985 825
rect 2735 775 2795 785
rect 2665 755 2795 775
rect 2520 505 2625 525
rect 2520 455 2555 505
rect 2605 455 2625 505
rect 2235 395 2430 455
rect 2370 375 2430 395
rect 2520 435 2625 455
rect 2735 455 2795 755
rect 2520 375 2580 435
rect 2735 395 2985 455
rect 2735 375 2795 395
rect 2925 375 2985 395
rect 165 30 225 95
rect 355 30 415 95
rect 545 30 605 95
rect 695 30 755 95
rect 965 30 1025 95
rect 1115 30 1175 95
rect 1310 30 1370 95
rect 1950 30 2010 95
rect 2100 30 2160 95
rect 2370 30 2430 95
rect 2520 30 2580 95
rect 2735 30 2795 95
rect 2925 30 2985 95
<< polycontact >>
rect 535 775 585 825
rect 685 775 735 825
rect 415 455 465 505
rect 970 615 1020 665
rect 1255 775 1305 825
rect 1925 775 1975 825
rect 970 455 1020 505
rect 1120 455 1170 505
rect 2090 615 2140 665
rect 2390 615 2440 665
rect 2090 455 2140 505
rect 2685 775 2735 825
rect 2555 455 2605 505
<< metal1 >>
rect 0 1395 3150 1485
rect 55 1315 145 1395
rect 55 1265 75 1315
rect 125 1265 145 1315
rect 55 1195 145 1265
rect 55 1145 75 1195
rect 125 1145 145 1195
rect 55 1070 145 1145
rect 55 1020 75 1070
rect 125 1020 145 1070
rect 55 945 145 1020
rect 55 895 75 945
rect 125 895 145 945
rect 55 875 145 895
rect 245 1315 335 1335
rect 245 1265 265 1315
rect 315 1265 335 1315
rect 245 1195 335 1265
rect 245 1145 265 1195
rect 315 1145 335 1195
rect 245 1070 335 1145
rect 245 1020 265 1070
rect 315 1020 335 1070
rect 245 945 335 1020
rect 245 895 265 945
rect 315 895 335 945
rect 435 1315 525 1395
rect 435 1265 455 1315
rect 505 1265 525 1315
rect 435 1200 525 1265
rect 435 1150 455 1200
rect 505 1150 525 1200
rect 435 1085 525 1150
rect 435 1035 455 1085
rect 505 1035 525 1085
rect 435 975 525 1035
rect 435 925 455 975
rect 505 925 525 975
rect 435 905 525 925
rect 815 1315 920 1335
rect 815 1265 845 1315
rect 895 1265 920 1315
rect 815 1195 920 1265
rect 815 1145 845 1195
rect 895 1145 920 1195
rect 815 1080 920 1145
rect 815 1030 845 1080
rect 895 1030 920 1080
rect 815 945 920 1030
rect 245 685 335 895
rect 815 895 845 945
rect 895 895 920 945
rect 1200 1315 1290 1395
rect 1200 1265 1220 1315
rect 1270 1265 1290 1315
rect 1200 1200 1290 1265
rect 1200 1150 1220 1200
rect 1270 1150 1290 1200
rect 1200 1085 1290 1150
rect 1200 1035 1220 1085
rect 1270 1035 1290 1085
rect 1200 975 1290 1035
rect 1200 925 1220 975
rect 1270 925 1290 975
rect 1200 905 1290 925
rect 1390 1315 1480 1335
rect 1390 1265 1410 1315
rect 1460 1265 1480 1315
rect 1390 1195 1480 1265
rect 1390 1145 1410 1195
rect 1460 1145 1480 1195
rect 1390 1070 1480 1145
rect 1390 1020 1410 1070
rect 1460 1020 1480 1070
rect 1390 945 1480 1020
rect 815 845 920 895
rect 1390 895 1410 945
rect 1460 895 1480 945
rect 1725 1315 1930 1395
rect 1725 1265 1860 1315
rect 1910 1265 1930 1315
rect 1725 1200 1930 1265
rect 1725 1175 1860 1200
rect 1725 1125 1745 1175
rect 1795 1150 1860 1175
rect 1910 1150 1930 1200
rect 1795 1125 1930 1150
rect 1725 1085 1930 1125
rect 1725 1075 1860 1085
rect 1725 1025 1745 1075
rect 1795 1035 1860 1075
rect 1910 1035 1930 1085
rect 1795 1025 1930 1035
rect 1725 975 1930 1025
rect 1725 925 1745 975
rect 1795 925 1860 975
rect 1910 925 1930 975
rect 1725 905 1930 925
rect 2220 1315 2310 1335
rect 2220 1265 2240 1315
rect 2290 1265 2310 1315
rect 2220 1195 2310 1265
rect 2220 1145 2240 1195
rect 2290 1145 2310 1195
rect 2220 1070 2310 1145
rect 2610 1315 2700 1395
rect 2610 1265 2630 1315
rect 2680 1265 2700 1315
rect 2610 1145 2700 1265
rect 2610 1095 2630 1145
rect 2680 1095 2700 1145
rect 2610 1075 2700 1095
rect 2815 1315 2905 1335
rect 2815 1265 2835 1315
rect 2885 1265 2905 1315
rect 2815 1195 2905 1265
rect 2815 1145 2835 1195
rect 2885 1145 2905 1195
rect 2220 1020 2240 1070
rect 2290 1020 2310 1070
rect 2220 945 2310 1020
rect 1390 845 1480 895
rect 2220 895 2240 945
rect 2290 895 2310 945
rect 2220 845 2310 895
rect 2815 1070 2905 1145
rect 2815 1020 2835 1070
rect 2885 1020 2905 1070
rect 2815 945 2905 1020
rect 2815 895 2835 945
rect 2885 895 2905 945
rect 405 825 605 845
rect 405 775 535 825
rect 585 775 605 825
rect 405 755 605 775
rect 665 825 755 845
rect 665 775 685 825
rect 735 775 755 825
rect 245 665 445 685
rect 245 615 265 665
rect 315 615 375 665
rect 425 615 445 665
rect 245 595 445 615
rect 55 345 145 365
rect 55 295 75 345
rect 125 295 145 345
rect 55 175 145 295
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 245 345 335 595
rect 665 525 755 775
rect 395 505 755 525
rect 395 455 415 505
rect 465 455 545 505
rect 595 455 685 505
rect 735 455 755 505
rect 395 435 755 455
rect 815 825 1325 845
rect 815 775 1255 825
rect 1305 775 1325 825
rect 815 755 1325 775
rect 1390 825 1995 845
rect 1390 775 1925 825
rect 1975 775 1995 825
rect 1390 755 1995 775
rect 2220 825 2755 845
rect 2220 775 2685 825
rect 2735 775 2755 825
rect 2220 755 2755 775
rect 815 365 890 755
rect 950 665 1150 685
rect 950 615 970 665
rect 1020 615 1080 665
rect 1130 615 1150 665
rect 950 595 1150 615
rect 1390 525 1480 755
rect 1960 665 2160 685
rect 1960 615 1980 665
rect 2030 615 2090 665
rect 2140 615 2160 665
rect 1960 595 2160 615
rect 950 505 1040 525
rect 950 455 970 505
rect 1020 455 1040 505
rect 950 435 1040 455
rect 1100 505 1480 525
rect 1100 455 1120 505
rect 1170 455 1480 505
rect 1100 435 1480 455
rect 1960 505 2160 525
rect 1960 455 1980 505
rect 2030 455 2090 505
rect 2140 455 2160 505
rect 1960 435 2160 455
rect 245 295 265 345
rect 315 295 335 345
rect 245 175 335 295
rect 245 125 265 175
rect 315 125 335 175
rect 245 105 335 125
rect 435 345 525 365
rect 435 295 455 345
rect 505 295 525 345
rect 435 175 525 295
rect 435 125 455 175
rect 505 125 525 175
rect 435 45 525 125
rect 815 345 935 365
rect 815 295 850 345
rect 900 295 935 345
rect 815 200 935 295
rect 815 150 850 200
rect 900 150 935 200
rect 815 105 935 150
rect 1200 345 1290 365
rect 1200 295 1220 345
rect 1270 295 1290 345
rect 1200 175 1290 295
rect 1200 125 1220 175
rect 1270 125 1290 175
rect 1200 45 1290 125
rect 1390 345 1480 435
rect 1390 295 1410 345
rect 1460 295 1480 345
rect 1390 175 1480 295
rect 1390 125 1410 175
rect 1460 125 1480 175
rect 1390 105 1480 125
rect 1730 345 1930 365
rect 1730 295 1750 345
rect 1800 295 1860 345
rect 1910 295 1930 345
rect 1730 245 1930 295
rect 1730 195 1750 245
rect 1800 195 1930 245
rect 1730 175 1930 195
rect 1730 125 1860 175
rect 1910 125 1930 175
rect 1730 45 1930 125
rect 2220 345 2310 755
rect 2370 665 2460 685
rect 2370 615 2390 665
rect 2440 615 2460 665
rect 2370 505 2460 615
rect 2815 525 2905 895
rect 3005 1315 3095 1395
rect 3005 1265 3025 1315
rect 3075 1265 3095 1315
rect 3005 1195 3095 1265
rect 3005 1145 3025 1195
rect 3075 1145 3095 1195
rect 3005 1070 3095 1145
rect 3005 1020 3025 1070
rect 3075 1020 3095 1070
rect 3005 945 3095 1020
rect 3005 895 3025 945
rect 3075 895 3095 945
rect 3005 875 3095 895
rect 2370 455 2390 505
rect 2440 455 2460 505
rect 2370 435 2460 455
rect 2520 505 2905 525
rect 2520 455 2555 505
rect 2605 455 2905 505
rect 2520 435 2905 455
rect 2220 295 2240 345
rect 2290 295 2310 345
rect 2220 175 2310 295
rect 2220 125 2240 175
rect 2290 125 2310 175
rect 2220 105 2310 125
rect 2615 345 2705 365
rect 2615 295 2635 345
rect 2685 295 2705 345
rect 2615 175 2705 295
rect 2615 125 2635 175
rect 2685 125 2705 175
rect 2615 45 2705 125
rect 2815 345 2905 435
rect 2815 295 2835 345
rect 2885 295 2905 345
rect 2815 175 2905 295
rect 2815 125 2835 175
rect 2885 125 2905 175
rect 2815 105 2905 125
rect 3005 345 3095 365
rect 3005 295 3025 345
rect 3075 295 3095 345
rect 3005 175 3095 295
rect 3005 125 3025 175
rect 3075 125 3095 175
rect 3005 45 3095 125
rect 0 -45 3150 45
<< via1 >>
rect 265 615 315 665
rect 375 615 425 665
rect 415 455 465 505
rect 545 455 595 505
rect 685 455 735 505
rect 970 615 1020 665
rect 1080 615 1130 665
rect 1980 615 2030 665
rect 2090 615 2140 665
rect 970 455 1020 505
rect 1980 455 2030 505
rect 2090 455 2140 505
rect 2390 455 2440 505
<< metal2 >>
rect 245 665 2220 685
rect 245 615 265 665
rect 315 615 375 665
rect 425 615 970 665
rect 1020 615 1080 665
rect 1130 615 1980 665
rect 2030 615 2090 665
rect 2140 615 2220 665
rect 245 595 2220 615
rect 395 505 2545 525
rect 395 455 415 505
rect 465 455 545 505
rect 595 455 685 505
rect 735 455 970 505
rect 1020 455 1980 505
rect 2030 455 2090 505
rect 2140 455 2390 505
rect 2440 455 2545 505
rect 395 435 2545 455
<< labels >>
flabel ndiffusion s 1055 195 1055 195 2 FreeSans 400 0 0 0 x6
flabel ndiffusion 635 195 635 195 2 FreeSans 400 0 0 0 x5
flabel metal1 s 845 165 845 165 2 FreeSans 400 0 0 0 nmas
flabel metal1 s 225 -15 225 -15 2 FreeSans 400 0 0 0 vss
port 5 s
flabel metal1 260 610 260 610 2 FreeSans 400 0 0 0 nck
flabel metal1 s 415 800 415 800 2 FreeSans 400 0 0 0 d
port 2 s
flabel metal1 s 455 1395 455 1395 2 FreeSans 400 0 0 0 vdd
port 4 n
flabel pdiffusion s 1055 1065 1055 1065 2 FreeSans 400 0 0 0 x2
flabel pdiffusion s 665 1065 665 1065 2 FreeSans 400 0 0 0 x1
flabel metal1 s 1115 770 1115 770 2 FreeSans 400 0 0 0 nmas
flabel metal1 s 1405 285 1405 285 2 FreeSans 400 0 0 0 mas
flabel metal1 s 1420 1065 1420 1065 2 FreeSans 400 0 0 0 mas
flabel metal1 s 950 465 950 465 2 FreeSans 400 0 0 0 ck
port 3 ne
flabel metal1 s 845 925 845 925 2 FreeSans 400 0 0 0 nmas
flabel pdiffusion s 2040 1065 2040 1065 2 FreeSans 400 0 0 0 x3
flabel ndiffusion s 2040 165 2040 165 2 FreeSans 400 0 0 0 x7
flabel nwell s 1770 600 1770 600 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 2085 610 2085 610 2 FreeSans 400 0 0 0 nck
flabel ndiffusion s 2460 165 2460 165 2 FreeSans 400 0 0 0 x8
flabel pdiffusion s 2460 1185 2460 1185 2 FreeSans 400 0 0 0 x4
flabel metal1 s 2835 710 2835 710 2 FreeSans 400 0 0 0 q
port 1 e
flabel metal1 s 2490 800 2490 800 2 FreeSans 400 0 0 0 nslv
<< end >>
