`celldefine
module inv_a (z, a);
  output z;
  input  a;

  not G1 (z, a);
endmodule
`endcelldefine
