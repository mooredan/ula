magic
tech scmos
timestamp 1511331171
<< error_p >>
rect 114 69 123 70
rect 257 54 261 55
rect 258 53 260 54
rect 8 42 16 43
rect 17 42 21 43
rect 22 42 24 48
rect 9 39 10 42
rect 15 39 16 42
rect 18 39 19 42
rect 21 39 24 42
rect 274 43 278 44
rect 274 41 275 43
rect 277 41 278 43
rect 274 40 278 41
rect 8 36 9 37
rect 9 30 10 36
rect 15 30 16 37
rect 17 36 18 37
rect 22 36 24 39
rect 258 37 260 38
rect 18 30 19 36
rect 21 30 24 36
rect 114 33 123 34
rect 258 33 260 34
rect 22 29 24 30
rect 7 27 24 29
rect 114 27 118 28
rect 212 27 215 29
rect 211 22 215 23
rect 211 20 212 22
rect 214 20 215 22
rect 211 19 215 20
rect 211 17 215 18
rect 206 16 210 17
rect 27 15 30 16
rect 3 12 7 13
rect 17 12 21 13
rect 30 12 31 15
rect 206 14 207 16
rect 209 14 210 16
rect 211 15 212 17
rect 214 15 215 17
rect 211 14 215 15
rect 255 15 256 16
rect 255 14 257 15
rect 206 13 210 14
rect 32 12 39 13
rect 6 9 7 12
rect 8 9 16 10
rect 18 9 19 12
rect 33 9 34 12
rect 205 10 209 11
rect 9 6 10 9
rect 15 6 16 9
rect 205 8 206 10
rect 208 8 209 10
rect 205 7 209 8
rect 212 10 216 11
rect 212 8 213 10
rect 215 8 216 10
rect 212 7 216 8
<< nwell >>
rect -3 24 27 54
rect 82 27 139 75
rect 146 27 205 65
rect 218 24 242 65
<< ntransistor >>
rect 6 6 9 15
rect 15 6 18 15
rect 30 6 33 15
rect 106 3 109 22
rect 171 4 173 21
rect 229 4 231 17
<< ptransistor >>
rect 6 27 9 48
rect 15 27 18 48
rect 105 33 108 70
rect 114 33 117 70
rect 170 33 172 59
rect 179 33 181 59
rect 229 30 231 59
<< ndiffusion >>
rect 0 12 6 15
rect 0 9 3 12
rect 0 6 6 9
rect 9 9 15 15
rect 18 12 27 15
rect 21 9 30 12
rect 18 6 30 9
rect 33 12 39 15
rect 33 6 39 9
rect 102 3 106 22
rect 109 3 112 22
rect 167 4 171 21
rect 173 4 177 21
rect 224 4 229 17
rect 231 4 236 17
rect 193 -13 197 -6
rect 200 -13 204 -6
<< pdiffusion >>
rect 0 42 6 48
rect 0 39 3 42
rect 0 36 6 39
rect 0 30 3 36
rect 0 27 6 30
rect 9 42 15 48
rect 9 36 15 39
rect 9 27 15 30
rect 18 42 24 48
rect 21 39 24 42
rect 18 36 24 39
rect 21 30 24 36
rect 99 33 105 70
rect 108 33 114 70
rect 117 33 123 70
rect 164 33 170 59
rect 172 33 179 59
rect 181 33 188 59
rect 211 47 215 51
rect 211 39 215 43
rect 211 31 215 35
rect 18 27 24 30
rect 224 30 229 59
rect 231 30 236 59
rect 254 25 264 56
rect 268 45 273 55
<< ndcontact >>
rect 3 9 6 12
rect 9 6 15 9
rect 27 12 30 15
rect 18 9 21 12
rect 33 9 39 12
<< pdcontact >>
rect 3 39 6 42
rect 3 30 6 36
rect 9 39 15 42
rect 9 30 15 36
rect 18 39 21 42
rect 18 30 21 36
rect 211 51 215 55
rect 211 43 215 47
rect 211 35 215 39
rect 211 27 215 31
<< polysilicon >>
rect 105 70 108 72
rect 114 70 117 72
rect 6 48 9 51
rect 15 48 18 51
rect 170 59 172 61
rect 179 59 181 61
rect 229 59 231 61
rect 105 31 108 33
rect 114 31 117 33
rect 170 31 172 33
rect 179 31 181 33
rect 229 27 231 30
rect 6 24 9 27
rect 15 24 18 27
rect 106 22 109 27
rect 6 15 9 18
rect 15 15 18 18
rect 30 15 33 18
rect 6 3 9 6
rect 15 3 18 6
rect 30 3 33 6
rect 171 21 173 27
rect 224 21 231 27
rect 229 17 231 21
rect 253 12 259 18
rect 106 1 109 3
rect 171 2 173 4
rect 229 2 231 4
rect 171 -13 173 -4
rect 176 -13 178 -4
<< polycontact >>
rect 3 24 6 27
<< genericcontact >>
rect 225 55 227 57
rect 233 54 235 56
rect 258 52 260 54
rect 225 49 227 51
rect 233 48 235 50
rect 258 47 260 49
rect 225 43 227 45
rect 233 43 235 45
rect 258 42 260 44
rect 275 41 277 43
rect 225 37 227 39
rect 233 38 235 40
rect 258 37 260 39
rect 225 32 227 34
rect 233 32 235 34
rect 258 33 260 35
rect 258 29 260 31
rect 226 23 228 25
rect 212 20 214 22
rect 207 14 209 16
rect 212 15 214 17
rect 225 13 227 15
rect 233 13 235 15
rect 255 14 257 16
rect 206 8 208 10
rect 213 8 215 10
rect 225 6 227 8
rect 233 7 235 9
<< metal1 >>
rect 85 70 136 73
rect 85 63 102 66
rect 122 63 136 66
rect 150 60 201 63
rect 222 60 238 63
rect 85 56 99 59
rect 122 56 136 59
rect 150 54 167 57
rect 187 54 201 57
rect 85 49 99 52
rect 122 49 136 52
rect 150 48 164 51
rect 187 48 201 51
rect -3 45 21 48
rect 211 47 215 51
rect 3 42 6 45
rect 18 42 21 45
rect 85 42 136 45
rect 150 42 164 45
rect 187 42 201 45
rect 3 36 6 39
rect 9 36 15 39
rect 211 39 215 43
rect 18 36 21 39
rect 85 35 136 38
rect 150 36 201 39
rect 9 24 15 30
rect 85 28 95 31
rect 126 28 136 31
rect 150 30 201 33
rect 211 31 215 35
rect 224 31 228 60
rect 150 24 160 27
rect 191 24 201 27
rect 85 21 102 24
rect 116 21 136 24
rect 225 22 229 26
rect 150 18 167 21
rect 181 18 201 21
rect 3 12 21 15
rect 85 14 136 17
rect 150 12 201 15
rect 18 6 39 9
rect 85 7 136 10
rect 150 6 201 9
rect 9 3 15 6
rect 224 3 228 16
rect 232 6 236 57
rect 257 26 261 54
rect 254 7 258 19
rect -3 0 39 3
rect 85 0 136 3
rect 150 0 201 3
rect 222 0 238 3
<< metal2 >>
rect 48 70 66 73
rect 48 63 66 66
rect 48 56 66 59
rect 48 49 66 52
rect 48 42 66 45
rect 48 35 66 38
rect 48 28 66 31
rect 27 24 36 27
rect 48 21 66 24
rect 48 14 66 17
rect 248 13 275 17
rect 48 7 66 10
rect 48 0 66 3
<< gv1 >>
rect 255 14 257 16
<< bb >>
rect 0 0 39 51
rect 85 0 136 73
rect 222 0 238 63
<< labels >>
rlabel metal1 -3 0 -3 0 2 Gnd
port 3 ne
rlabel polycontact 3 24 3 24 2 a
port 1 ne
rlabel metal1 -3 45 -3 45 2 Vdd
port 2 ne
rlabel nwell 0 24 0 24 2 Vdd
rlabel metal1 12 30 12 30 2 z
port 0 ne
rlabel nwell 85 27 85 27 2 Vdd
rlabel metal1 85 70 85 70 2 Vdd
port 2 ne
rlabel metal1 85 0 85 0 2 Gnd
port 3 ne
rlabel metal1 150 0 150 0 2 Gnd
port 3 ne
rlabel nwell 150 27 150 27 2 Vdd
rlabel metal1 150 60 150 60 2 Vdd
port 2 ne
rlabel metal1 222 60 222 60 2 Vdd
port 2 ne
rlabel metal1 222 0 222 0 2 Gnd
port 3 ne
<< end >>
