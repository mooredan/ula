magic
tech scmos
magscale 1 2
timestamp 1572801428
<< error_p >>
rect 94 700 96 701
rect 126 700 128 701
rect 132 700 134 701
rect 158 700 160 701
rect 164 700 166 701
rect 222 700 224 701
rect 228 700 230 701
rect 549 683 550 684
rect 555 670 556 671
rect 158 533 160 535
rect 164 533 166 535
rect 392 533 394 535
rect 482 533 484 535
rect 488 533 490 535
rect 578 533 580 535
<< nwell >>
rect 30 1208 572 1304
rect 28 950 572 1208
rect 28 850 570 950
rect 284 848 570 850
rect -12 507 606 677
rect -6 498 606 507
rect -6 22 22 498
rect 572 22 606 498
rect -6 -6 606 22
<< ntransistor >>
rect 38 706 42 766
rect 54 706 58 766
rect 88 706 92 766
rect 104 706 108 766
rect 120 706 124 766
rect 136 706 140 766
rect 152 706 156 766
rect 168 706 172 766
rect 184 706 188 766
rect 200 706 204 766
rect 216 706 220 766
rect 232 706 236 766
rect 248 706 252 766
rect 264 706 268 766
rect 280 706 284 766
rect 296 706 300 766
rect 396 707 400 767
rect 412 707 416 767
rect 428 707 432 767
rect 444 707 448 767
rect 460 707 464 767
rect 476 707 480 767
rect 492 707 496 767
rect 508 707 512 767
rect 524 707 528 767
rect 540 707 544 767
rect 556 707 560 767
rect 572 707 576 767
rect 76 432 276 438
rect 76 342 276 348
rect 76 300 276 306
rect 76 212 276 218
rect 76 170 276 176
rect 76 82 276 88
rect 324 432 524 438
rect 324 342 524 348
rect 324 300 524 306
rect 324 212 524 218
rect 324 170 524 176
rect 324 82 524 88
<< ptransistor >>
rect 76 1248 276 1254
rect 76 1160 276 1166
rect 76 1118 276 1124
rect 76 1032 276 1038
rect 76 990 276 996
rect 76 902 276 908
rect 324 1248 524 1254
rect 324 1160 524 1166
rect 324 1118 524 1124
rect 324 1032 524 1038
rect 324 990 524 996
rect 324 902 524 908
rect 38 539 42 643
rect 54 539 58 643
rect 88 539 92 643
rect 104 539 108 643
rect 120 539 124 643
rect 136 539 140 643
rect 152 539 156 643
rect 168 539 172 643
rect 184 539 188 643
rect 200 539 204 643
rect 216 539 220 643
rect 232 539 236 643
rect 248 539 252 643
rect 264 539 268 643
rect 280 539 284 643
rect 296 539 300 643
rect 396 539 400 643
rect 412 539 416 643
rect 428 539 432 643
rect 444 539 448 643
rect 460 539 464 643
rect 476 539 480 643
rect 492 539 496 643
rect 508 539 512 643
rect 524 539 528 643
rect 540 539 544 643
rect 556 539 560 643
rect 572 539 576 643
<< ndiffusion >>
rect 26 706 38 766
rect 42 706 54 766
rect 58 706 70 766
rect 76 706 88 766
rect 92 706 104 766
rect 108 706 120 766
rect 124 706 136 766
rect 140 706 152 766
rect 156 706 168 766
rect 172 706 184 766
rect 188 706 200 766
rect 204 706 216 766
rect 220 706 232 766
rect 236 706 248 766
rect 252 706 264 766
rect 268 706 280 766
rect 284 706 296 766
rect 300 706 312 766
rect 384 707 396 767
rect 400 707 412 767
rect 416 707 428 767
rect 432 707 444 767
rect 448 707 460 767
rect 464 707 476 767
rect 480 707 492 767
rect 496 707 508 767
rect 512 707 524 767
rect 528 707 540 767
rect 544 707 556 767
rect 560 707 572 767
rect 576 761 582 767
rect 576 707 586 761
rect 94 701 100 706
rect 126 701 134 706
rect 158 701 166 706
rect 222 701 230 706
rect 384 701 394 707
rect 418 701 426 707
rect 450 701 456 707
rect 482 701 490 707
rect 514 701 522 707
rect 546 701 552 707
rect 578 701 586 707
rect 76 438 276 456
rect 76 348 276 432
rect 76 306 276 342
rect 76 218 276 300
rect 76 176 276 212
rect 76 88 276 170
rect 76 64 276 82
rect 324 438 524 456
rect 324 348 524 432
rect 324 306 524 342
rect 324 218 524 300
rect 324 176 524 212
rect 324 88 524 170
rect 324 64 524 82
<< pdiffusion >>
rect 72 1260 280 1272
rect 76 1258 280 1260
rect 320 1260 528 1272
rect 320 1258 524 1260
rect 76 1254 276 1258
rect 76 1166 276 1248
rect 76 1124 276 1160
rect 76 1038 276 1118
rect 76 996 276 1032
rect 76 908 276 990
rect 76 884 276 902
rect 324 1254 524 1258
rect 324 1166 524 1248
rect 324 1124 524 1160
rect 324 1038 524 1118
rect 324 996 524 1032
rect 324 908 524 990
rect 324 884 524 902
rect 126 643 134 649
rect 158 643 166 649
rect 222 643 230 649
rect 384 643 394 649
rect 418 643 426 649
rect 450 643 456 649
rect 482 643 490 649
rect 514 643 522 649
rect 546 643 552 649
rect 578 643 586 649
rect 26 539 38 643
rect 42 539 54 643
rect 58 539 70 643
rect 76 539 88 643
rect 92 539 104 643
rect 108 539 120 643
rect 124 539 136 643
rect 140 539 152 643
rect 156 539 168 643
rect 172 539 184 643
rect 188 539 200 643
rect 204 539 216 643
rect 220 539 232 643
rect 236 539 248 643
rect 252 539 264 643
rect 268 539 280 643
rect 284 539 296 643
rect 300 539 312 643
rect 384 539 396 643
rect 400 539 412 643
rect 416 539 428 643
rect 432 539 444 643
rect 448 539 460 643
rect 464 539 476 643
rect 480 539 492 643
rect 496 539 508 643
rect 512 539 524 643
rect 528 539 540 643
rect 544 539 556 643
rect 560 539 572 643
rect 576 539 586 643
rect 158 535 166 539
rect 384 535 394 539
rect 482 535 490 539
rect 578 535 586 539
<< psubstratepdiff >>
rect 0 1314 600 1340
rect 0 840 22 1314
rect 234 840 294 842
rect 306 840 366 842
rect 578 840 600 1314
rect 0 820 600 840
rect 0 697 12 820
rect 586 767 600 820
rect 582 761 600 767
rect 0 690 14 697
rect 30 690 46 697
rect 94 695 100 701
rect 62 690 100 695
rect 126 695 134 701
rect 158 695 166 701
rect 0 689 100 690
rect 126 690 168 695
rect 222 697 230 701
rect 194 690 270 697
rect 384 697 394 701
rect 418 697 426 701
rect 450 697 456 701
rect 296 691 456 697
rect 482 697 490 701
rect 514 697 522 701
rect 546 697 552 701
rect 482 691 552 697
rect 586 701 600 761
rect 578 691 600 701
rect 296 690 600 691
rect 126 689 600 690
rect 0 683 600 689
rect 28 460 562 492
rect 28 60 60 460
rect 76 456 276 460
rect 76 60 276 64
rect 286 60 314 460
rect 324 456 524 460
rect 324 60 524 64
rect 540 60 562 460
rect 28 28 562 60
<< nsubstratendiff >>
rect 38 1272 562 1296
rect 38 1260 72 1272
rect 38 880 60 1260
rect 280 1258 320 1272
rect 528 1260 562 1272
rect 76 880 276 884
rect 284 880 316 1258
rect 324 880 524 884
rect 540 880 562 1260
rect 38 860 562 880
rect 0 659 600 665
rect 0 653 14 659
rect 0 523 12 653
rect 30 653 46 659
rect 62 653 100 659
rect 126 653 168 659
rect 126 649 134 653
rect 158 649 166 653
rect 194 653 244 659
rect 222 649 230 653
rect 270 653 456 659
rect 384 649 394 653
rect 418 649 426 653
rect 450 649 456 653
rect 482 653 552 659
rect 482 649 490 653
rect 514 649 522 653
rect 546 649 552 653
rect 578 649 600 659
rect 72 523 86 531
rect 158 531 166 535
rect 384 531 394 535
rect 482 531 490 535
rect 586 535 600 649
rect 578 531 600 535
rect 112 523 600 531
rect 0 504 600 523
rect 0 16 16 504
rect 578 16 600 504
rect 0 0 600 16
<< polysilicon >>
rect 62 1248 76 1254
rect 276 1248 282 1254
rect 62 1166 74 1248
rect 278 1166 282 1248
rect 62 1160 76 1166
rect 276 1160 282 1166
rect 62 1124 74 1160
rect 278 1124 282 1160
rect 62 1118 76 1124
rect 276 1118 282 1124
rect 62 1038 74 1118
rect 278 1038 282 1118
rect 62 1032 76 1038
rect 276 1032 282 1038
rect 62 996 74 1032
rect 278 996 282 1032
rect 62 990 76 996
rect 276 990 282 996
rect 62 908 74 990
rect 278 908 282 990
rect 62 902 76 908
rect 276 902 282 908
rect 318 1248 324 1254
rect 524 1248 538 1254
rect 318 1166 322 1248
rect 526 1166 538 1248
rect 318 1160 324 1166
rect 524 1160 538 1166
rect 318 1124 322 1160
rect 526 1124 538 1160
rect 318 1118 324 1124
rect 524 1118 538 1124
rect 318 1038 322 1118
rect 526 1038 538 1118
rect 318 1032 324 1038
rect 524 1032 538 1038
rect 318 996 322 1032
rect 526 996 538 1032
rect 318 990 324 996
rect 524 990 538 996
rect 318 908 322 990
rect 526 908 538 990
rect 318 902 324 908
rect 524 902 538 908
rect 222 790 580 810
rect 386 780 416 790
rect 38 766 42 770
rect 48 768 70 780
rect 88 768 156 772
rect 54 766 58 768
rect 88 766 92 768
rect 104 766 108 768
rect 120 766 124 768
rect 136 766 140 768
rect 152 766 156 768
rect 168 768 236 772
rect 168 766 172 768
rect 184 766 188 768
rect 200 766 204 768
rect 216 766 220 768
rect 232 766 236 768
rect 248 766 252 770
rect 264 766 268 770
rect 280 766 284 770
rect 296 766 300 770
rect 396 767 400 780
rect 412 770 432 774
rect 412 767 416 770
rect 428 767 432 770
rect 444 769 464 773
rect 444 767 448 769
rect 460 767 464 769
rect 476 767 480 771
rect 492 767 496 771
rect 508 769 528 773
rect 508 767 512 769
rect 524 767 528 769
rect 540 769 560 773
rect 540 767 544 769
rect 556 767 560 769
rect 572 767 576 772
rect 38 704 42 706
rect 54 704 58 706
rect 16 700 42 704
rect 16 692 28 700
rect 48 692 60 704
rect 88 700 92 706
rect 104 703 108 706
rect 120 703 124 706
rect 102 691 124 703
rect 136 701 140 706
rect 152 701 156 706
rect 168 704 172 706
rect 184 704 188 706
rect 168 699 192 704
rect 200 701 204 706
rect 216 701 220 706
rect 232 701 236 706
rect 248 704 252 706
rect 264 704 268 706
rect 280 704 284 706
rect 296 704 300 706
rect 170 692 192 699
rect 248 700 300 704
rect 396 705 400 707
rect 412 705 416 707
rect 396 701 416 705
rect 428 705 432 707
rect 444 705 448 707
rect 428 701 448 705
rect 460 705 464 707
rect 476 705 480 707
rect 272 692 294 700
rect 458 693 480 705
rect 492 705 496 707
rect 508 705 512 707
rect 492 701 512 705
rect 524 705 528 707
rect 540 705 544 707
rect 524 701 544 705
rect 556 705 560 707
rect 572 705 576 707
rect 554 693 576 705
rect 62 668 294 680
rect 16 649 28 657
rect 16 645 42 649
rect 48 645 60 657
rect 38 643 42 645
rect 54 643 58 645
rect 88 643 92 647
rect 102 645 124 657
rect 104 643 108 645
rect 120 643 124 645
rect 170 649 192 657
rect 136 643 140 647
rect 152 643 156 647
rect 168 645 192 649
rect 168 643 172 645
rect 184 643 188 645
rect 200 643 204 647
rect 216 643 220 647
rect 246 649 268 657
rect 232 643 236 647
rect 246 645 300 649
rect 248 643 252 645
rect 264 643 268 645
rect 280 643 284 645
rect 296 643 300 645
rect 396 647 416 651
rect 396 643 400 647
rect 412 643 416 647
rect 428 647 448 651
rect 428 643 432 647
rect 444 643 448 647
rect 458 645 480 657
rect 460 643 464 645
rect 476 643 480 645
rect 492 645 512 649
rect 492 643 496 645
rect 508 643 512 645
rect 524 645 544 649
rect 524 643 528 645
rect 540 643 544 645
rect 554 645 576 657
rect 556 643 560 645
rect 572 643 576 645
rect 38 537 42 539
rect 54 537 58 539
rect 88 537 92 539
rect 104 537 108 539
rect 120 537 124 539
rect 136 537 140 539
rect 152 537 156 539
rect 20 525 42 537
rect 48 525 70 537
rect 88 533 156 537
rect 88 525 110 533
rect 168 537 172 539
rect 184 537 188 539
rect 200 537 204 539
rect 216 537 220 539
rect 232 537 236 539
rect 168 533 236 537
rect 248 535 252 539
rect 264 535 268 539
rect 280 535 284 539
rect 296 535 300 539
rect 396 535 400 539
rect 412 537 416 539
rect 428 537 432 539
rect 412 533 432 537
rect 444 537 448 539
rect 460 537 464 539
rect 444 533 464 537
rect 476 535 480 539
rect 492 535 496 539
rect 508 537 512 539
rect 524 537 528 539
rect 508 533 528 537
rect 540 537 544 539
rect 556 537 560 539
rect 540 533 560 537
rect 572 535 576 539
rect 62 432 76 438
rect 276 432 284 438
rect 62 348 74 432
rect 278 348 284 432
rect 62 342 76 348
rect 276 342 284 348
rect 62 306 74 342
rect 278 306 284 342
rect 62 300 76 306
rect 276 300 284 306
rect 62 218 74 300
rect 278 218 284 300
rect 62 212 76 218
rect 276 212 284 218
rect 62 176 74 212
rect 278 176 284 212
rect 62 170 76 176
rect 276 170 284 176
rect 62 88 74 170
rect 278 88 284 170
rect 62 82 76 88
rect 276 82 284 88
rect 316 432 324 438
rect 524 432 538 438
rect 316 348 322 432
rect 526 348 538 432
rect 316 342 324 348
rect 524 342 538 348
rect 316 306 322 342
rect 526 306 538 342
rect 316 300 324 306
rect 524 300 538 306
rect 316 218 322 300
rect 526 218 538 300
rect 316 212 324 218
rect 524 212 538 218
rect 316 176 322 212
rect 526 176 538 212
rect 316 170 324 176
rect 524 170 538 176
rect 316 88 322 170
rect 526 88 538 170
rect 316 82 324 88
rect 524 82 538 88
<< metal1 >>
rect 124 1400 476 1480
rect 204 1380 396 1400
rect 224 1360 376 1380
rect 0 1316 232 1338
rect 0 850 20 1316
rect 28 1234 234 1310
rect 240 1308 360 1360
rect 368 1316 600 1338
rect 28 1184 58 1234
rect 64 1190 72 1228
rect 78 1184 104 1234
rect 240 1224 286 1308
rect 112 1191 286 1224
rect 28 1104 234 1184
rect 28 1054 58 1104
rect 64 1060 72 1098
rect 78 1054 104 1104
rect 240 1096 286 1191
rect 111 1061 286 1096
rect 28 976 234 1054
rect 28 860 58 976
rect 64 872 72 963
rect 78 924 104 976
rect 240 966 286 1061
rect 111 933 286 966
rect 78 878 232 924
rect 64 860 82 872
rect 88 860 232 878
rect 0 808 58 850
rect 0 708 22 808
rect 64 796 72 860
rect 78 820 231 850
rect 78 808 216 820
rect 240 814 286 933
rect 294 860 306 1296
rect 314 1224 360 1308
rect 366 1232 572 1310
rect 314 1191 489 1224
rect 314 1096 360 1191
rect 497 1181 522 1232
rect 528 1187 536 1225
rect 542 1181 572 1232
rect 366 1104 572 1181
rect 314 1061 489 1096
rect 314 966 360 1061
rect 497 1054 522 1104
rect 528 1060 536 1098
rect 542 1054 572 1104
rect 366 976 572 1054
rect 314 933 489 966
rect 296 820 304 850
rect 314 814 360 933
rect 497 924 522 976
rect 368 878 522 924
rect 368 860 512 878
rect 528 872 536 968
rect 518 860 536 872
rect 542 860 572 976
rect 580 850 600 1316
rect 368 820 600 850
rect 222 806 580 814
rect 64 787 83 796
rect 74 780 83 787
rect 222 786 380 806
rect 28 770 68 778
rect 74 774 262 780
rect 268 776 380 786
rect 386 780 416 800
rect 422 790 580 806
rect 422 780 457 790
rect 586 784 600 820
rect 254 770 262 774
rect 300 774 380 776
rect 422 774 430 780
rect 576 776 600 784
rect 300 770 430 774
rect 28 720 36 770
rect 44 714 52 764
rect 38 708 52 714
rect 60 716 68 764
rect 78 762 246 768
rect 78 721 86 762
rect 60 708 70 716
rect 94 714 102 756
rect 0 683 12 708
rect 18 694 26 702
rect 38 696 44 708
rect 0 640 12 665
rect 18 655 24 694
rect 32 684 44 696
rect 50 694 58 702
rect 50 678 56 694
rect 64 678 70 708
rect 76 708 102 714
rect 110 711 118 762
rect 126 708 134 756
rect 142 711 150 762
rect 76 685 98 708
rect 128 704 134 708
rect 158 704 166 756
rect 174 711 182 762
rect 190 708 198 756
rect 206 708 214 762
rect 104 693 122 701
rect 40 670 58 678
rect 64 670 82 678
rect 18 647 26 655
rect 32 653 44 664
rect 38 641 44 653
rect 50 655 56 670
rect 50 647 58 655
rect 64 641 70 670
rect 0 544 22 640
rect 38 635 52 641
rect 28 547 36 629
rect 44 553 52 635
rect 60 632 70 641
rect 76 641 98 663
rect 106 655 112 693
rect 128 685 166 704
rect 172 694 190 702
rect 222 697 230 756
rect 238 720 246 762
rect 254 764 294 770
rect 316 766 430 770
rect 436 767 474 773
rect 254 714 262 764
rect 184 678 190 694
rect 196 684 230 697
rect 236 708 262 714
rect 270 714 278 758
rect 286 720 294 764
rect 302 714 310 764
rect 270 708 310 714
rect 160 670 178 678
rect 184 670 202 678
rect 104 647 122 655
rect 128 646 166 664
rect 172 655 178 670
rect 172 647 190 655
rect 196 653 230 664
rect 76 635 103 641
rect 128 640 134 646
rect 0 12 16 544
rect 28 541 54 547
rect 60 541 68 632
rect 78 547 86 629
rect 93 553 103 635
rect 110 549 118 640
rect 125 555 134 640
rect 110 547 120 549
rect 78 541 120 547
rect 48 535 54 541
rect 114 539 120 541
rect 142 539 150 640
rect 157 637 166 646
rect 157 545 167 637
rect 174 539 182 641
rect 189 545 199 637
rect 206 539 214 640
rect 222 553 230 653
rect 236 640 242 708
rect 248 686 268 697
rect 274 694 292 702
rect 280 678 286 694
rect 248 670 266 678
rect 274 670 292 678
rect 254 655 260 670
rect 248 647 266 655
rect 272 653 296 664
rect 302 641 308 708
rect 236 634 278 640
rect 236 629 246 634
rect 238 547 246 629
rect 221 541 246 547
rect 254 550 262 627
rect 270 556 278 634
rect 286 635 308 641
rect 286 550 294 635
rect 254 542 294 550
rect 221 539 228 541
rect 22 527 40 535
rect 48 527 68 535
rect 90 527 108 535
rect 114 533 228 539
rect 254 535 262 542
rect 302 541 310 629
rect 234 529 262 535
rect 316 532 380 766
rect 436 760 442 767
rect 386 709 394 760
rect 402 754 442 760
rect 402 709 410 754
rect 388 697 394 709
rect 418 697 426 748
rect 388 673 426 697
rect 434 709 442 754
rect 448 709 458 761
rect 466 709 474 767
rect 498 767 570 773
rect 482 709 490 765
rect 498 709 506 767
rect 434 678 440 709
rect 448 694 454 709
rect 460 695 478 703
rect 484 697 490 709
rect 514 697 522 761
rect 446 686 454 694
rect 434 670 452 678
rect 388 653 426 665
rect 388 637 394 653
rect 22 521 28 527
rect 22 494 72 521
rect 22 26 28 494
rect 34 443 72 486
rect 78 484 84 514
rect 78 464 86 484
rect 34 75 58 443
rect 78 434 84 464
rect 64 428 84 434
rect 64 86 72 428
rect 34 32 86 75
rect 46 28 80 32
rect 94 26 100 527
rect 114 521 228 527
rect 106 508 228 521
rect 106 506 216 508
rect 106 494 214 506
rect 234 502 240 529
rect 269 523 380 532
rect 222 494 240 502
rect 246 492 380 523
rect 386 521 394 637
rect 402 535 410 641
rect 418 545 426 653
rect 434 641 440 670
rect 446 655 454 663
rect 466 655 472 695
rect 484 685 522 697
rect 530 713 538 767
rect 448 641 454 655
rect 460 647 478 655
rect 484 653 522 665
rect 484 641 490 653
rect 434 535 442 641
rect 448 545 458 641
rect 466 535 474 641
rect 402 527 474 535
rect 386 494 460 521
rect 466 500 474 527
rect 482 521 490 641
rect 498 535 506 641
rect 514 545 522 653
rect 530 641 536 713
rect 544 710 554 761
rect 544 697 550 710
rect 562 709 570 767
rect 578 709 600 776
rect 542 683 550 697
rect 556 695 574 703
rect 561 678 567 695
rect 580 683 600 709
rect 555 670 573 678
rect 542 653 550 665
rect 561 655 567 670
rect 544 641 550 653
rect 556 647 574 655
rect 580 641 600 665
rect 530 535 538 641
rect 544 545 554 641
rect 562 535 570 641
rect 498 527 570 535
rect 480 507 508 521
rect 466 492 506 500
rect 246 488 352 492
rect 106 419 240 486
rect 246 411 286 488
rect 106 371 286 411
rect 106 286 240 365
rect 246 278 286 371
rect 112 241 286 278
rect 106 157 240 234
rect 246 148 286 241
rect 106 112 286 148
rect 107 36 238 105
rect 114 28 238 36
rect 246 98 286 112
rect 294 108 306 481
rect 314 411 352 488
rect 359 419 494 486
rect 314 371 494 411
rect 314 278 352 371
rect 360 286 494 365
rect 314 241 494 278
rect 314 148 352 241
rect 360 157 494 234
rect 314 112 494 148
rect 314 98 352 112
rect 22 18 40 26
rect 88 18 106 26
rect 246 25 352 98
rect 360 32 494 105
rect 360 28 482 32
rect 500 26 506 492
rect 488 18 506 26
rect 514 26 520 527
rect 578 521 600 641
rect 527 494 600 521
rect 527 464 535 484
rect 528 434 535 464
rect 528 86 536 434
rect 542 75 572 486
rect 526 32 572 75
rect 538 28 572 32
rect 514 18 532 26
rect 578 16 600 494
rect 48 12 82 16
rect 113 12 482 16
rect 538 12 600 16
rect 0 0 600 12
<< metal2 >>
rect 0 1190 600 1340
rect 0 1180 104 1190
rect 284 1180 316 1190
rect 497 1180 600 1190
rect 0 1040 600 1180
rect 0 1030 104 1040
rect 284 1030 316 1040
rect 500 1030 600 1040
rect 0 880 600 1030
rect 0 878 58 880
rect 90 874 510 880
rect 542 878 600 880
rect 64 866 82 872
rect 518 866 536 872
rect 64 860 536 866
rect 72 858 536 860
rect 20 845 576 850
rect 0 777 600 845
rect 0 767 68 777
rect 123 767 163 777
rect 238 767 280 777
rect 381 767 421 777
rect 500 767 600 777
rect 0 737 600 767
rect 0 710 230 737
rect 238 720 278 728
rect 286 710 600 737
rect 0 686 600 710
rect 273 683 426 686
rect 484 685 522 686
rect 40 677 58 678
rect 184 677 202 678
rect 248 677 266 678
rect 40 671 266 677
rect 388 673 426 683
rect 434 677 452 678
rect 555 677 573 678
rect 40 670 58 671
rect 184 670 202 671
rect 248 670 266 671
rect 434 671 573 677
rect 434 670 452 671
rect 555 670 573 671
rect 16 662 36 663
rect 62 662 180 663
rect 206 662 230 663
rect 16 652 230 662
rect 273 659 426 665
rect 484 659 522 663
rect 273 652 522 659
rect 0 637 600 652
rect 0 612 262 637
rect 270 621 310 629
rect 318 612 600 637
rect 0 582 600 612
rect 0 572 36 582
rect 92 572 136 582
rect 188 572 232 582
rect 336 572 379 582
rect 447 572 490 582
rect 561 572 600 582
rect 0 510 600 572
rect 0 492 214 510
rect 222 484 240 502
rect 248 492 600 510
rect 78 476 535 484
rect 78 464 86 476
rect 0 456 70 460
rect 108 456 492 466
rect 527 464 535 476
rect 542 456 600 460
rect 0 310 600 456
rect 0 300 100 310
rect 286 300 314 310
rect 500 300 600 310
rect 0 160 600 300
rect 0 150 100 160
rect 286 150 314 160
rect 500 150 600 160
rect 0 47 600 150
rect 0 38 246 47
rect 0 0 14 38
rect 22 0 40 26
rect 48 0 80 38
rect 88 0 106 26
rect 114 0 246 38
rect 256 0 344 39
rect 352 35 600 47
rect 352 0 480 35
rect 488 0 506 26
rect 514 0 532 26
rect 540 0 600 35
<< labels >>
flabel nwell 0 -6 0 -6 4 FreeSans 20 0 0 0 VddNW
flabel nwell 600 -6 600 -6 6 FreeSans 20 0 0 0 VddNW
flabel psubstratepdiff 600 686 600 686 6 FreeSans 20 0 0 0 GndAct
flabel psubstratepdiff 0 686 0 686 4 FreeSans 20 0 0 0 GndAct
flabel metal2 600 0 600 0 6 FreeSans 20 0 0 0 VddAct
flabel metal2 0 0 0 0 4 FreeSans 20 0 0 0 VddAct
flabel metal1 466 683 466 683 4 FreeSans 80 0 0 0 DIunbuf
flabel metal1 434 683 434 683 6 FreeSans 80 0 0 0 DIB
flabel metal1 530 683 530 683 4 FreeSans 80 0 0 0 DI
flabel psubstratepdiff 31 683 31 683 6 FreeSans 64 0 0 0 OEN
flabel metal1 54 683 54 683 6 FreeSans 64 0 0 0 OEB
flabel metal1 69 667 69 667 2 FreeSans 64 0 0 0 OE
flabel metal2 88 0 88 0 2 FreeSans 80 0 0 0 DO
flabel metal2 256 0 256 0 2 FreeSans 80 0 0 0 DATA
flabel metal2 22 0 22 0 2 FreeSans 80 0 0 0 OEN
flabel metal2 514 0 514 0 2 FreeSans 80 0 0 0 DI
flabel metal2 488 0 488 0 8 FreeSans 80 0 0 0 DIB
flabel metal2 88 0 88 0 6 FreeSans 80 0 0 0 DO
flabel metal2 600 492 600 492 6 FreeSans 20 0 0 0 VddM2B
flabel metal2 0 492 0 492 4 FreeSans 20 0 0 0 VddM2B
flabel metal2 600 880 600 880 6 FreeSans 20 0 0 0 VddM2A
flabel metal2 0 880 0 880 4 FreeSans 20 0 0 0 VddM2A
flabel metal2 0 688 0 688 4 FreeSans 20 0 0 0 GndM2B
flabel metal2 600 688 600 688 6 FreeSans 20 0 0 0 GndM2B
flabel metal2 600 0 600 0 6 FreeSans 20 0 0 0 GndM2A
flabel metal2 0 0 0 0 4 FreeSans 20 0 0 0 GndM2A
<< end >>
