magic
tech amic5n
timestamp 1621830667
<< nwell >>
rect -120 870 1320 2430
<< ntransistor >>
rect 210 120 270 690
rect 450 120 510 690
rect 930 120 990 690
<< ptransistor >>
rect 210 1210 270 1780
rect 450 1210 510 1780
rect 930 1050 990 2250
<< nselect >>
rect 0 60 1200 750
<< pselect >>
rect 0 990 1200 2310
<< ndiffusion >>
rect 60 655 210 690
rect 60 605 95 655
rect 145 605 210 655
rect 60 505 210 605
rect 60 455 95 505
rect 145 455 210 505
rect 60 355 210 455
rect 60 305 95 355
rect 145 305 210 355
rect 60 205 210 305
rect 60 155 95 205
rect 145 155 210 205
rect 60 120 210 155
rect 270 120 450 690
rect 510 655 660 690
rect 510 605 575 655
rect 625 605 660 655
rect 510 475 660 605
rect 510 425 575 475
rect 625 425 660 475
rect 510 265 660 425
rect 510 215 575 265
rect 625 215 660 265
rect 510 120 660 215
rect 780 475 930 690
rect 780 425 815 475
rect 865 425 930 475
rect 780 205 930 425
rect 780 155 815 205
rect 865 155 930 205
rect 780 120 930 155
rect 990 655 1140 690
rect 990 605 1055 655
rect 1105 605 1140 655
rect 990 445 1140 605
rect 990 395 1055 445
rect 1105 395 1140 445
rect 990 265 1140 395
rect 990 215 1055 265
rect 1105 215 1140 265
rect 990 120 1140 215
<< pdiffusion >>
rect 660 2215 930 2250
rect 660 2165 815 2215
rect 865 2165 930 2215
rect 660 2035 930 2165
rect 660 1985 815 2035
rect 865 1985 930 2035
rect 660 1885 930 1985
rect 660 1835 815 1885
rect 865 1835 930 1885
rect 660 1780 930 1835
rect 60 1745 210 1780
rect 60 1695 95 1745
rect 145 1695 210 1745
rect 60 1595 210 1695
rect 60 1545 95 1595
rect 145 1545 210 1595
rect 60 1445 210 1545
rect 60 1395 95 1445
rect 145 1395 210 1445
rect 60 1295 210 1395
rect 60 1245 95 1295
rect 145 1245 210 1295
rect 60 1210 210 1245
rect 270 1745 450 1780
rect 270 1695 335 1745
rect 385 1695 450 1745
rect 270 1595 450 1695
rect 270 1545 335 1595
rect 385 1545 450 1595
rect 270 1445 450 1545
rect 270 1395 335 1445
rect 385 1395 450 1445
rect 270 1295 450 1395
rect 270 1245 335 1295
rect 385 1245 450 1295
rect 270 1210 450 1245
rect 510 1745 930 1780
rect 510 1695 575 1745
rect 625 1735 930 1745
rect 625 1695 815 1735
rect 510 1685 815 1695
rect 865 1685 930 1735
rect 510 1595 930 1685
rect 510 1545 575 1595
rect 625 1585 930 1595
rect 625 1545 815 1585
rect 510 1535 815 1545
rect 865 1535 930 1585
rect 510 1445 930 1535
rect 510 1395 575 1445
rect 625 1435 930 1445
rect 625 1395 815 1435
rect 510 1385 815 1395
rect 865 1385 930 1435
rect 510 1295 930 1385
rect 510 1245 575 1295
rect 625 1285 930 1295
rect 625 1245 815 1285
rect 510 1235 815 1245
rect 865 1235 930 1285
rect 510 1210 930 1235
rect 640 1135 930 1210
rect 640 1085 815 1135
rect 865 1085 930 1135
rect 640 1050 930 1085
rect 990 2155 1140 2250
rect 990 2105 1055 2155
rect 1105 2105 1140 2155
rect 990 2005 1140 2105
rect 990 1955 1055 2005
rect 1105 1955 1140 2005
rect 990 1825 1140 1955
rect 990 1775 1055 1825
rect 1105 1775 1140 1825
rect 990 1645 1140 1775
rect 990 1595 1055 1645
rect 1105 1595 1140 1645
rect 990 1465 1140 1595
rect 990 1415 1055 1465
rect 1105 1415 1140 1465
rect 990 1285 1140 1415
rect 990 1235 1055 1285
rect 1105 1235 1140 1285
rect 990 1135 1140 1235
rect 990 1085 1055 1135
rect 1105 1085 1140 1135
rect 990 1050 1140 1085
<< ndcontact >>
rect 95 605 145 655
rect 95 455 145 505
rect 95 305 145 355
rect 95 155 145 205
rect 575 605 625 655
rect 575 425 625 475
rect 575 215 625 265
rect 815 425 865 475
rect 815 155 865 205
rect 1055 605 1105 655
rect 1055 395 1105 445
rect 1055 215 1105 265
<< pdcontact >>
rect 815 2165 865 2215
rect 815 1985 865 2035
rect 815 1835 865 1885
rect 95 1695 145 1745
rect 95 1545 145 1595
rect 95 1395 145 1445
rect 95 1245 145 1295
rect 335 1695 385 1745
rect 335 1545 385 1595
rect 335 1395 385 1445
rect 335 1245 385 1295
rect 575 1695 625 1745
rect 815 1685 865 1735
rect 575 1545 625 1595
rect 815 1535 865 1585
rect 575 1395 625 1445
rect 815 1385 865 1435
rect 575 1245 625 1295
rect 815 1235 865 1285
rect 815 1085 865 1135
rect 1055 2105 1105 2155
rect 1055 1955 1105 2005
rect 1055 1775 1105 1825
rect 1055 1595 1105 1645
rect 1055 1415 1105 1465
rect 1055 1235 1105 1285
rect 1055 1085 1105 1135
<< polysilicon >>
rect 930 2250 990 2315
rect 210 1780 270 1845
rect 450 1780 510 1845
rect 210 1120 270 1210
rect 60 1055 270 1120
rect 60 1005 125 1055
rect 175 1005 270 1055
rect 60 940 270 1005
rect 210 690 270 940
rect 450 960 510 1210
rect 930 960 990 1050
rect 450 895 660 960
rect 450 845 545 895
rect 595 845 660 895
rect 450 780 660 845
rect 750 895 990 960
rect 750 845 815 895
rect 865 845 990 895
rect 750 780 990 845
rect 450 690 510 780
rect 930 690 990 780
rect 210 55 270 120
rect 450 55 510 120
rect 930 55 990 120
<< polycontact >>
rect 125 1005 175 1055
rect 545 845 595 895
rect 815 845 865 895
<< metal1 >>
rect 0 2280 1200 2370
rect 60 1745 180 2280
rect 660 2215 900 2280
rect 660 2165 815 2215
rect 865 2165 900 2215
rect 660 2035 900 2165
rect 660 1985 815 2035
rect 865 1985 900 2035
rect 660 1885 900 1985
rect 660 1835 815 1885
rect 865 1835 900 1885
rect 660 1780 900 1835
rect 60 1695 95 1745
rect 145 1695 180 1745
rect 60 1595 180 1695
rect 60 1545 95 1595
rect 145 1545 180 1595
rect 60 1445 180 1545
rect 60 1395 95 1445
rect 145 1395 180 1445
rect 60 1295 180 1395
rect 60 1245 95 1295
rect 145 1245 180 1295
rect 60 1210 180 1245
rect 300 1745 420 1780
rect 300 1695 335 1745
rect 385 1695 420 1745
rect 300 1595 420 1695
rect 300 1545 335 1595
rect 385 1545 420 1595
rect 300 1445 420 1545
rect 300 1395 335 1445
rect 385 1395 420 1445
rect 300 1295 420 1395
rect 300 1245 335 1295
rect 385 1245 420 1295
rect 90 1055 210 1090
rect 90 1005 125 1055
rect 175 1005 210 1055
rect 90 970 210 1005
rect 300 720 420 1245
rect 540 1745 900 1780
rect 540 1695 575 1745
rect 625 1735 900 1745
rect 625 1695 815 1735
rect 540 1685 815 1695
rect 865 1685 900 1735
rect 540 1595 900 1685
rect 540 1545 575 1595
rect 625 1585 900 1595
rect 625 1545 815 1585
rect 540 1535 815 1545
rect 865 1535 900 1585
rect 540 1445 900 1535
rect 540 1395 575 1445
rect 625 1435 900 1445
rect 625 1395 815 1435
rect 540 1385 815 1395
rect 865 1385 900 1435
rect 540 1295 900 1385
rect 540 1245 575 1295
rect 625 1285 900 1295
rect 625 1245 815 1285
rect 540 1235 815 1245
rect 865 1235 900 1285
rect 540 1210 900 1235
rect 640 1135 900 1210
rect 640 1085 815 1135
rect 865 1085 900 1135
rect 640 1050 900 1085
rect 1020 2155 1140 2190
rect 1020 2105 1055 2155
rect 1105 2105 1140 2155
rect 1020 2005 1140 2105
rect 1020 1955 1055 2005
rect 1105 1955 1140 2005
rect 1020 1825 1140 1955
rect 1020 1775 1055 1825
rect 1105 1775 1140 1825
rect 1020 1645 1140 1775
rect 1020 1595 1055 1645
rect 1105 1595 1140 1645
rect 1020 1465 1140 1595
rect 1020 1415 1055 1465
rect 1105 1415 1140 1465
rect 1020 1285 1140 1415
rect 1020 1235 1055 1285
rect 1105 1235 1140 1285
rect 1020 1135 1140 1235
rect 1020 1085 1055 1135
rect 1105 1085 1140 1135
rect 510 895 630 930
rect 510 845 545 895
rect 595 845 630 895
rect 510 810 630 845
rect 780 895 900 930
rect 780 845 815 895
rect 865 845 900 895
rect 780 720 900 845
rect 60 655 180 690
rect 60 605 95 655
rect 145 605 180 655
rect 60 505 180 605
rect 300 655 900 720
rect 300 605 575 655
rect 625 605 900 655
rect 300 600 900 605
rect 1020 655 1140 1085
rect 1020 605 1055 655
rect 1105 605 1140 655
rect 300 570 660 600
rect 60 455 95 505
rect 145 455 180 505
rect 60 355 180 455
rect 60 305 95 355
rect 145 305 180 355
rect 60 205 180 305
rect 60 155 95 205
rect 145 155 180 205
rect 540 475 660 570
rect 540 425 575 475
rect 625 425 660 475
rect 540 265 660 425
rect 540 215 575 265
rect 625 215 660 265
rect 540 180 660 215
rect 780 475 900 510
rect 780 425 815 475
rect 865 425 900 475
rect 780 205 900 425
rect 60 90 180 155
rect 780 155 815 205
rect 865 155 900 205
rect 1020 445 1140 605
rect 1020 395 1055 445
rect 1105 395 1140 445
rect 1020 265 1140 395
rect 1020 215 1055 265
rect 1105 215 1140 265
rect 1020 180 1140 215
rect 780 90 900 155
rect 0 0 1200 90
<< labels >>
flabel nwell 0 930 0 930 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 30 30 30 30 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 30 2310 30 2310 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel ndiffusion s 360 330 360 330 2 FreeSans 400 0 0 0 x1
flabel metal1 s 570 870 570 870 2 FreeSans 400 0 0 0 b
port 3 ne
flabel metal1 s 1080 810 1080 810 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 690 630 690 630 2 FreeSans 400 0 0 0 n1
flabel metal1 s 150 1030 150 1030 2 FreeSans 400 0 0 0 a
port 2 ne
<< end >>
