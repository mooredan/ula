`celldefine
module tie1_b (z);
  output z;

  assign z = 1'b1;
endmodule
`endcelldefine
