magic
tech amic5n
timestamp 1624142566
<< nwell >>
rect -130 550 2080 1495
<< ntransistor >>
rect 225 275 285 400
rect 615 95 675 400
rect 1250 95 1310 400
rect 1665 205 1725 330
<< ptransistor >>
rect 225 745 285 930
rect 615 700 675 1345
rect 805 700 865 1345
rect 1060 700 1120 1345
rect 1250 700 1310 1345
rect 1665 745 1725 930
<< nselect >>
rect 110 1090 320 1300
rect 1630 1090 1840 1300
rect -10 295 1960 430
rect -10 100 850 295
rect 1080 100 1960 295
rect -10 0 1960 100
<< pselect >>
rect -10 1300 1960 1440
rect -10 1090 110 1300
rect 320 1090 1630 1300
rect 1840 1090 1960 1300
rect -10 670 1960 1090
rect 850 100 1080 295
<< ndiffusion >>
rect 75 370 225 400
rect 75 320 115 370
rect 165 320 225 370
rect 75 275 225 320
rect 285 370 405 400
rect 285 320 325 370
rect 375 320 405 370
rect 285 275 405 320
rect 495 370 615 400
rect 495 320 525 370
rect 575 320 615 370
rect 75 270 195 275
rect 75 220 115 270
rect 165 220 195 270
rect 75 190 195 220
rect 495 175 615 320
rect 495 125 525 175
rect 575 125 615 175
rect 495 95 615 125
rect 675 370 795 400
rect 675 320 715 370
rect 765 320 795 370
rect 675 175 795 320
rect 1130 370 1250 400
rect 1130 320 1160 370
rect 1210 320 1250 370
rect 675 125 715 175
rect 765 125 795 175
rect 1130 175 1250 320
rect 675 95 795 125
rect 1130 125 1160 175
rect 1210 125 1250 175
rect 1130 95 1250 125
rect 1310 355 1430 400
rect 1310 305 1350 355
rect 1400 305 1430 355
rect 1310 175 1430 305
rect 1545 300 1665 330
rect 1545 250 1575 300
rect 1625 250 1665 300
rect 1545 205 1665 250
rect 1725 300 1875 330
rect 1725 250 1785 300
rect 1835 250 1875 300
rect 1725 205 1875 250
rect 1310 125 1350 175
rect 1400 125 1430 175
rect 1755 200 1875 205
rect 1755 150 1785 200
rect 1835 150 1875 200
rect 1310 95 1430 125
rect 1755 120 1875 150
<< pdiffusion >>
rect 495 1315 615 1345
rect 495 1265 525 1315
rect 575 1265 615 1315
rect 495 1200 615 1265
rect 495 1150 525 1200
rect 575 1150 615 1200
rect 495 1065 615 1150
rect 495 1015 525 1065
rect 575 1015 615 1065
rect 75 930 195 955
rect 495 945 615 1015
rect 75 925 225 930
rect 75 875 115 925
rect 165 875 225 925
rect 75 825 225 875
rect 75 775 115 825
rect 165 775 225 825
rect 75 745 225 775
rect 285 860 405 930
rect 285 810 325 860
rect 375 810 405 860
rect 285 745 405 810
rect 495 895 525 945
rect 575 895 615 945
rect 495 825 615 895
rect 495 775 525 825
rect 575 775 615 825
rect 495 700 615 775
rect 675 1315 805 1345
rect 675 1265 715 1315
rect 765 1265 805 1315
rect 675 1215 805 1265
rect 675 1165 715 1215
rect 765 1165 805 1215
rect 675 1115 805 1165
rect 675 1065 715 1115
rect 765 1065 805 1115
rect 675 985 805 1065
rect 675 935 715 985
rect 765 935 805 985
rect 675 700 805 935
rect 865 1315 1060 1345
rect 865 1265 925 1315
rect 975 1265 1060 1315
rect 865 1200 1060 1265
rect 865 1150 925 1200
rect 975 1150 1060 1200
rect 865 1065 1060 1150
rect 865 1015 925 1065
rect 975 1015 1060 1065
rect 865 945 1060 1015
rect 865 895 925 945
rect 975 895 1060 945
rect 865 825 1060 895
rect 865 775 925 825
rect 975 775 1060 825
rect 865 700 1060 775
rect 1120 1155 1250 1345
rect 1120 1105 1160 1155
rect 1210 1105 1250 1155
rect 1120 1015 1250 1105
rect 1120 965 1160 1015
rect 1210 965 1250 1015
rect 1120 915 1250 965
rect 1120 865 1160 915
rect 1210 865 1250 915
rect 1120 815 1250 865
rect 1120 765 1160 815
rect 1210 765 1250 815
rect 1120 700 1250 765
rect 1310 1315 1430 1345
rect 1310 1265 1350 1315
rect 1400 1265 1430 1315
rect 1310 1180 1430 1265
rect 1310 1130 1350 1180
rect 1400 1130 1430 1180
rect 1310 1080 1430 1130
rect 1310 1030 1350 1080
rect 1400 1030 1430 1080
rect 1310 980 1430 1030
rect 1310 930 1350 980
rect 1400 930 1430 980
rect 1755 930 1875 955
rect 1310 880 1430 930
rect 1310 830 1350 880
rect 1400 830 1430 880
rect 1310 780 1430 830
rect 1310 730 1350 780
rect 1400 730 1430 780
rect 1545 860 1665 930
rect 1545 810 1575 860
rect 1625 810 1665 860
rect 1545 745 1665 810
rect 1725 925 1875 930
rect 1725 875 1785 925
rect 1835 875 1875 925
rect 1725 825 1875 875
rect 1725 775 1785 825
rect 1835 775 1875 825
rect 1725 745 1875 775
rect 1310 700 1430 730
<< psubstratepdiff >>
rect 905 220 1015 250
rect 905 170 935 220
rect 985 170 1015 220
rect 905 140 1015 170
<< nsubstratendiff >>
rect 140 1225 280 1255
rect 140 1175 185 1225
rect 235 1175 280 1225
rect 140 1145 280 1175
rect 1670 1225 1810 1255
rect 1670 1175 1715 1225
rect 1765 1175 1810 1225
rect 1670 1145 1810 1175
<< nsubstratencontact >>
rect 185 1175 235 1225
rect 1715 1175 1765 1225
<< psubstratepcontact >>
rect 935 170 985 220
<< ndcontact >>
rect 115 320 165 370
rect 325 320 375 370
rect 525 320 575 370
rect 115 220 165 270
rect 525 125 575 175
rect 715 320 765 370
rect 1160 320 1210 370
rect 715 125 765 175
rect 1160 125 1210 175
rect 1350 305 1400 355
rect 1575 250 1625 300
rect 1785 250 1835 300
rect 1350 125 1400 175
rect 1785 150 1835 200
<< pdcontact >>
rect 525 1265 575 1315
rect 525 1150 575 1200
rect 525 1015 575 1065
rect 115 875 165 925
rect 115 775 165 825
rect 325 810 375 860
rect 525 895 575 945
rect 525 775 575 825
rect 715 1265 765 1315
rect 715 1165 765 1215
rect 715 1065 765 1115
rect 715 935 765 985
rect 925 1265 975 1315
rect 925 1150 975 1200
rect 925 1015 975 1065
rect 925 895 975 945
rect 925 775 975 825
rect 1160 1105 1210 1155
rect 1160 965 1210 1015
rect 1160 865 1210 915
rect 1160 765 1210 815
rect 1350 1265 1400 1315
rect 1350 1130 1400 1180
rect 1350 1030 1400 1080
rect 1350 930 1400 980
rect 1350 830 1400 880
rect 1350 730 1400 780
rect 1575 810 1625 860
rect 1785 875 1835 925
rect 1785 775 1835 825
<< polysilicon >>
rect 615 1345 675 1410
rect 805 1345 865 1410
rect 1060 1345 1120 1410
rect 1250 1345 1310 1410
rect 225 930 285 995
rect 225 685 285 745
rect 1665 930 1725 995
rect 115 665 285 685
rect 115 615 135 665
rect 185 615 285 665
rect 115 595 285 615
rect 225 400 285 595
rect 615 630 675 700
rect 805 630 865 700
rect 615 610 865 630
rect 615 560 675 610
rect 725 560 865 610
rect 615 540 865 560
rect 1060 560 1120 700
rect 1250 560 1310 700
rect 1060 540 1470 560
rect 615 400 675 540
rect 1060 490 1400 540
rect 1450 490 1470 540
rect 1060 470 1470 490
rect 1665 525 1725 745
rect 1665 505 1835 525
rect 1250 400 1310 470
rect 1665 455 1765 505
rect 1815 455 1835 505
rect 1665 435 1835 455
rect 225 210 285 275
rect 1665 330 1725 435
rect 1665 140 1725 205
rect 615 30 675 95
rect 1250 30 1310 95
<< polycontact >>
rect 135 615 185 665
rect 675 560 725 610
rect 1400 490 1450 540
rect 1765 455 1815 505
<< metal1 >>
rect 0 1395 1950 1485
rect 95 1245 185 1395
rect 505 1315 595 1335
rect 505 1265 525 1315
rect 575 1265 595 1315
rect 95 1225 255 1245
rect 95 1175 185 1225
rect 235 1175 255 1225
rect 95 1155 255 1175
rect 505 1200 595 1265
rect 95 925 185 1155
rect 95 875 115 925
rect 165 875 185 925
rect 505 1150 525 1200
rect 575 1150 595 1200
rect 505 1065 595 1150
rect 505 1015 525 1065
rect 575 1015 595 1065
rect 505 945 595 1015
rect 505 895 525 945
rect 575 895 595 945
rect 695 1315 785 1395
rect 695 1265 715 1315
rect 765 1265 785 1315
rect 695 1215 785 1265
rect 695 1165 715 1215
rect 765 1165 785 1215
rect 695 1115 785 1165
rect 695 1065 715 1115
rect 765 1065 785 1115
rect 695 985 785 1065
rect 695 935 715 985
rect 765 935 785 985
rect 695 915 785 935
rect 905 1325 995 1335
rect 1330 1325 1420 1335
rect 905 1315 1420 1325
rect 905 1265 925 1315
rect 975 1265 1350 1315
rect 1400 1265 1420 1315
rect 905 1235 1420 1265
rect 1765 1245 1855 1395
rect 905 1200 995 1235
rect 905 1150 925 1200
rect 975 1150 995 1200
rect 1330 1180 1420 1235
rect 905 1065 995 1150
rect 905 1015 925 1065
rect 975 1015 995 1065
rect 905 945 995 1015
rect 95 825 185 875
rect 95 775 115 825
rect 165 775 185 825
rect 95 745 185 775
rect 305 860 395 890
rect 305 810 325 860
rect 375 810 395 860
rect 30 665 205 685
rect 30 615 135 665
rect 185 615 205 665
rect 30 595 205 615
rect 305 630 395 810
rect 505 845 595 895
rect 905 895 925 945
rect 975 895 995 945
rect 905 845 995 895
rect 505 825 995 845
rect 505 775 525 825
rect 575 775 925 825
rect 975 775 995 825
rect 505 755 995 775
rect 1140 1155 1230 1175
rect 1140 1105 1160 1155
rect 1210 1105 1230 1155
rect 1140 1015 1230 1105
rect 1140 965 1160 1015
rect 1210 965 1230 1015
rect 1140 915 1230 965
rect 1140 865 1160 915
rect 1210 865 1230 915
rect 1140 815 1230 865
rect 1140 765 1160 815
rect 1210 765 1230 815
rect 305 610 745 630
rect 305 560 675 610
rect 725 560 745 610
rect 305 540 745 560
rect 95 370 185 390
rect 95 320 115 370
rect 165 320 185 370
rect 95 270 185 320
rect 305 370 395 540
rect 1140 390 1230 765
rect 1330 1130 1350 1180
rect 1400 1130 1420 1180
rect 1695 1225 1855 1245
rect 1695 1175 1715 1225
rect 1765 1175 1855 1225
rect 1695 1155 1855 1175
rect 1330 1080 1420 1130
rect 1330 1030 1350 1080
rect 1400 1030 1420 1080
rect 1330 980 1420 1030
rect 1330 930 1350 980
rect 1400 930 1420 980
rect 1330 880 1420 930
rect 1765 925 1855 1155
rect 1330 830 1350 880
rect 1400 830 1420 880
rect 1330 780 1420 830
rect 1330 730 1350 780
rect 1400 730 1420 780
rect 1330 710 1420 730
rect 1555 860 1645 890
rect 1555 810 1575 860
rect 1625 810 1645 860
rect 1555 560 1645 810
rect 1765 875 1785 925
rect 1835 875 1855 925
rect 1765 825 1855 875
rect 1765 775 1785 825
rect 1835 775 1855 825
rect 1765 745 1855 775
rect 1380 540 1645 560
rect 1380 490 1400 540
rect 1450 490 1645 540
rect 1380 470 1645 490
rect 305 320 325 370
rect 375 320 395 370
rect 305 285 395 320
rect 505 370 595 390
rect 505 320 525 370
rect 575 320 595 370
rect 95 220 115 270
rect 165 220 185 270
rect 95 45 185 220
rect 505 175 595 320
rect 505 125 525 175
rect 575 125 595 175
rect 505 45 595 125
rect 695 370 1230 390
rect 695 320 715 370
rect 765 320 1160 370
rect 1210 320 1230 370
rect 695 300 1230 320
rect 695 175 785 300
rect 695 125 715 175
rect 765 125 785 175
rect 695 105 785 125
rect 915 220 1005 240
rect 915 170 935 220
rect 985 170 1005 220
rect 915 45 1005 170
rect 1140 175 1230 300
rect 1140 125 1160 175
rect 1210 125 1230 175
rect 1140 105 1230 125
rect 1330 355 1420 375
rect 1330 305 1350 355
rect 1400 305 1420 355
rect 1330 175 1420 305
rect 1555 300 1645 470
rect 1745 505 1920 525
rect 1745 455 1765 505
rect 1815 455 1920 505
rect 1745 435 1920 455
rect 1555 250 1575 300
rect 1625 250 1645 300
rect 1555 215 1645 250
rect 1765 300 1855 320
rect 1765 250 1785 300
rect 1835 250 1855 300
rect 1330 125 1350 175
rect 1400 125 1420 175
rect 1330 45 1420 125
rect 1765 200 1855 250
rect 1765 150 1785 200
rect 1835 150 1855 200
rect 1765 45 1855 150
rect 0 -45 1950 45
<< labels >>
flabel metal1 s 1170 1045 1170 1045 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 50 615 50 615 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 206 1415 206 1415 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 1860 465 1860 465 2 FreeSans 400 0 0 0 b
port 2 ne
flabel nwell 10 555 10 555 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 6 5 6 5 2 FreeSans 400 0 0 0 vss
port 4 ne
<< properties >>
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
<< end >>
