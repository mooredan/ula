magic
tech amic5n
timestamp 1626102302
<< nwell >>
rect -130 550 3580 1495
<< ntransistor >>
rect 265 95 325 375
rect 455 95 515 375
rect 645 95 705 375
rect 795 95 855 375
rect 1065 95 1125 375
rect 1215 95 1275 375
rect 1410 95 1470 375
rect 1650 95 1710 375
rect 2170 95 2230 375
rect 2570 95 2630 375
rect 2730 95 2790 375
rect 2935 95 2995 375
rect 3125 95 3185 375
<< ptransistor >>
rect 265 865 325 1345
rect 455 865 515 1345
rect 645 865 705 1345
rect 825 865 885 1345
rect 1065 865 1125 1345
rect 1215 865 1275 1345
rect 1410 865 1470 1345
rect 1650 865 1710 1345
rect 2170 865 2230 1345
rect 2570 865 2630 1345
rect 2730 865 2790 1345
rect 2935 865 2995 1345
rect 3125 865 3185 1345
<< nselect >>
rect 10 835 145 1440
rect 1905 835 2040 1440
rect 3305 835 3440 1440
rect -10 320 1905 430
rect 145 45 1905 320
rect 245 0 1905 45
rect 2050 320 3460 430
rect 2050 0 3305 320
<< pselect >>
rect 145 835 1905 1440
rect 2040 835 3305 1440
rect 10 45 145 320
rect 1905 0 2050 430
rect 3305 0 3440 320
<< ndiffusion >>
rect 145 345 265 375
rect 145 295 175 345
rect 225 295 265 345
rect 145 175 265 295
rect 145 125 175 175
rect 225 125 265 175
rect 145 95 265 125
rect 325 345 455 375
rect 325 295 365 345
rect 415 295 455 345
rect 325 175 455 295
rect 325 125 365 175
rect 415 125 455 175
rect 325 95 455 125
rect 515 345 645 375
rect 515 295 555 345
rect 605 295 645 345
rect 515 175 645 295
rect 515 125 555 175
rect 605 125 645 175
rect 515 95 645 125
rect 705 95 795 375
rect 855 345 1065 375
rect 855 295 950 345
rect 1000 295 1065 345
rect 855 200 1065 295
rect 855 150 950 200
rect 1000 150 1065 200
rect 855 95 1065 150
rect 1125 95 1215 375
rect 1275 345 1410 375
rect 1275 295 1320 345
rect 1370 295 1410 345
rect 1275 175 1410 295
rect 1275 125 1320 175
rect 1370 125 1410 175
rect 1275 95 1410 125
rect 1470 345 1650 375
rect 1470 295 1535 345
rect 1585 295 1650 345
rect 1470 175 1650 295
rect 1470 125 1535 175
rect 1585 125 1650 175
rect 1470 95 1650 125
rect 1710 345 1830 375
rect 1710 295 1750 345
rect 1800 295 1830 345
rect 1710 175 1830 295
rect 1710 125 1750 175
rect 1800 125 1830 175
rect 1710 95 1830 125
rect 2050 345 2170 375
rect 2050 295 2080 345
rect 2130 295 2170 345
rect 2050 175 2170 295
rect 2050 125 2080 175
rect 2130 125 2170 175
rect 2050 95 2170 125
rect 2230 345 2360 375
rect 2230 295 2280 345
rect 2330 295 2360 345
rect 2230 175 2360 295
rect 2230 125 2280 175
rect 2330 125 2360 175
rect 2230 95 2360 125
rect 2450 345 2570 375
rect 2450 295 2480 345
rect 2530 295 2570 345
rect 2450 95 2570 295
rect 2630 95 2730 375
rect 2790 345 2935 375
rect 2790 295 2845 345
rect 2895 295 2935 345
rect 2790 175 2935 295
rect 2790 125 2845 175
rect 2895 125 2935 175
rect 2790 95 2935 125
rect 2995 345 3125 375
rect 2995 295 3035 345
rect 3085 295 3125 345
rect 2995 175 3125 295
rect 2995 125 3035 175
rect 3085 125 3125 175
rect 2995 95 3125 125
rect 3185 345 3305 375
rect 3185 295 3225 345
rect 3275 295 3305 345
rect 3185 175 3305 295
rect 3185 125 3225 175
rect 3275 125 3305 175
rect 3185 95 3305 125
<< pdiffusion >>
rect 145 1315 265 1345
rect 145 1265 175 1315
rect 225 1265 265 1315
rect 145 1195 265 1265
rect 145 1145 175 1195
rect 225 1145 265 1195
rect 145 1070 265 1145
rect 145 1020 175 1070
rect 225 1020 265 1070
rect 145 945 265 1020
rect 145 895 175 945
rect 225 895 265 945
rect 145 865 265 895
rect 325 1315 455 1345
rect 325 1265 365 1315
rect 415 1265 455 1315
rect 325 1195 455 1265
rect 325 1145 365 1195
rect 415 1145 455 1195
rect 325 1070 455 1145
rect 325 1020 365 1070
rect 415 1020 455 1070
rect 325 945 455 1020
rect 325 895 365 945
rect 415 895 455 945
rect 325 865 455 895
rect 515 1315 645 1345
rect 515 1265 555 1315
rect 605 1265 645 1315
rect 515 1200 645 1265
rect 515 1150 555 1200
rect 605 1150 645 1200
rect 515 1085 645 1150
rect 515 1035 555 1085
rect 605 1035 645 1085
rect 515 975 645 1035
rect 515 925 555 975
rect 605 925 645 975
rect 515 865 645 925
rect 705 865 825 1345
rect 885 1315 1065 1345
rect 885 1265 945 1315
rect 995 1265 1065 1315
rect 885 1195 1065 1265
rect 885 1145 945 1195
rect 995 1145 1065 1195
rect 885 1080 1065 1145
rect 885 1030 945 1080
rect 995 1030 1065 1080
rect 885 945 1065 1030
rect 885 895 945 945
rect 995 895 1065 945
rect 885 865 1065 895
rect 1125 865 1215 1345
rect 1275 1315 1410 1345
rect 1275 1265 1320 1315
rect 1370 1265 1410 1315
rect 1275 1200 1410 1265
rect 1275 1150 1320 1200
rect 1370 1150 1410 1200
rect 1275 1085 1410 1150
rect 1275 1035 1320 1085
rect 1370 1035 1410 1085
rect 1275 975 1410 1035
rect 1275 925 1320 975
rect 1370 925 1410 975
rect 1275 865 1410 925
rect 1470 1315 1650 1345
rect 1470 1265 1535 1315
rect 1585 1265 1650 1315
rect 1470 1195 1650 1265
rect 1470 1145 1535 1195
rect 1585 1145 1650 1195
rect 1470 1070 1650 1145
rect 1470 1020 1535 1070
rect 1585 1020 1650 1070
rect 1470 945 1650 1020
rect 1470 895 1535 945
rect 1585 895 1650 945
rect 1470 865 1650 895
rect 1710 1315 1830 1345
rect 1710 1265 1750 1315
rect 1800 1265 1830 1315
rect 1710 1195 1830 1265
rect 1710 1145 1750 1195
rect 1800 1145 1830 1195
rect 1710 1070 1830 1145
rect 1710 1020 1750 1070
rect 1800 1020 1830 1070
rect 1710 945 1830 1020
rect 1710 895 1750 945
rect 1800 895 1830 945
rect 1710 865 1830 895
rect 2040 1315 2170 1345
rect 2040 1265 2080 1315
rect 2130 1265 2170 1315
rect 2040 1200 2170 1265
rect 2040 1150 2080 1200
rect 2130 1150 2170 1200
rect 2040 1085 2170 1150
rect 2040 1035 2080 1085
rect 2130 1035 2170 1085
rect 2040 975 2170 1035
rect 2040 925 2080 975
rect 2130 925 2170 975
rect 2040 865 2170 925
rect 2230 1315 2360 1345
rect 2230 1265 2280 1315
rect 2330 1265 2360 1315
rect 2230 1195 2360 1265
rect 2230 1145 2280 1195
rect 2330 1145 2360 1195
rect 2230 1070 2360 1145
rect 2230 1020 2280 1070
rect 2330 1020 2360 1070
rect 2230 945 2360 1020
rect 2230 895 2280 945
rect 2330 895 2360 945
rect 2230 865 2360 895
rect 2450 1315 2570 1345
rect 2450 1265 2480 1315
rect 2530 1265 2570 1315
rect 2450 1195 2570 1265
rect 2450 1145 2480 1195
rect 2530 1145 2570 1195
rect 2450 1070 2570 1145
rect 2450 1020 2480 1070
rect 2530 1020 2570 1070
rect 2450 865 2570 1020
rect 2630 865 2730 1345
rect 2790 1315 2935 1345
rect 2790 1265 2845 1315
rect 2895 1265 2935 1315
rect 2790 1195 2935 1265
rect 2790 1145 2845 1195
rect 2895 1145 2935 1195
rect 2790 1070 2935 1145
rect 2790 1020 2845 1070
rect 2895 1020 2935 1070
rect 2790 945 2935 1020
rect 2790 895 2845 945
rect 2895 895 2935 945
rect 2790 865 2935 895
rect 2995 1315 3125 1345
rect 2995 1265 3035 1315
rect 3085 1265 3125 1315
rect 2995 1195 3125 1265
rect 2995 1145 3035 1195
rect 3085 1145 3125 1195
rect 2995 1070 3125 1145
rect 2995 1020 3035 1070
rect 3085 1020 3125 1070
rect 2995 945 3125 1020
rect 2995 895 3035 945
rect 3085 895 3125 945
rect 2995 865 3125 895
rect 3185 1315 3305 1345
rect 3185 1265 3225 1315
rect 3275 1265 3305 1315
rect 3185 1195 3305 1265
rect 3185 1145 3225 1195
rect 3275 1145 3305 1195
rect 3185 1070 3305 1145
rect 3185 1020 3225 1070
rect 3275 1020 3305 1070
rect 3185 945 3305 1020
rect 3185 895 3225 945
rect 3275 895 3305 945
rect 3185 865 3305 895
<< psubstratepdiff >>
rect 45 290 145 320
rect 45 240 75 290
rect 125 240 145 290
rect 45 175 145 240
rect 45 125 75 175
rect 125 125 145 175
rect 45 95 145 125
rect 1940 345 2050 375
rect 1940 295 1970 345
rect 2020 295 2050 345
rect 1940 175 2050 295
rect 1940 125 1970 175
rect 2020 125 2050 175
rect 1940 95 2050 125
rect 3305 290 3405 320
rect 3305 240 3325 290
rect 3375 240 3405 290
rect 3305 175 3405 240
rect 3305 125 3325 175
rect 3375 125 3405 175
rect 3305 95 3405 125
<< nsubstratendiff >>
rect 45 1315 145 1345
rect 45 1265 75 1315
rect 125 1265 145 1315
rect 45 1195 145 1265
rect 45 1145 75 1195
rect 125 1145 145 1195
rect 45 1070 145 1145
rect 45 1020 75 1070
rect 125 1020 145 1070
rect 45 945 145 1020
rect 45 895 75 945
rect 125 895 145 945
rect 45 865 145 895
rect 1940 1315 2040 1345
rect 1940 1265 1970 1315
rect 2020 1265 2040 1315
rect 1940 1195 2040 1265
rect 1940 1145 1970 1195
rect 2020 1145 2040 1195
rect 1940 1085 2040 1145
rect 1940 1035 1970 1085
rect 2020 1035 2040 1085
rect 1940 985 2040 1035
rect 1940 935 1970 985
rect 2020 935 2040 985
rect 1940 865 2040 935
rect 3305 1315 3405 1345
rect 3305 1265 3325 1315
rect 3375 1265 3405 1315
rect 3305 1195 3405 1265
rect 3305 1145 3325 1195
rect 3375 1145 3405 1195
rect 3305 1070 3405 1145
rect 3305 1020 3325 1070
rect 3375 1020 3405 1070
rect 3305 945 3405 1020
rect 3305 895 3325 945
rect 3375 895 3405 945
rect 3305 865 3405 895
<< nsubstratencontact >>
rect 75 1265 125 1315
rect 75 1145 125 1195
rect 75 1020 125 1070
rect 75 895 125 945
rect 1970 1265 2020 1315
rect 1970 1145 2020 1195
rect 1970 1035 2020 1085
rect 1970 935 2020 985
rect 3325 1265 3375 1315
rect 3325 1145 3375 1195
rect 3325 1020 3375 1070
rect 3325 895 3375 945
<< psubstratepcontact >>
rect 75 240 125 290
rect 75 125 125 175
rect 1970 295 2020 345
rect 1970 125 2020 175
rect 3325 240 3375 290
rect 3325 125 3375 175
<< ndcontact >>
rect 175 295 225 345
rect 175 125 225 175
rect 365 295 415 345
rect 365 125 415 175
rect 555 295 605 345
rect 555 125 605 175
rect 950 295 1000 345
rect 950 150 1000 200
rect 1320 295 1370 345
rect 1320 125 1370 175
rect 1535 295 1585 345
rect 1535 125 1585 175
rect 1750 295 1800 345
rect 1750 125 1800 175
rect 2080 295 2130 345
rect 2080 125 2130 175
rect 2280 295 2330 345
rect 2280 125 2330 175
rect 2480 295 2530 345
rect 2845 295 2895 345
rect 2845 125 2895 175
rect 3035 295 3085 345
rect 3035 125 3085 175
rect 3225 295 3275 345
rect 3225 125 3275 175
<< pdcontact >>
rect 175 1265 225 1315
rect 175 1145 225 1195
rect 175 1020 225 1070
rect 175 895 225 945
rect 365 1265 415 1315
rect 365 1145 415 1195
rect 365 1020 415 1070
rect 365 895 415 945
rect 555 1265 605 1315
rect 555 1150 605 1200
rect 555 1035 605 1085
rect 555 925 605 975
rect 945 1265 995 1315
rect 945 1145 995 1195
rect 945 1030 995 1080
rect 945 895 995 945
rect 1320 1265 1370 1315
rect 1320 1150 1370 1200
rect 1320 1035 1370 1085
rect 1320 925 1370 975
rect 1535 1265 1585 1315
rect 1535 1145 1585 1195
rect 1535 1020 1585 1070
rect 1535 895 1585 945
rect 1750 1265 1800 1315
rect 1750 1145 1800 1195
rect 1750 1020 1800 1070
rect 1750 895 1800 945
rect 2080 1265 2130 1315
rect 2080 1150 2130 1200
rect 2080 1035 2130 1085
rect 2080 925 2130 975
rect 2280 1265 2330 1315
rect 2280 1145 2330 1195
rect 2280 1020 2330 1070
rect 2280 895 2330 945
rect 2480 1265 2530 1315
rect 2480 1145 2530 1195
rect 2480 1020 2530 1070
rect 2845 1265 2895 1315
rect 2845 1145 2895 1195
rect 2845 1020 2895 1070
rect 2845 895 2895 945
rect 3035 1265 3085 1315
rect 3035 1145 3085 1195
rect 3035 1020 3085 1070
rect 3035 895 3085 945
rect 3225 1265 3275 1315
rect 3225 1145 3275 1195
rect 3225 1020 3275 1070
rect 3225 895 3275 945
<< polysilicon >>
rect 265 1345 325 1410
rect 455 1345 515 1410
rect 645 1345 705 1410
rect 825 1345 885 1410
rect 1065 1345 1125 1410
rect 1215 1345 1275 1410
rect 1410 1345 1470 1410
rect 1650 1345 1710 1410
rect 2170 1345 2230 1410
rect 2570 1345 2630 1410
rect 2730 1345 2790 1410
rect 2935 1345 2995 1410
rect 3125 1345 3185 1410
rect 265 845 325 865
rect 455 845 515 865
rect 645 845 705 865
rect 825 845 885 865
rect 265 785 515 845
rect 615 825 705 845
rect 265 525 325 785
rect 615 775 635 825
rect 685 775 705 825
rect 615 755 705 775
rect 765 825 885 845
rect 765 775 785 825
rect 835 775 885 825
rect 765 755 885 775
rect 265 505 585 525
rect 265 455 515 505
rect 565 455 585 505
rect 265 435 585 455
rect 265 375 325 435
rect 455 375 515 435
rect 645 375 705 755
rect 1065 685 1125 865
rect 1050 665 1140 685
rect 1050 655 1070 665
rect 795 615 1070 655
rect 1120 615 1140 665
rect 795 595 1140 615
rect 795 375 855 595
rect 1215 525 1275 865
rect 1410 845 1470 865
rect 1335 825 1470 845
rect 1335 775 1355 825
rect 1405 775 1470 825
rect 1335 755 1470 775
rect 1050 505 1140 525
rect 1050 455 1070 505
rect 1120 455 1140 505
rect 1050 435 1140 455
rect 1200 505 1290 525
rect 1200 455 1220 505
rect 1270 455 1290 505
rect 1200 435 1290 455
rect 1065 375 1125 435
rect 1215 375 1275 435
rect 1410 375 1470 755
rect 1650 685 1710 865
rect 2170 845 2230 865
rect 2080 825 2230 845
rect 2080 775 2100 825
rect 2150 775 2230 825
rect 2080 755 2230 775
rect 2570 845 2630 865
rect 2570 825 2670 845
rect 2570 775 2600 825
rect 2650 775 2670 825
rect 2570 755 2670 775
rect 1635 665 1725 685
rect 1635 615 1655 665
rect 1705 615 1725 665
rect 1635 595 1725 615
rect 1635 505 1725 525
rect 1635 455 1655 505
rect 1705 455 1725 505
rect 1635 435 1725 455
rect 1650 375 1710 435
rect 2170 375 2230 755
rect 2730 685 2790 865
rect 2935 845 2995 865
rect 3125 845 3185 865
rect 2935 785 3185 845
rect 2935 685 2995 785
rect 2570 665 2660 685
rect 2570 615 2590 665
rect 2640 615 2660 665
rect 2570 595 2660 615
rect 2730 665 2995 685
rect 2730 615 2765 665
rect 2815 615 2885 665
rect 2935 615 2995 665
rect 2730 595 2995 615
rect 2570 375 2630 595
rect 2730 375 2790 595
rect 2935 455 2995 595
rect 2935 395 3185 455
rect 2935 375 2995 395
rect 3125 375 3185 395
rect 265 30 325 95
rect 455 30 515 95
rect 645 30 705 95
rect 795 30 855 95
rect 1065 30 1125 95
rect 1215 30 1275 95
rect 1410 30 1470 95
rect 1650 30 1710 95
rect 2170 30 2230 95
rect 2570 30 2630 95
rect 2730 30 2790 95
rect 2935 30 2995 95
rect 3125 30 3185 95
<< polycontact >>
rect 635 775 685 825
rect 785 775 835 825
rect 515 455 565 505
rect 1070 615 1120 665
rect 1355 775 1405 825
rect 1070 455 1120 505
rect 1220 455 1270 505
rect 2100 775 2150 825
rect 2600 775 2650 825
rect 1655 615 1705 665
rect 1655 455 1705 505
rect 2590 615 2640 665
rect 2765 615 2815 665
rect 2885 615 2935 665
<< metal1 >>
rect 0 1395 3450 1485
rect 55 1315 245 1395
rect 55 1265 75 1315
rect 125 1265 175 1315
rect 225 1265 245 1315
rect 55 1195 245 1265
rect 55 1145 75 1195
rect 125 1145 175 1195
rect 225 1145 245 1195
rect 55 1070 245 1145
rect 55 1020 75 1070
rect 125 1020 175 1070
rect 225 1020 245 1070
rect 55 945 245 1020
rect 55 895 75 945
rect 125 895 175 945
rect 225 895 245 945
rect 55 875 245 895
rect 345 1315 435 1335
rect 345 1265 365 1315
rect 415 1265 435 1315
rect 345 1195 435 1265
rect 345 1145 365 1195
rect 415 1145 435 1195
rect 345 1070 435 1145
rect 345 1020 365 1070
rect 415 1020 435 1070
rect 345 945 435 1020
rect 345 895 365 945
rect 415 895 435 945
rect 535 1315 625 1395
rect 535 1265 555 1315
rect 605 1265 625 1315
rect 535 1200 625 1265
rect 535 1150 555 1200
rect 605 1150 625 1200
rect 535 1085 625 1150
rect 535 1035 555 1085
rect 605 1035 625 1085
rect 535 975 625 1035
rect 535 925 555 975
rect 605 925 625 975
rect 535 905 625 925
rect 915 1315 1020 1335
rect 915 1265 945 1315
rect 995 1265 1020 1315
rect 915 1195 1020 1265
rect 915 1145 945 1195
rect 995 1145 1020 1195
rect 915 1080 1020 1145
rect 915 1030 945 1080
rect 995 1030 1020 1080
rect 915 945 1020 1030
rect 345 685 435 895
rect 915 895 945 945
rect 995 895 1020 945
rect 1300 1315 1390 1395
rect 1300 1265 1320 1315
rect 1370 1265 1390 1315
rect 1300 1200 1390 1265
rect 1300 1150 1320 1200
rect 1370 1150 1390 1200
rect 1300 1085 1390 1150
rect 1300 1035 1320 1085
rect 1370 1035 1390 1085
rect 1300 975 1390 1035
rect 1300 925 1320 975
rect 1370 925 1390 975
rect 1300 905 1390 925
rect 1485 1315 1605 1335
rect 1485 1265 1535 1315
rect 1585 1265 1605 1315
rect 1485 1195 1605 1265
rect 1485 1145 1535 1195
rect 1585 1145 1605 1195
rect 1485 1070 1605 1145
rect 1485 1020 1535 1070
rect 1585 1020 1605 1070
rect 1485 945 1605 1020
rect 915 845 1020 895
rect 1485 895 1535 945
rect 1585 895 1605 945
rect 1485 865 1605 895
rect 1730 1330 1830 1335
rect 1730 1315 1865 1330
rect 1730 1265 1750 1315
rect 1800 1265 1865 1315
rect 1730 1195 1865 1265
rect 1730 1145 1750 1195
rect 1800 1145 1865 1195
rect 1730 1070 1865 1145
rect 1730 1020 1750 1070
rect 1800 1020 1865 1070
rect 1730 945 1865 1020
rect 1730 895 1750 945
rect 1800 895 1865 945
rect 1950 1315 2150 1395
rect 1950 1265 1970 1315
rect 2020 1265 2080 1315
rect 2130 1265 2150 1315
rect 1950 1200 2150 1265
rect 1950 1195 2080 1200
rect 1950 1145 1970 1195
rect 2020 1150 2080 1195
rect 2130 1150 2150 1200
rect 2020 1145 2150 1150
rect 1950 1085 2150 1145
rect 1950 1035 1970 1085
rect 2020 1035 2080 1085
rect 2130 1035 2150 1085
rect 1950 985 2150 1035
rect 1950 935 1970 985
rect 2020 975 2150 985
rect 2020 935 2080 975
rect 1950 925 2080 935
rect 2130 925 2150 975
rect 1950 905 2150 925
rect 2260 1315 2360 1335
rect 2260 1265 2280 1315
rect 2330 1265 2360 1315
rect 2260 1195 2360 1265
rect 2260 1145 2280 1195
rect 2330 1145 2360 1195
rect 2260 1070 2360 1145
rect 2260 1020 2280 1070
rect 2330 1020 2360 1070
rect 2260 945 2360 1020
rect 505 825 705 845
rect 505 775 635 825
rect 685 775 705 825
rect 505 755 705 775
rect 765 825 855 845
rect 765 775 785 825
rect 835 775 855 825
rect 345 665 545 685
rect 345 615 365 665
rect 415 615 475 665
rect 525 615 545 665
rect 345 595 545 615
rect 145 345 245 365
rect 145 310 175 345
rect 55 295 175 310
rect 225 295 245 345
rect 55 290 245 295
rect 55 240 75 290
rect 125 240 245 290
rect 55 175 245 240
rect 55 125 75 175
rect 125 125 175 175
rect 225 125 245 175
rect 55 45 245 125
rect 345 345 435 595
rect 765 525 855 775
rect 495 505 855 525
rect 495 455 515 505
rect 565 455 645 505
rect 695 455 785 505
rect 835 455 855 505
rect 495 435 855 455
rect 915 825 1425 845
rect 915 775 1355 825
rect 1405 775 1425 825
rect 915 755 1425 775
rect 915 365 990 755
rect 1485 685 1575 865
rect 1730 845 1865 895
rect 2260 895 2280 945
rect 2330 895 2360 945
rect 1730 825 2170 845
rect 1730 775 1775 825
rect 1825 775 2100 825
rect 2150 775 2170 825
rect 1730 755 2170 775
rect 1050 665 1250 685
rect 1050 615 1070 665
rect 1120 615 1180 665
rect 1230 615 1250 665
rect 1050 595 1250 615
rect 1310 595 1575 685
rect 1635 665 1725 685
rect 1635 615 1655 665
rect 1705 615 1725 665
rect 1635 595 1725 615
rect 1310 525 1400 595
rect 1050 505 1140 525
rect 1050 455 1070 505
rect 1120 455 1140 505
rect 1050 435 1140 455
rect 1200 505 1400 525
rect 1200 455 1220 505
rect 1270 455 1400 505
rect 1200 435 1400 455
rect 1485 375 1575 595
rect 1635 505 1725 525
rect 1635 455 1655 505
rect 1705 455 1725 505
rect 1635 435 1725 455
rect 1785 375 1865 755
rect 345 295 365 345
rect 415 295 435 345
rect 345 175 435 295
rect 345 125 365 175
rect 415 125 435 175
rect 345 105 435 125
rect 535 345 625 365
rect 535 295 555 345
rect 605 295 625 345
rect 535 175 625 295
rect 535 125 555 175
rect 605 125 625 175
rect 535 45 625 125
rect 915 345 1035 365
rect 915 295 950 345
rect 1000 295 1035 345
rect 915 200 1035 295
rect 915 150 950 200
rect 1000 150 1035 200
rect 915 105 1035 150
rect 1300 345 1390 365
rect 1300 295 1320 345
rect 1370 295 1390 345
rect 1300 175 1390 295
rect 1300 125 1320 175
rect 1370 125 1390 175
rect 1300 45 1390 125
rect 1485 345 1605 375
rect 1485 295 1535 345
rect 1585 295 1605 345
rect 1485 175 1605 295
rect 1485 125 1535 175
rect 1585 125 1605 175
rect 1485 105 1605 125
rect 1730 345 1865 375
rect 1730 295 1750 345
rect 1800 295 1865 345
rect 1730 175 1865 295
rect 1730 125 1750 175
rect 1800 125 1865 175
rect 1730 105 1865 125
rect 1950 345 2150 365
rect 1950 295 1970 345
rect 2020 295 2080 345
rect 2130 295 2150 345
rect 1950 175 2150 295
rect 1950 125 1970 175
rect 2020 125 2080 175
rect 2130 125 2150 175
rect 1950 45 2150 125
rect 2260 345 2360 895
rect 2260 295 2280 345
rect 2330 295 2360 345
rect 2260 195 2360 295
rect 2420 1315 2550 1335
rect 2420 1265 2480 1315
rect 2530 1265 2550 1315
rect 2420 1195 2550 1265
rect 2420 1145 2480 1195
rect 2530 1145 2550 1195
rect 2420 1070 2550 1145
rect 2420 1020 2480 1070
rect 2530 1020 2550 1070
rect 2420 925 2550 1020
rect 2825 1315 2915 1395
rect 2825 1265 2845 1315
rect 2895 1265 2915 1315
rect 2825 1195 2915 1265
rect 2825 1145 2845 1195
rect 2895 1145 2915 1195
rect 2825 1070 2915 1145
rect 2825 1020 2845 1070
rect 2895 1020 2915 1070
rect 2825 945 2915 1020
rect 2420 825 2510 925
rect 2825 895 2845 945
rect 2895 895 2915 945
rect 2825 875 2915 895
rect 3015 1315 3105 1335
rect 3015 1265 3035 1315
rect 3085 1265 3105 1315
rect 3015 1195 3105 1265
rect 3015 1145 3035 1195
rect 3085 1145 3105 1195
rect 3015 1070 3105 1145
rect 3015 1020 3035 1070
rect 3085 1020 3105 1070
rect 3015 945 3105 1020
rect 3015 895 3035 945
rect 3085 895 3105 945
rect 2420 775 2440 825
rect 2490 775 2510 825
rect 2420 375 2510 775
rect 2570 825 2670 845
rect 2570 775 2600 825
rect 2650 775 2670 825
rect 2570 755 2670 775
rect 2570 665 2660 685
rect 2570 615 2590 665
rect 2640 615 2660 665
rect 2570 595 2660 615
rect 2730 665 2955 685
rect 2730 615 2765 665
rect 2815 615 2885 665
rect 2935 615 2955 665
rect 2730 595 2955 615
rect 2730 525 2825 595
rect 2610 435 2825 525
rect 2420 345 2550 375
rect 2420 295 2480 345
rect 2530 295 2550 345
rect 2420 275 2550 295
rect 2610 195 2705 435
rect 2260 175 2705 195
rect 2260 125 2280 175
rect 2330 125 2705 175
rect 2260 105 2705 125
rect 2825 345 2915 365
rect 2825 295 2845 345
rect 2895 295 2915 345
rect 2825 175 2915 295
rect 2825 125 2845 175
rect 2895 125 2915 175
rect 2825 45 2915 125
rect 3015 345 3105 895
rect 3205 1315 3395 1395
rect 3205 1265 3225 1315
rect 3275 1265 3325 1315
rect 3375 1265 3395 1315
rect 3205 1195 3395 1265
rect 3205 1145 3225 1195
rect 3275 1145 3325 1195
rect 3375 1145 3395 1195
rect 3205 1070 3395 1145
rect 3205 1020 3225 1070
rect 3275 1020 3325 1070
rect 3375 1020 3395 1070
rect 3205 945 3395 1020
rect 3205 895 3225 945
rect 3275 895 3325 945
rect 3375 895 3395 945
rect 3205 875 3395 895
rect 3015 295 3035 345
rect 3085 295 3105 345
rect 3015 175 3105 295
rect 3015 125 3035 175
rect 3085 125 3105 175
rect 3015 105 3105 125
rect 3205 345 3305 365
rect 3205 295 3225 345
rect 3275 310 3305 345
rect 3275 295 3395 310
rect 3205 290 3395 295
rect 3205 240 3325 290
rect 3375 240 3395 290
rect 3205 175 3395 240
rect 3205 125 3225 175
rect 3275 125 3325 175
rect 3375 125 3395 175
rect 3205 45 3395 125
rect 0 -45 3450 45
<< via1 >>
rect 365 615 415 665
rect 475 615 525 665
rect 515 455 565 505
rect 645 455 695 505
rect 785 455 835 505
rect 1775 775 1825 825
rect 1070 615 1120 665
rect 1180 615 1230 665
rect 1655 615 1705 665
rect 1070 455 1120 505
rect 1655 455 1705 505
rect 2440 775 2490 825
rect 2600 775 2650 825
rect 2590 615 2640 665
<< metal2 >>
rect 1730 825 2510 845
rect 1730 775 1775 825
rect 1825 775 2440 825
rect 2490 775 2510 825
rect 1730 755 2510 775
rect 2580 825 2820 845
rect 2580 775 2600 825
rect 2650 775 2820 825
rect 2580 755 2820 775
rect 345 665 2660 685
rect 345 615 365 665
rect 415 615 475 665
rect 525 615 1070 665
rect 1120 615 1180 665
rect 1230 615 1655 665
rect 1705 615 2590 665
rect 2640 615 2660 665
rect 345 595 2660 615
rect 2730 525 2820 755
rect 495 505 2820 525
rect 495 455 515 505
rect 565 455 645 505
rect 695 455 785 505
rect 835 455 1070 505
rect 1120 455 1655 505
rect 1705 455 2820 505
rect 495 435 2820 455
<< labels >>
flabel ndiffusion s 1155 195 1155 195 2 FreeSans 400 0 0 0 x6
flabel ndiffusion 735 195 735 195 2 FreeSans 400 0 0 0 x5
flabel metal1 360 610 360 610 2 FreeSans 400 0 0 0 nck
flabel metal1 s 515 800 515 800 2 FreeSans 400 0 0 0 d
port 1 s
flabel metal1 s 555 1395 555 1395 2 FreeSans 400 0 0 0 vdd
port 3 n
flabel pdiffusion s 1155 1065 1155 1065 2 FreeSans 400 0 0 0 x2
flabel pdiffusion s 765 1065 765 1065 2 FreeSans 400 0 0 0 x1
flabel metal1 s 1050 465 1050 465 2 FreeSans 400 0 0 0 ck
port 2 ne
flabel metal1 s 945 925 945 925 2 FreeSans 400 0 0 0 nmas
flabel metal1 s 175 15 175 15 2 FreeSans 400 0 0 0 vss
port 4 s
flabel metal1 s 1791 940 1791 940 8 FreeSans 400 180 0 0 slv
flabel metal1 s 1545 1065 1545 1065 2 FreeSans 400 0 0 0 mas
flabel metal1 s 2800 640 2800 640 2 FreeSans 400 0 0 0 nslv
flabel pdiffusion s 2660 1185 2660 1185 2 FreeSans 400 0 0 0 x4
flabel metal1 s 3035 710 3035 710 2 FreeSans 400 0 0 0 q
port 0 e
flabel ndiffusion s 2715 150 2715 150 2 FreeSans 400 0 0 0 x8
<< properties >>
string LEFsite core
string LEFclass CORE
string FIXED_BBOX 0 0 3450 1440
string LEFsymmetry X Y
<< end >>
