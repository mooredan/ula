magic
tech amic5n
timestamp 1622288771
<< metal1 >>
rect 1145 2220 1205 2270
rect 1130 2200 1220 2220
rect 1130 2150 1150 2200
rect 1200 2150 1220 2200
rect 1130 2130 1220 2150
rect 1145 1900 1205 2130
rect 1280 2060 1340 2270
rect 1415 2220 1475 2270
rect 1400 2200 1490 2220
rect 1400 2150 1420 2200
rect 1470 2150 1490 2200
rect 1400 2130 1490 2150
rect 1265 2040 1355 2060
rect 1265 1990 1285 2040
rect 1335 1990 1355 2040
rect 1265 1970 1355 1990
rect 1130 1880 1220 1900
rect 1130 1830 1150 1880
rect 1200 1830 1220 1880
rect 1130 1810 1220 1830
rect 1145 1580 1205 1810
rect 1280 1740 1340 1970
rect 1415 1900 1475 2130
rect 1550 2060 1610 2270
rect 1685 2220 1745 2270
rect 1670 2200 1760 2220
rect 1670 2150 1690 2200
rect 1740 2150 1760 2200
rect 1670 2130 1760 2150
rect 1535 2040 1625 2060
rect 1535 1990 1555 2040
rect 1605 1990 1625 2040
rect 1535 1970 1625 1990
rect 1400 1880 1490 1900
rect 1400 1830 1420 1880
rect 1470 1830 1490 1880
rect 1400 1810 1490 1830
rect 1265 1720 1355 1740
rect 1265 1670 1285 1720
rect 1335 1670 1355 1720
rect 1265 1650 1355 1670
rect 1130 1560 1220 1580
rect 1130 1510 1150 1560
rect 1200 1510 1220 1560
rect 1130 1490 1220 1510
rect 1145 1260 1205 1490
rect 1280 1420 1340 1650
rect 1415 1580 1475 1810
rect 1550 1740 1610 1970
rect 1685 1900 1745 2130
rect 1820 2060 1880 2270
rect 1955 2220 2015 2270
rect 1940 2200 2030 2220
rect 1940 2150 1960 2200
rect 2010 2150 2030 2200
rect 1940 2130 2030 2150
rect 1805 2040 1895 2060
rect 1805 1990 1825 2040
rect 1875 1990 1895 2040
rect 1805 1970 1895 1990
rect 1670 1880 1760 1900
rect 1670 1830 1690 1880
rect 1740 1830 1760 1880
rect 1670 1810 1760 1830
rect 1535 1720 1625 1740
rect 1535 1670 1555 1720
rect 1605 1670 1625 1720
rect 1535 1650 1625 1670
rect 1400 1560 1490 1580
rect 1400 1510 1420 1560
rect 1470 1510 1490 1560
rect 1400 1490 1490 1510
rect 1265 1400 1355 1420
rect 1265 1350 1285 1400
rect 1335 1350 1355 1400
rect 1265 1330 1355 1350
rect 1130 1240 1220 1260
rect 1130 1190 1150 1240
rect 1200 1190 1220 1240
rect 1130 1170 1220 1190
rect 1145 940 1205 1170
rect 1280 1100 1340 1330
rect 1415 1260 1475 1490
rect 1550 1420 1610 1650
rect 1685 1580 1745 1810
rect 1820 1740 1880 1970
rect 1955 1900 2015 2130
rect 2090 2060 2150 2270
rect 2225 2220 2285 2270
rect 2210 2200 2300 2220
rect 2210 2150 2230 2200
rect 2280 2150 2300 2200
rect 2210 2130 2300 2150
rect 2075 2040 2165 2060
rect 2075 1990 2095 2040
rect 2145 1990 2165 2040
rect 2075 1970 2165 1990
rect 1940 1880 2030 1900
rect 1940 1830 1960 1880
rect 2010 1830 2030 1880
rect 1940 1810 2030 1830
rect 1805 1720 1895 1740
rect 1805 1670 1825 1720
rect 1875 1670 1895 1720
rect 1805 1650 1895 1670
rect 1670 1560 1760 1580
rect 1670 1510 1690 1560
rect 1740 1510 1760 1560
rect 1670 1490 1760 1510
rect 1535 1400 1625 1420
rect 1535 1350 1555 1400
rect 1605 1350 1625 1400
rect 1535 1330 1625 1350
rect 1400 1240 1490 1260
rect 1400 1190 1420 1240
rect 1470 1190 1490 1240
rect 1400 1170 1490 1190
rect 1265 1080 1355 1100
rect 1265 1030 1285 1080
rect 1335 1030 1355 1080
rect 1265 1010 1355 1030
rect 1130 920 1220 940
rect 1130 870 1150 920
rect 1200 870 1220 920
rect 1130 850 1220 870
rect 1145 620 1205 850
rect 1280 780 1340 1010
rect 1415 940 1475 1170
rect 1550 1100 1610 1330
rect 1685 1260 1745 1490
rect 1820 1420 1880 1650
rect 1955 1580 2015 1810
rect 2090 1740 2150 1970
rect 2225 1900 2285 2130
rect 2360 2060 2420 2270
rect 2495 2220 2555 2270
rect 2480 2200 2570 2220
rect 2480 2150 2500 2200
rect 2550 2150 2570 2200
rect 2480 2130 2570 2150
rect 2345 2040 2435 2060
rect 2345 1990 2365 2040
rect 2415 1990 2435 2040
rect 2345 1970 2435 1990
rect 2210 1880 2300 1900
rect 2210 1830 2230 1880
rect 2280 1830 2300 1880
rect 2210 1810 2300 1830
rect 2075 1720 2165 1740
rect 2075 1670 2095 1720
rect 2145 1670 2165 1720
rect 2075 1650 2165 1670
rect 1940 1560 2030 1580
rect 1940 1510 1960 1560
rect 2010 1510 2030 1560
rect 1940 1490 2030 1510
rect 1805 1400 1895 1420
rect 1805 1350 1825 1400
rect 1875 1350 1895 1400
rect 1805 1330 1895 1350
rect 1670 1240 1760 1260
rect 1670 1190 1690 1240
rect 1740 1190 1760 1240
rect 1670 1170 1760 1190
rect 1535 1080 1625 1100
rect 1535 1030 1555 1080
rect 1605 1030 1625 1080
rect 1535 1010 1625 1030
rect 1400 920 1490 940
rect 1400 870 1420 920
rect 1470 870 1490 920
rect 1400 850 1490 870
rect 1265 760 1355 780
rect 1265 710 1285 760
rect 1335 710 1355 760
rect 1265 690 1355 710
rect 1130 600 1220 620
rect 1130 550 1150 600
rect 1200 550 1220 600
rect 1130 530 1220 550
rect 1145 300 1205 530
rect 1280 460 1340 690
rect 1415 620 1475 850
rect 1550 780 1610 1010
rect 1685 940 1745 1170
rect 1820 1100 1880 1330
rect 1955 1260 2015 1490
rect 2090 1420 2150 1650
rect 2225 1580 2285 1810
rect 2360 1740 2420 1970
rect 2495 1900 2555 2130
rect 2630 2060 2690 2270
rect 2765 2220 2825 2270
rect 2750 2200 2840 2220
rect 2750 2150 2770 2200
rect 2820 2150 2840 2200
rect 2750 2130 2840 2150
rect 2615 2040 2705 2060
rect 2615 1990 2635 2040
rect 2685 1990 2705 2040
rect 2615 1970 2705 1990
rect 2480 1880 2570 1900
rect 2480 1830 2500 1880
rect 2550 1830 2570 1880
rect 2480 1810 2570 1830
rect 2345 1720 2435 1740
rect 2345 1670 2365 1720
rect 2415 1670 2435 1720
rect 2345 1650 2435 1670
rect 2210 1560 2300 1580
rect 2210 1510 2230 1560
rect 2280 1510 2300 1560
rect 2210 1490 2300 1510
rect 2075 1400 2165 1420
rect 2075 1350 2095 1400
rect 2145 1350 2165 1400
rect 2075 1330 2165 1350
rect 1940 1240 2030 1260
rect 1940 1190 1960 1240
rect 2010 1190 2030 1240
rect 1940 1170 2030 1190
rect 1805 1080 1895 1100
rect 1805 1030 1825 1080
rect 1875 1030 1895 1080
rect 1805 1010 1895 1030
rect 1670 920 1760 940
rect 1670 870 1690 920
rect 1740 870 1760 920
rect 1670 850 1760 870
rect 1535 760 1625 780
rect 1535 710 1555 760
rect 1605 710 1625 760
rect 1535 690 1625 710
rect 1400 600 1490 620
rect 1400 550 1420 600
rect 1470 550 1490 600
rect 1400 530 1490 550
rect 1265 440 1355 460
rect 1265 390 1285 440
rect 1335 390 1355 440
rect 1265 370 1355 390
rect 1130 280 1220 300
rect 1130 230 1150 280
rect 1200 230 1220 280
rect 1130 210 1220 230
rect 1145 -20 1205 210
rect 1280 140 1340 370
rect 1415 300 1475 530
rect 1550 460 1610 690
rect 1685 620 1745 850
rect 1820 780 1880 1010
rect 1955 940 2015 1170
rect 2090 1100 2150 1330
rect 2225 1260 2285 1490
rect 2360 1420 2420 1650
rect 2495 1580 2555 1810
rect 2630 1740 2690 1970
rect 2765 1900 2825 2130
rect 2900 2060 2960 2270
rect 3035 2220 3095 2275
rect 3020 2200 3110 2220
rect 3020 2150 3040 2200
rect 3090 2150 3110 2200
rect 3020 2130 3110 2150
rect 2885 2040 2975 2060
rect 2885 1990 2905 2040
rect 2955 1990 2975 2040
rect 2885 1970 2975 1990
rect 2750 1880 2840 1900
rect 2750 1830 2770 1880
rect 2820 1830 2840 1880
rect 2750 1810 2840 1830
rect 2615 1720 2705 1740
rect 2615 1670 2635 1720
rect 2685 1670 2705 1720
rect 2615 1650 2705 1670
rect 2480 1560 2570 1580
rect 2480 1510 2500 1560
rect 2550 1510 2570 1560
rect 2480 1490 2570 1510
rect 2345 1400 2435 1420
rect 2345 1350 2365 1400
rect 2415 1350 2435 1400
rect 2345 1330 2435 1350
rect 2210 1240 2300 1260
rect 2210 1190 2230 1240
rect 2280 1190 2300 1240
rect 2210 1170 2300 1190
rect 2075 1080 2165 1100
rect 2075 1030 2095 1080
rect 2145 1030 2165 1080
rect 2075 1010 2165 1030
rect 1940 920 2030 940
rect 1940 870 1960 920
rect 2010 870 2030 920
rect 1940 850 2030 870
rect 1805 760 1895 780
rect 1805 710 1825 760
rect 1875 710 1895 760
rect 1805 690 1895 710
rect 1670 600 1760 620
rect 1670 550 1690 600
rect 1740 550 1760 600
rect 1670 530 1760 550
rect 1535 440 1625 460
rect 1535 390 1555 440
rect 1605 390 1625 440
rect 1535 370 1625 390
rect 1400 280 1490 300
rect 1400 230 1420 280
rect 1470 230 1490 280
rect 1400 210 1490 230
rect 1265 120 1355 140
rect 1265 70 1285 120
rect 1335 70 1355 120
rect 1265 50 1355 70
rect 1130 -40 1220 -20
rect 1130 -90 1150 -40
rect 1200 -90 1220 -40
rect 1130 -110 1220 -90
rect 1145 -265 1205 -110
rect 1280 -265 1340 50
rect 1415 -20 1475 210
rect 1550 140 1610 370
rect 1685 300 1745 530
rect 1820 460 1880 690
rect 1955 620 2015 850
rect 2090 780 2150 1010
rect 2225 940 2285 1170
rect 2360 1100 2420 1330
rect 2495 1260 2555 1490
rect 2630 1420 2690 1650
rect 2765 1580 2825 1810
rect 2900 1740 2960 1970
rect 3035 1900 3095 2130
rect 3020 1880 3110 1900
rect 3020 1830 3040 1880
rect 3090 1830 3110 1880
rect 3020 1810 3110 1830
rect 2885 1720 2975 1740
rect 2885 1670 2905 1720
rect 2955 1670 2975 1720
rect 2885 1650 2975 1670
rect 2750 1560 2840 1580
rect 2750 1510 2770 1560
rect 2820 1510 2840 1560
rect 2750 1490 2840 1510
rect 2615 1400 2705 1420
rect 2615 1350 2635 1400
rect 2685 1350 2705 1400
rect 2615 1330 2705 1350
rect 2480 1240 2570 1260
rect 2480 1190 2500 1240
rect 2550 1190 2570 1240
rect 2480 1170 2570 1190
rect 2345 1080 2435 1100
rect 2345 1030 2365 1080
rect 2415 1030 2435 1080
rect 2345 1010 2435 1030
rect 2210 920 2300 940
rect 2210 870 2230 920
rect 2280 870 2300 920
rect 2210 850 2300 870
rect 2075 760 2165 780
rect 2075 710 2095 760
rect 2145 710 2165 760
rect 2075 690 2165 710
rect 1940 600 2030 620
rect 1940 550 1960 600
rect 2010 550 2030 600
rect 1940 530 2030 550
rect 1805 440 1895 460
rect 1805 390 1825 440
rect 1875 390 1895 440
rect 1805 370 1895 390
rect 1670 280 1760 300
rect 1670 230 1690 280
rect 1740 230 1760 280
rect 1670 210 1760 230
rect 1535 120 1625 140
rect 1535 70 1555 120
rect 1605 70 1625 120
rect 1535 50 1625 70
rect 1400 -40 1490 -20
rect 1400 -90 1420 -40
rect 1470 -90 1490 -40
rect 1400 -110 1490 -90
rect 1415 -265 1475 -110
rect 1550 -265 1610 50
rect 1685 -20 1745 210
rect 1820 140 1880 370
rect 1955 300 2015 530
rect 2090 460 2150 690
rect 2225 620 2285 850
rect 2360 780 2420 1010
rect 2495 940 2555 1170
rect 2630 1100 2690 1330
rect 2765 1260 2825 1490
rect 2900 1420 2960 1650
rect 3035 1580 3095 1810
rect 3020 1560 3110 1580
rect 3020 1510 3040 1560
rect 3090 1510 3110 1560
rect 3020 1490 3110 1510
rect 2885 1400 2975 1420
rect 2885 1350 2905 1400
rect 2955 1350 2975 1400
rect 2885 1330 2975 1350
rect 2750 1240 2840 1260
rect 2750 1190 2770 1240
rect 2820 1190 2840 1240
rect 2750 1170 2840 1190
rect 2615 1080 2705 1100
rect 2615 1030 2635 1080
rect 2685 1030 2705 1080
rect 2615 1010 2705 1030
rect 2480 920 2570 940
rect 2480 870 2500 920
rect 2550 870 2570 920
rect 2480 850 2570 870
rect 2345 760 2435 780
rect 2345 710 2365 760
rect 2415 710 2435 760
rect 2345 690 2435 710
rect 2210 600 2300 620
rect 2210 550 2230 600
rect 2280 550 2300 600
rect 2210 530 2300 550
rect 2075 440 2165 460
rect 2075 390 2095 440
rect 2145 390 2165 440
rect 2075 370 2165 390
rect 1940 280 2030 300
rect 1940 230 1960 280
rect 2010 230 2030 280
rect 1940 210 2030 230
rect 1805 120 1895 140
rect 1805 70 1825 120
rect 1875 70 1895 120
rect 1805 50 1895 70
rect 1670 -40 1760 -20
rect 1670 -90 1690 -40
rect 1740 -90 1760 -40
rect 1670 -110 1760 -90
rect 1685 -265 1745 -110
rect 1820 -265 1880 50
rect 1955 -20 2015 210
rect 2090 140 2150 370
rect 2225 300 2285 530
rect 2360 460 2420 690
rect 2495 620 2555 850
rect 2630 780 2690 1010
rect 2765 940 2825 1170
rect 2900 1100 2960 1330
rect 3035 1260 3095 1490
rect 3020 1240 3110 1260
rect 3020 1190 3040 1240
rect 3090 1190 3110 1240
rect 3020 1170 3110 1190
rect 2885 1080 2975 1100
rect 2885 1030 2905 1080
rect 2955 1030 2975 1080
rect 2885 1010 2975 1030
rect 2750 920 2840 940
rect 2750 870 2770 920
rect 2820 870 2840 920
rect 2750 850 2840 870
rect 2615 760 2705 780
rect 2615 710 2635 760
rect 2685 710 2705 760
rect 2615 690 2705 710
rect 2480 600 2570 620
rect 2480 550 2500 600
rect 2550 550 2570 600
rect 2480 530 2570 550
rect 2345 440 2435 460
rect 2345 390 2365 440
rect 2415 390 2435 440
rect 2345 370 2435 390
rect 2210 280 2300 300
rect 2210 230 2230 280
rect 2280 230 2300 280
rect 2210 210 2300 230
rect 2075 120 2165 140
rect 2075 70 2095 120
rect 2145 70 2165 120
rect 2075 50 2165 70
rect 1940 -40 2030 -20
rect 1940 -90 1960 -40
rect 2010 -90 2030 -40
rect 1940 -110 2030 -90
rect 1955 -265 2015 -110
rect 2090 -265 2150 50
rect 2225 -20 2285 210
rect 2360 140 2420 370
rect 2495 300 2555 530
rect 2630 460 2690 690
rect 2765 620 2825 850
rect 2900 780 2960 1010
rect 3035 940 3095 1170
rect 3020 920 3110 940
rect 3020 870 3040 920
rect 3090 870 3110 920
rect 3020 850 3110 870
rect 2885 760 2975 780
rect 2885 710 2905 760
rect 2955 710 2975 760
rect 2885 690 2975 710
rect 2750 600 2840 620
rect 2750 550 2770 600
rect 2820 550 2840 600
rect 2750 530 2840 550
rect 2615 440 2705 460
rect 2615 390 2635 440
rect 2685 390 2705 440
rect 2615 370 2705 390
rect 2480 280 2570 300
rect 2480 230 2500 280
rect 2550 230 2570 280
rect 2480 210 2570 230
rect 2345 120 2435 140
rect 2345 70 2365 120
rect 2415 70 2435 120
rect 2345 50 2435 70
rect 2210 -40 2300 -20
rect 2210 -90 2230 -40
rect 2280 -90 2300 -40
rect 2210 -110 2300 -90
rect 2225 -265 2285 -110
rect 2360 -265 2420 50
rect 2495 -20 2555 210
rect 2630 140 2690 370
rect 2765 300 2825 530
rect 2900 460 2960 690
rect 3035 620 3095 850
rect 3020 600 3110 620
rect 3020 550 3040 600
rect 3090 550 3110 600
rect 3020 530 3110 550
rect 2885 440 2975 460
rect 2885 390 2905 440
rect 2955 390 2975 440
rect 2885 370 2975 390
rect 2750 280 2840 300
rect 2750 230 2770 280
rect 2820 230 2840 280
rect 2750 210 2840 230
rect 2615 120 2705 140
rect 2615 70 2635 120
rect 2685 70 2705 120
rect 2615 50 2705 70
rect 2480 -40 2570 -20
rect 2480 -90 2500 -40
rect 2550 -90 2570 -40
rect 2480 -110 2570 -90
rect 2495 -265 2555 -110
rect 2630 -265 2690 50
rect 2765 -20 2825 210
rect 2900 140 2960 370
rect 3035 300 3095 530
rect 3020 280 3110 300
rect 3020 230 3040 280
rect 3090 230 3110 280
rect 3020 210 3110 230
rect 3885 215 3945 515
rect 4020 485 4080 515
rect 4005 465 4095 485
rect 4005 415 4025 465
rect 4075 415 4095 465
rect 4005 395 4095 415
rect 4020 325 4080 395
rect 4005 305 4095 325
rect 4005 255 4025 305
rect 4075 255 4095 305
rect 4005 235 4095 255
rect 4020 215 4080 235
rect 4155 215 4215 515
rect 2885 120 2975 140
rect 2885 70 2905 120
rect 2955 70 2975 120
rect 2885 50 2975 70
rect 2750 -40 2840 -20
rect 2750 -90 2770 -40
rect 2820 -90 2840 -40
rect 2750 -110 2840 -90
rect 2765 -265 2825 -110
rect 2900 -265 2960 50
rect 3035 -20 3095 210
rect 3020 -40 3110 -20
rect 3020 -90 3040 -40
rect 3090 -90 3110 -40
rect 3020 -110 3110 -90
rect 3035 -265 3095 -110
<< via1 >>
rect 1150 2150 1200 2200
rect 1420 2150 1470 2200
rect 1285 1990 1335 2040
rect 1150 1830 1200 1880
rect 1690 2150 1740 2200
rect 1555 1990 1605 2040
rect 1420 1830 1470 1880
rect 1285 1670 1335 1720
rect 1150 1510 1200 1560
rect 1960 2150 2010 2200
rect 1825 1990 1875 2040
rect 1690 1830 1740 1880
rect 1555 1670 1605 1720
rect 1420 1510 1470 1560
rect 1285 1350 1335 1400
rect 1150 1190 1200 1240
rect 2230 2150 2280 2200
rect 2095 1990 2145 2040
rect 1960 1830 2010 1880
rect 1825 1670 1875 1720
rect 1690 1510 1740 1560
rect 1555 1350 1605 1400
rect 1420 1190 1470 1240
rect 1285 1030 1335 1080
rect 1150 870 1200 920
rect 2500 2150 2550 2200
rect 2365 1990 2415 2040
rect 2230 1830 2280 1880
rect 2095 1670 2145 1720
rect 1960 1510 2010 1560
rect 1825 1350 1875 1400
rect 1690 1190 1740 1240
rect 1555 1030 1605 1080
rect 1420 870 1470 920
rect 1285 710 1335 760
rect 1150 550 1200 600
rect 2770 2150 2820 2200
rect 2635 1990 2685 2040
rect 2500 1830 2550 1880
rect 2365 1670 2415 1720
rect 2230 1510 2280 1560
rect 2095 1350 2145 1400
rect 1960 1190 2010 1240
rect 1825 1030 1875 1080
rect 1690 870 1740 920
rect 1555 710 1605 760
rect 1420 550 1470 600
rect 1285 390 1335 440
rect 1150 230 1200 280
rect 3040 2150 3090 2200
rect 2905 1990 2955 2040
rect 2770 1830 2820 1880
rect 2635 1670 2685 1720
rect 2500 1510 2550 1560
rect 2365 1350 2415 1400
rect 2230 1190 2280 1240
rect 2095 1030 2145 1080
rect 1960 870 2010 920
rect 1825 710 1875 760
rect 1690 550 1740 600
rect 1555 390 1605 440
rect 1420 230 1470 280
rect 1285 70 1335 120
rect 1150 -90 1200 -40
rect 3040 1830 3090 1880
rect 2905 1670 2955 1720
rect 2770 1510 2820 1560
rect 2635 1350 2685 1400
rect 2500 1190 2550 1240
rect 2365 1030 2415 1080
rect 2230 870 2280 920
rect 2095 710 2145 760
rect 1960 550 2010 600
rect 1825 390 1875 440
rect 1690 230 1740 280
rect 1555 70 1605 120
rect 1420 -90 1470 -40
rect 3040 1510 3090 1560
rect 2905 1350 2955 1400
rect 2770 1190 2820 1240
rect 2635 1030 2685 1080
rect 2500 870 2550 920
rect 2365 710 2415 760
rect 2230 550 2280 600
rect 2095 390 2145 440
rect 1960 230 2010 280
rect 1825 70 1875 120
rect 1690 -90 1740 -40
rect 3040 1190 3090 1240
rect 2905 1030 2955 1080
rect 2770 870 2820 920
rect 2635 710 2685 760
rect 2500 550 2550 600
rect 2365 390 2415 440
rect 2230 230 2280 280
rect 2095 70 2145 120
rect 1960 -90 2010 -40
rect 3040 870 3090 920
rect 2905 710 2955 760
rect 2770 550 2820 600
rect 2635 390 2685 440
rect 2500 230 2550 280
rect 2365 70 2415 120
rect 2230 -90 2280 -40
rect 3040 550 3090 600
rect 2905 390 2955 440
rect 2770 230 2820 280
rect 2635 70 2685 120
rect 2500 -90 2550 -40
rect 3040 230 3090 280
rect 4025 415 4075 465
rect 4025 255 4075 305
rect 2905 70 2955 120
rect 2770 -90 2820 -40
rect 3040 -90 3090 -40
<< metal2 >>
rect 1130 2210 1220 2220
rect 1400 2210 1490 2220
rect 1670 2210 1760 2220
rect 1940 2210 2030 2220
rect 2210 2210 2300 2220
rect 2480 2210 2570 2220
rect 2750 2210 2840 2220
rect 3020 2210 3110 2220
rect 1085 2200 3220 2210
rect 1085 2150 1150 2200
rect 1200 2150 1420 2200
rect 1470 2150 1690 2200
rect 1740 2150 1960 2200
rect 2010 2150 2230 2200
rect 2280 2150 2500 2200
rect 2550 2150 2770 2200
rect 2820 2150 3040 2200
rect 3090 2150 3220 2200
rect 1085 2140 3220 2150
rect 1130 2130 1220 2140
rect 1400 2130 1490 2140
rect 1670 2130 1760 2140
rect 1940 2130 2030 2140
rect 2210 2130 2300 2140
rect 2480 2130 2570 2140
rect 2750 2130 2840 2140
rect 3020 2130 3110 2140
rect 1265 2050 1355 2060
rect 1535 2050 1625 2060
rect 1805 2050 1895 2060
rect 2075 2050 2165 2060
rect 2345 2050 2435 2060
rect 2615 2050 2705 2060
rect 2885 2050 2975 2060
rect 1085 2040 3215 2050
rect 1085 1990 1285 2040
rect 1335 1990 1555 2040
rect 1605 1990 1825 2040
rect 1875 1990 2095 2040
rect 2145 1990 2365 2040
rect 2415 1990 2635 2040
rect 2685 1990 2905 2040
rect 2955 1990 3215 2040
rect 1085 1980 3215 1990
rect 1265 1970 1355 1980
rect 1535 1970 1625 1980
rect 1805 1970 1895 1980
rect 2075 1970 2165 1980
rect 2345 1970 2435 1980
rect 2615 1970 2705 1980
rect 2885 1970 2975 1980
rect 1130 1890 1220 1900
rect 1400 1890 1490 1900
rect 1670 1890 1760 1900
rect 1940 1890 2030 1900
rect 2210 1890 2300 1900
rect 2480 1890 2570 1900
rect 2750 1890 2840 1900
rect 3020 1890 3110 1900
rect 1085 1880 3220 1890
rect 1085 1830 1150 1880
rect 1200 1830 1420 1880
rect 1470 1830 1690 1880
rect 1740 1830 1960 1880
rect 2010 1830 2230 1880
rect 2280 1830 2500 1880
rect 2550 1830 2770 1880
rect 2820 1830 3040 1880
rect 3090 1830 3220 1880
rect 1085 1820 3220 1830
rect 1130 1810 1220 1820
rect 1400 1810 1490 1820
rect 1670 1810 1760 1820
rect 1940 1810 2030 1820
rect 2210 1810 2300 1820
rect 2480 1810 2570 1820
rect 2750 1810 2840 1820
rect 3020 1810 3110 1820
rect 1265 1730 1355 1740
rect 1535 1730 1625 1740
rect 1805 1730 1895 1740
rect 2075 1730 2165 1740
rect 2345 1730 2435 1740
rect 2615 1730 2705 1740
rect 2885 1730 2975 1740
rect 1085 1720 3215 1730
rect 1085 1670 1285 1720
rect 1335 1670 1555 1720
rect 1605 1670 1825 1720
rect 1875 1670 2095 1720
rect 2145 1670 2365 1720
rect 2415 1670 2635 1720
rect 2685 1670 2905 1720
rect 2955 1670 3215 1720
rect 1085 1660 3215 1670
rect 1265 1650 1355 1660
rect 1535 1650 1625 1660
rect 1805 1650 1895 1660
rect 2075 1650 2165 1660
rect 2345 1650 2435 1660
rect 2615 1650 2705 1660
rect 2885 1650 2975 1660
rect 1130 1570 1220 1580
rect 1400 1570 1490 1580
rect 1670 1570 1760 1580
rect 1940 1570 2030 1580
rect 2210 1570 2300 1580
rect 2480 1570 2570 1580
rect 2750 1570 2840 1580
rect 3020 1570 3110 1580
rect 1085 1560 3220 1570
rect 1085 1510 1150 1560
rect 1200 1510 1420 1560
rect 1470 1510 1690 1560
rect 1740 1510 1960 1560
rect 2010 1510 2230 1560
rect 2280 1510 2500 1560
rect 2550 1510 2770 1560
rect 2820 1510 3040 1560
rect 3090 1510 3220 1560
rect 1085 1500 3220 1510
rect 1130 1490 1220 1500
rect 1400 1490 1490 1500
rect 1670 1490 1760 1500
rect 1940 1490 2030 1500
rect 2210 1490 2300 1500
rect 2480 1490 2570 1500
rect 2750 1490 2840 1500
rect 3020 1490 3110 1500
rect -210 1410 -120 1420
rect 100 1410 190 1420
rect 410 1410 500 1420
rect 720 1410 810 1420
rect 1265 1410 1355 1420
rect 1535 1410 1625 1420
rect 1805 1410 1895 1420
rect 2075 1410 2165 1420
rect 2345 1410 2435 1420
rect 2615 1410 2705 1420
rect 2885 1410 2975 1420
rect -335 1400 980 1410
rect -335 1350 -190 1400
rect -140 1350 120 1400
rect 170 1350 430 1400
rect 480 1350 740 1400
rect 790 1350 980 1400
rect -335 1340 980 1350
rect 1085 1400 3215 1410
rect 1085 1350 1285 1400
rect 1335 1350 1555 1400
rect 1605 1350 1825 1400
rect 1875 1350 2095 1400
rect 2145 1350 2365 1400
rect 2415 1350 2635 1400
rect 2685 1350 2905 1400
rect 2955 1350 3215 1400
rect 1085 1340 3215 1350
rect -210 1330 -120 1340
rect 100 1330 190 1340
rect 410 1330 500 1340
rect 720 1330 810 1340
rect 1265 1330 1355 1340
rect 1535 1330 1625 1340
rect 1805 1330 1895 1340
rect 2075 1330 2165 1340
rect 2345 1330 2435 1340
rect 2615 1330 2705 1340
rect 2885 1330 2975 1340
rect -55 1250 35 1260
rect 255 1250 345 1260
rect 565 1250 655 1260
rect 875 1250 965 1260
rect 1130 1250 1220 1260
rect 1400 1250 1490 1260
rect 1670 1250 1760 1260
rect 1940 1250 2030 1260
rect 2210 1250 2300 1260
rect 2480 1250 2570 1260
rect 2750 1250 2840 1260
rect 3020 1250 3110 1260
rect -335 1240 980 1250
rect -335 1190 -35 1240
rect 15 1190 275 1240
rect 325 1190 585 1240
rect 635 1190 895 1240
rect 945 1190 980 1240
rect -335 1180 980 1190
rect 1085 1240 3220 1250
rect 1085 1190 1150 1240
rect 1200 1190 1420 1240
rect 1470 1190 1690 1240
rect 1740 1190 1960 1240
rect 2010 1190 2230 1240
rect 2280 1190 2500 1240
rect 2550 1190 2770 1240
rect 2820 1190 3040 1240
rect 3090 1190 3220 1240
rect 1085 1180 3220 1190
rect -55 1170 35 1180
rect 255 1170 345 1180
rect 565 1170 655 1180
rect 875 1170 965 1180
rect 1130 1170 1220 1180
rect 1400 1170 1490 1180
rect 1670 1170 1760 1180
rect 1940 1170 2030 1180
rect 2210 1170 2300 1180
rect 2480 1170 2570 1180
rect 2750 1170 2840 1180
rect 3020 1170 3110 1180
rect -210 1090 -120 1100
rect 100 1090 190 1100
rect 410 1090 500 1100
rect 720 1090 810 1100
rect 1265 1090 1355 1100
rect 1535 1090 1625 1100
rect 1805 1090 1895 1100
rect 2075 1090 2165 1100
rect 2345 1090 2435 1100
rect 2615 1090 2705 1100
rect 2885 1090 2975 1100
rect -335 1080 980 1090
rect -335 1030 -190 1080
rect -140 1030 120 1080
rect 170 1030 430 1080
rect 480 1030 740 1080
rect 790 1030 980 1080
rect -335 1020 980 1030
rect 1085 1080 3215 1090
rect 1085 1030 1285 1080
rect 1335 1030 1555 1080
rect 1605 1030 1825 1080
rect 1875 1030 2095 1080
rect 2145 1030 2365 1080
rect 2415 1030 2635 1080
rect 2685 1030 2905 1080
rect 2955 1030 3215 1080
rect 1085 1020 3215 1030
rect -210 1010 -120 1020
rect 100 1010 190 1020
rect 410 1010 500 1020
rect 720 1010 810 1020
rect 1265 1010 1355 1020
rect 1535 1010 1625 1020
rect 1805 1010 1895 1020
rect 2075 1010 2165 1020
rect 2345 1010 2435 1020
rect 2615 1010 2705 1020
rect 2885 1010 2975 1020
rect -55 930 35 940
rect 255 930 345 940
rect 565 930 655 940
rect 875 930 965 940
rect 1130 930 1220 940
rect 1400 930 1490 940
rect 1670 930 1760 940
rect 1940 930 2030 940
rect 2210 930 2300 940
rect 2480 930 2570 940
rect 2750 930 2840 940
rect 3020 930 3110 940
rect -335 920 980 930
rect -335 870 -35 920
rect 15 870 275 920
rect 325 870 585 920
rect 635 870 895 920
rect 945 870 980 920
rect -335 860 980 870
rect 1085 920 3220 930
rect 1085 870 1150 920
rect 1200 870 1420 920
rect 1470 870 1690 920
rect 1740 870 1960 920
rect 2010 870 2230 920
rect 2280 870 2500 920
rect 2550 870 2770 920
rect 2820 870 3040 920
rect 3090 870 3220 920
rect 1085 860 3220 870
rect -55 850 35 860
rect 255 850 345 860
rect 565 850 655 860
rect 875 850 965 860
rect 1130 850 1220 860
rect 1400 850 1490 860
rect 1670 850 1760 860
rect 1940 850 2030 860
rect 2210 850 2300 860
rect 2480 850 2570 860
rect 2750 850 2840 860
rect 3020 850 3110 860
rect -210 770 -120 780
rect 100 770 190 780
rect 410 770 500 780
rect 720 770 810 780
rect 1265 770 1355 780
rect 1535 770 1625 780
rect 1805 770 1895 780
rect 2075 770 2165 780
rect 2345 770 2435 780
rect 2615 770 2705 780
rect 2885 770 2975 780
rect -335 760 980 770
rect -335 710 -190 760
rect -140 710 120 760
rect 170 710 430 760
rect 480 710 740 760
rect 790 710 980 760
rect -335 700 980 710
rect 1085 760 3215 770
rect 1085 710 1285 760
rect 1335 710 1555 760
rect 1605 710 1825 760
rect 1875 710 2095 760
rect 2145 710 2365 760
rect 2415 710 2635 760
rect 2685 710 2905 760
rect 2955 710 3215 760
rect 1085 700 3215 710
rect -210 690 -120 700
rect 100 690 190 700
rect 410 690 500 700
rect 720 690 810 700
rect 1265 690 1355 700
rect 1535 690 1625 700
rect 1805 690 1895 700
rect 2075 690 2165 700
rect 2345 690 2435 700
rect 2615 690 2705 700
rect 2885 690 2975 700
rect -55 610 35 620
rect 255 610 345 620
rect 565 610 655 620
rect 875 610 965 620
rect 1130 610 1220 620
rect 1400 610 1490 620
rect 1670 610 1760 620
rect 1940 610 2030 620
rect 2210 610 2300 620
rect 2480 610 2570 620
rect 2750 610 2840 620
rect 3020 610 3110 620
rect -335 600 980 610
rect -335 550 -35 600
rect 15 550 275 600
rect 325 550 585 600
rect 635 550 895 600
rect 945 550 980 600
rect -335 540 980 550
rect 1085 600 3220 610
rect 1085 550 1150 600
rect 1200 550 1420 600
rect 1470 550 1690 600
rect 1740 550 1960 600
rect 2010 550 2230 600
rect 2280 550 2500 600
rect 2550 550 2770 600
rect 2820 550 3040 600
rect 3090 550 3220 600
rect 1085 540 3220 550
rect -55 530 35 540
rect 255 530 345 540
rect 565 530 655 540
rect 875 530 965 540
rect 1130 530 1220 540
rect 1400 530 1490 540
rect 1670 530 1760 540
rect 1940 530 2030 540
rect 2210 530 2300 540
rect 2480 530 2570 540
rect 2750 530 2840 540
rect 3020 530 3110 540
rect 4005 475 4095 485
rect 3850 465 4335 475
rect -210 450 -120 460
rect 100 450 190 460
rect 410 450 500 460
rect 720 450 810 460
rect 1265 450 1355 460
rect 1535 450 1625 460
rect 1805 450 1895 460
rect 2075 450 2165 460
rect 2345 450 2435 460
rect 2615 450 2705 460
rect 2885 450 2975 460
rect -335 440 980 450
rect -335 390 -190 440
rect -140 390 120 440
rect 170 390 430 440
rect 480 390 740 440
rect 790 390 980 440
rect -335 380 980 390
rect 1085 440 3215 450
rect 1085 390 1285 440
rect 1335 390 1555 440
rect 1605 390 1825 440
rect 1875 390 2095 440
rect 2145 390 2365 440
rect 2415 390 2635 440
rect 2685 390 2905 440
rect 2955 390 3215 440
rect 3850 415 4025 465
rect 4075 415 4335 465
rect 3850 405 4335 415
rect 4005 395 4095 405
rect 1085 380 3215 390
rect -210 370 -120 380
rect 100 370 190 380
rect 410 370 500 380
rect 720 370 810 380
rect 1265 370 1355 380
rect 1535 370 1625 380
rect 1805 370 1895 380
rect 2075 370 2165 380
rect 2345 370 2435 380
rect 2615 370 2705 380
rect 2885 370 2975 380
rect 4005 315 4095 325
rect 3850 305 4340 315
rect -55 290 35 300
rect 255 290 345 300
rect 565 290 655 300
rect 875 290 965 300
rect 1130 290 1220 300
rect 1400 290 1490 300
rect 1670 290 1760 300
rect 1940 290 2030 300
rect 2210 290 2300 300
rect 2480 290 2570 300
rect 2750 290 2840 300
rect 3020 290 3110 300
rect -335 280 980 290
rect -335 230 -35 280
rect 15 230 275 280
rect 325 230 585 280
rect 635 230 895 280
rect 945 230 980 280
rect -335 220 980 230
rect 1085 280 3220 290
rect 1085 230 1150 280
rect 1200 230 1420 280
rect 1470 230 1690 280
rect 1740 230 1960 280
rect 2010 230 2230 280
rect 2280 230 2500 280
rect 2550 230 2770 280
rect 2820 230 3040 280
rect 3090 230 3220 280
rect 3850 255 4025 305
rect 4075 255 4340 305
rect 3850 245 4340 255
rect 4005 235 4095 245
rect 1085 220 3220 230
rect -55 210 35 220
rect 255 210 345 220
rect 565 210 655 220
rect 875 210 965 220
rect 1130 210 1220 220
rect 1400 210 1490 220
rect 1670 210 1760 220
rect 1940 210 2030 220
rect 2210 210 2300 220
rect 2480 210 2570 220
rect 2750 210 2840 220
rect 3020 210 3110 220
rect -210 130 -120 140
rect 100 130 190 140
rect 410 130 500 140
rect 720 130 810 140
rect 1265 130 1355 140
rect 1535 130 1625 140
rect 1805 130 1895 140
rect 2075 130 2165 140
rect 2345 130 2435 140
rect 2615 130 2705 140
rect 2885 130 2975 140
rect -335 120 980 130
rect -335 70 -190 120
rect -140 70 120 120
rect 170 70 430 120
rect 480 70 740 120
rect 790 70 980 120
rect -335 60 980 70
rect 1085 120 3215 130
rect 1085 70 1285 120
rect 1335 70 1555 120
rect 1605 70 1825 120
rect 1875 70 2095 120
rect 2145 70 2365 120
rect 2415 70 2635 120
rect 2685 70 2905 120
rect 2955 70 3215 120
rect 1085 60 3215 70
rect -210 50 -120 60
rect 100 50 190 60
rect 410 50 500 60
rect 720 50 810 60
rect 1265 50 1355 60
rect 1535 50 1625 60
rect 1805 50 1895 60
rect 2075 50 2165 60
rect 2345 50 2435 60
rect 2615 50 2705 60
rect 2885 50 2975 60
rect -55 -30 35 -20
rect 255 -30 345 -20
rect 565 -30 655 -20
rect 875 -30 965 -20
rect 1130 -30 1220 -20
rect 1400 -30 1490 -20
rect 1670 -30 1760 -20
rect 1940 -30 2030 -20
rect 2210 -30 2300 -20
rect 2480 -30 2570 -20
rect 2750 -30 2840 -20
rect 3020 -30 3110 -20
rect -335 -40 980 -30
rect -335 -90 -35 -40
rect 15 -90 275 -40
rect 325 -90 585 -40
rect 635 -90 895 -40
rect 945 -90 980 -40
rect -335 -100 980 -90
rect 1085 -40 3220 -30
rect 1085 -90 1150 -40
rect 1200 -90 1420 -40
rect 1470 -90 1690 -40
rect 1740 -90 1960 -40
rect 2010 -90 2230 -40
rect 2280 -90 2500 -40
rect 2550 -90 2770 -40
rect 2820 -90 3040 -40
rect 3090 -90 3220 -40
rect 1085 -100 3220 -90
rect -55 -110 35 -100
rect 255 -110 345 -100
rect 565 -110 655 -100
rect 875 -110 965 -100
rect 1130 -110 1220 -100
rect 1400 -110 1490 -100
rect 1670 -110 1760 -100
rect 1940 -110 2030 -100
rect 2210 -110 2300 -100
rect 2480 -110 2570 -100
rect 2750 -110 2840 -100
rect 3020 -110 3110 -100
<< via2 >>
rect -190 1350 -140 1400
rect 120 1350 170 1400
rect 430 1350 480 1400
rect 740 1350 790 1400
rect -35 1190 15 1240
rect 275 1190 325 1240
rect 585 1190 635 1240
rect 895 1190 945 1240
rect -190 1030 -140 1080
rect 120 1030 170 1080
rect 430 1030 480 1080
rect 740 1030 790 1080
rect -35 870 15 920
rect 275 870 325 920
rect 585 870 635 920
rect 895 870 945 920
rect -190 710 -140 760
rect 120 710 170 760
rect 430 710 480 760
rect 740 710 790 760
rect -35 550 15 600
rect 275 550 325 600
rect 585 550 635 600
rect 895 550 945 600
rect -190 390 -140 440
rect 120 390 170 440
rect 430 390 480 440
rect 740 390 790 440
rect -35 230 15 280
rect 275 230 325 280
rect 585 230 635 280
rect 895 230 945 280
rect -190 70 -140 120
rect 120 70 170 120
rect 430 70 480 120
rect 740 70 790 120
rect -35 -90 15 -40
rect 275 -90 325 -40
rect 585 -90 635 -40
rect 895 -90 945 -40
<< metal3 >>
rect -205 1420 -125 1595
rect -210 1400 -120 1420
rect -210 1350 -190 1400
rect -140 1350 -120 1400
rect -210 1330 -120 1350
rect -205 1100 -125 1330
rect -50 1260 30 1595
rect 105 1420 185 1595
rect 100 1400 190 1420
rect 100 1350 120 1400
rect 170 1350 190 1400
rect 100 1330 190 1350
rect -55 1240 35 1260
rect -55 1190 -35 1240
rect 15 1190 35 1240
rect -55 1170 35 1190
rect -210 1080 -120 1100
rect -210 1030 -190 1080
rect -140 1030 -120 1080
rect -210 1010 -120 1030
rect -205 780 -125 1010
rect -50 940 30 1170
rect 105 1100 185 1330
rect 260 1260 340 1595
rect 415 1420 495 1595
rect 410 1400 500 1420
rect 410 1350 430 1400
rect 480 1350 500 1400
rect 410 1330 500 1350
rect 255 1240 345 1260
rect 255 1190 275 1240
rect 325 1190 345 1240
rect 255 1170 345 1190
rect 100 1080 190 1100
rect 100 1030 120 1080
rect 170 1030 190 1080
rect 100 1010 190 1030
rect -55 920 35 940
rect -55 870 -35 920
rect 15 870 35 920
rect -55 850 35 870
rect -210 760 -120 780
rect -210 710 -190 760
rect -140 710 -120 760
rect -210 690 -120 710
rect -205 460 -125 690
rect -50 620 30 850
rect 105 780 185 1010
rect 260 940 340 1170
rect 415 1100 495 1330
rect 570 1260 650 1595
rect 725 1420 805 1595
rect 720 1400 810 1420
rect 720 1350 740 1400
rect 790 1350 810 1400
rect 720 1330 810 1350
rect 565 1240 655 1260
rect 565 1190 585 1240
rect 635 1190 655 1240
rect 565 1170 655 1190
rect 410 1080 500 1100
rect 410 1030 430 1080
rect 480 1030 500 1080
rect 410 1010 500 1030
rect 255 920 345 940
rect 255 870 275 920
rect 325 870 345 920
rect 255 850 345 870
rect 100 760 190 780
rect 100 710 120 760
rect 170 710 190 760
rect 100 690 190 710
rect -55 600 35 620
rect -55 550 -35 600
rect 15 550 35 600
rect -55 530 35 550
rect -210 440 -120 460
rect -210 390 -190 440
rect -140 390 -120 440
rect -210 370 -120 390
rect -205 140 -125 370
rect -50 300 30 530
rect 105 460 185 690
rect 260 620 340 850
rect 415 780 495 1010
rect 570 940 650 1170
rect 725 1100 805 1330
rect 880 1260 960 1595
rect 875 1240 965 1260
rect 875 1190 895 1240
rect 945 1190 965 1240
rect 875 1170 965 1190
rect 720 1080 810 1100
rect 720 1030 740 1080
rect 790 1030 810 1080
rect 720 1010 810 1030
rect 565 920 655 940
rect 565 870 585 920
rect 635 870 655 920
rect 565 850 655 870
rect 410 760 500 780
rect 410 710 430 760
rect 480 710 500 760
rect 410 690 500 710
rect 255 600 345 620
rect 255 550 275 600
rect 325 550 345 600
rect 255 530 345 550
rect 100 440 190 460
rect 100 390 120 440
rect 170 390 190 440
rect 100 370 190 390
rect -55 280 35 300
rect -55 230 -35 280
rect 15 230 35 280
rect -55 210 35 230
rect -210 120 -120 140
rect -210 70 -190 120
rect -140 70 -120 120
rect -210 50 -120 70
rect -205 -150 -125 50
rect -50 -20 30 210
rect 105 140 185 370
rect 260 300 340 530
rect 415 460 495 690
rect 570 620 650 850
rect 725 780 805 1010
rect 880 940 960 1170
rect 875 920 965 940
rect 875 870 895 920
rect 945 870 965 920
rect 875 850 965 870
rect 720 760 810 780
rect 720 710 740 760
rect 790 710 810 760
rect 720 690 810 710
rect 565 600 655 620
rect 565 550 585 600
rect 635 550 655 600
rect 565 530 655 550
rect 410 440 500 460
rect 410 390 430 440
rect 480 390 500 440
rect 410 370 500 390
rect 255 280 345 300
rect 255 230 275 280
rect 325 230 345 280
rect 255 210 345 230
rect 100 120 190 140
rect 100 70 120 120
rect 170 70 190 120
rect 100 50 190 70
rect -55 -40 35 -20
rect -55 -90 -35 -40
rect 15 -90 35 -40
rect -55 -110 35 -90
rect -50 -150 30 -110
rect 105 -150 185 50
rect 260 -20 340 210
rect 415 140 495 370
rect 570 300 650 530
rect 725 460 805 690
rect 880 620 960 850
rect 875 600 965 620
rect 875 550 895 600
rect 945 550 965 600
rect 875 530 965 550
rect 720 440 810 460
rect 720 390 740 440
rect 790 390 810 440
rect 720 370 810 390
rect 565 280 655 300
rect 565 230 585 280
rect 635 230 655 280
rect 565 210 655 230
rect 410 120 500 140
rect 410 70 430 120
rect 480 70 500 120
rect 410 50 500 70
rect 255 -40 345 -20
rect 255 -90 275 -40
rect 325 -90 345 -40
rect 255 -110 345 -90
rect 260 -150 340 -110
rect 415 -150 495 50
rect 570 -20 650 210
rect 725 140 805 370
rect 880 300 960 530
rect 875 280 965 300
rect 875 230 895 280
rect 945 230 965 280
rect 875 210 965 230
rect 720 120 810 140
rect 720 70 740 120
rect 790 70 810 120
rect 720 50 810 70
rect 565 -40 655 -20
rect 565 -90 585 -40
rect 635 -90 655 -40
rect 565 -110 655 -90
rect 570 -150 650 -110
rect 725 -150 805 50
rect 880 -20 960 210
rect 875 -40 965 -20
rect 875 -90 895 -40
rect 945 -90 965 -40
rect 875 -110 965 -90
rect 880 -150 960 -110
<< end >>
