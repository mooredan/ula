* Functional simulation of pad_x0_top and pad_in_top

* .include mag/pad_xtal.cir
.include mag/pad_x0_top.cir
.include mag/pad_in_top.cir

.lib device_models/AMI_C5N.lib TT
.lib device_models/AMI_C5N_rmodels.lib NOM 

.param VDD_VAL=5
+      FREQ=6.5Meg
+      PER={1 / FREQ}
+      PH={PER / 2.0}
+      TRF={PER * 0.1}


* power supply
Vvdd vdd 0 DC VDD_VAL
Vvss vss 0 DC 0

* input signal
* with 50 ohm output impedance
* SIN(VO VA FREQ) VO=offset VA=amplitude
* Voffset indc 0 DC {VDD_VAL/2.0}

* Vin x1 0 SIN({VDD_VAL/2.0} 0.5 {FREQ})
Voffset offset 0 DC {VDD_VAL/2.0}
Vin x1 offset DC 0 AC {VDD_VAL/10.0} 
* Vin x1 0 DC 0

* Vdout dout indc  DC 0
* + PULSE({VDD_VAL/-2.0} {VDD_VAL/2.0} {PER/2.0} {TRF} {TRF} {PH-TRF} {PER}) 

* Voe oe 0 DC {VDD_VAL} PWL(0 {VDD_VAL} 400n {VDD_VAL} 401n 0 3u 0 3.005u {VDD_VAL})

* .subckt pad_xtal x0 x1 vdd vss
Xdut x0 x1 vdd vss pad_xtal
Rf x0 x1 5Meg

* output load
* Cx0 x0 0 1p
Rl x0 rn 10k
Vl rn 0 DC 0

* .save all @r.xdut.rin1[i] @Cout[i]
* .save all @m.xdut.xpad_io_top_0.m1002[id]
* +         @m.xdut.xpad_io_top_0.m1010[id]
.save all

.op

* .tran 0.1n {PER*5}
* .dc Vin 0 {VDD_VAL} 0.01
.ac lin 100 0.100Meg 10.000Meg



.control
destroy all
run

* setplot dc1 
* plot v(a) v(pad)
* plot i(vvdd)

* setplot tran1
* plot v(x1) v(x0)
* let freq = 6.5e6
* let per = 1.0 / freq

setplot ac1
plot vdb(x1) vdb(x0)

let zin = v(x1) / -i(Vin)
let zout = v(x0) / i(Vl)

* plot re(zin)

* meas tran x0_avg avg v(x0) from={PER} to={2.0*PER}
* meas tran x1_avg avg v(x1) from={PER} to={2.0*PER}
* meas tran x0_rms rms v(x0) from={PER} to={2.0*PER}
* meas tran x1_rms rms v(x1) from={PER} to={2.0*PER}

* let x0_amp = x0_rms - x0_avg
* let x1_amp = x1_rms - x1_avg

* let AV = x0_amp / x1_amp
* print x0_amp
* print x1_amp
* print AV


* setplot dc1
* plot v(x1) v(x0)
* plot @m.xdut.xpad_io_top_0.m1002[id] @m.xdut.xpad_io_top_0.m1010[id]

* setplot ac1
* plot vdb(pad)

let idx = 64 
* 
while idx <=  64 
*   let zin = v(in) / l.xdut.xpk14.l1#branch
   print idx
   print zin[idx]
   print abs(zin[idx])
   print abs(frequency[idx])
   print real(zin[idx])
   print imag(zin[idx])
   let Xin = imag(zin[idx])
   print mag(zin[idx])
   print ph(zin[idx]) * 180 / pi
   let omega = 2 * pi * abs(frequency[idx])
   let Xcin = -Xin
   let Cin = 1 / (omega * Xcin)
   print Cin
* 
* *  let zout = v(pad) / l.xdut.lout2#branch
  print zout[idx]
  print abs(zout[idx])
  print real(zout[idx])
  print imag(zout[idx])
  let Xout = imag(zout[idx])
  print mag(zout[idx])
  print ph(zout[idx]) * 180 / pi
  if ( Xout < 0 ) 
     let Xcout = -Xout
     let Cout = 1 / (omega * Xcout)
     print Cout
  else 
     let Xlout = Xout
     let Lout = (omega * Xlout)
     print Lout
  end
*   
*  
  let idx = idx + 1
end
.endc

.end
