`celldefine
module inv_c (z, a);
  output z;
  input  a;

  not G1 (z, a);
endmodule
`endcelldefine
