* Output transition times
* .include mag/dly_test.cir
* .include mag/dly_c.cir
.include mag/nand2_b.cir
.include mag/nand2_c.cir
.include mag/nor2_c.cir
.include mag/nor2_b.cir
.include mag/subc_2.cir
.include mag/schmitt.cir
.include mag/inv_d.cir
.include mag/inv_e.cir
.include mag/pad_io_bot.cir

.lib device_models/AMI_C5N.lib TT
.lib device_models/AMI_C5N_rmodels.lib NOM 

.temp 25

.param VDD_VAL=5

* power supply
vvdd vdd 0 DC VDD_VAL
vvss vss 0 DC 0


*************************************
* .subckt pad_io_bot tri ntri xpad din pd npu vdd vss

Xdut tri ntri xpad din pd npu vdd vss pad_io_bot

*************************************
* vnpd  npd 0 DC 0 PULSE(0 {VDD_VAL} 10n 4.8n 4.8n 80n 220n)
va  xdut.a 0 DC 0 PULSE(0 {VDD_VAL} 10n 4.8n 4.8n 80n 220n)
vadly  xdut.adly 0 DC 0 PULSE(0 {VDD_VAL} 10n 4.8n 4.8n 80n 220n)
* vdin    din 0 DC 0 PULSE(0 {VDD_VAL} 10n 4.8n 4.8n 45.2n 100n)
Vxpad xpad 0 DC 0
Vntri ntri 0 DC 5
Vtri tri 0 DC 0


* output load
* cpad pad vgnd 50p
* vvgnd vgnd 0 DC 0

* add small load to core side of the
* input series resistor


.save all

.op
* .tran 0.1n 900n

.control
destroy all
run

* setplot tran1
* plot v(a) v(zout)
* plot  v(node1)  v(node2)

print v(vdd)

* let vdd_max = maximum(v(vdd))
* let vol = vdd_max * 0.1
* let voh = vdd_max * 0.9
* 
* print vdd_max
* print vol
* print voh
* 
* 
* meas tran nputlh TRIG v(xdut.npu) VAL=vol RISE=1 TARG v(xdut.npu) VAL=voh RISE=1
* meas tran nputhl TRIG v(xdut.npu) VAL=voh FALL=2 TARG v(xdut.npu) VAL=vol FALL=2
* meas tran padtlh TRIG v(pad) VAL=vol RISE=2 TARG v(pad) VAL=voh RISE=2
* 
* meas tran pdtlh TRIG v(xdut.pd) VAL=vol RISE=1 TARG v(xdut.pd) VAL=voh RISE=1
* meas tran pdthl TRIG v(xdut.pd) VAL=voh FALL=2 TARG v(xdut.pd) VAL=vol FALL=2
* meas tran padthl TRIG v(pad) VAL=voh FALL=1 TARG v(pad) VAL=vol FALL=1

.endc

.end
