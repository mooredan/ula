magic
tech amic5n
timestamp 1622329769
<< nwell >>
rect 895 805 2065 2455
<< ntransistor >>
rect 1165 95 1225 655
rect 1355 95 1415 655
rect 1545 95 1605 655
rect 1735 95 1795 655
<< ptransistor >>
rect 1165 955 1225 2305
rect 1355 955 1415 2305
rect 1545 955 1605 2305
rect 1735 955 1795 2305
<< nselect >>
rect 1000 0 1960 685
<< pselect >>
rect 1000 925 1960 2400
<< ndiffusion >>
rect 1045 625 1165 655
rect 1045 575 1075 625
rect 1125 575 1165 625
rect 1045 475 1165 575
rect 1045 425 1075 475
rect 1125 425 1165 475
rect 1045 375 1165 425
rect 1045 325 1075 375
rect 1125 325 1165 375
rect 1045 275 1165 325
rect 1045 225 1075 275
rect 1125 225 1165 275
rect 1045 175 1165 225
rect 1045 125 1075 175
rect 1125 125 1165 175
rect 1045 95 1165 125
rect 1225 625 1355 655
rect 1225 575 1265 625
rect 1315 575 1355 625
rect 1225 475 1355 575
rect 1225 425 1265 475
rect 1315 425 1355 475
rect 1225 375 1355 425
rect 1225 325 1265 375
rect 1315 325 1355 375
rect 1225 275 1355 325
rect 1225 225 1265 275
rect 1315 225 1355 275
rect 1225 175 1355 225
rect 1225 125 1265 175
rect 1315 125 1355 175
rect 1225 95 1355 125
rect 1415 625 1545 655
rect 1415 575 1455 625
rect 1505 575 1545 625
rect 1415 475 1545 575
rect 1415 425 1455 475
rect 1505 425 1545 475
rect 1415 375 1545 425
rect 1415 325 1455 375
rect 1505 325 1545 375
rect 1415 275 1545 325
rect 1415 225 1455 275
rect 1505 225 1545 275
rect 1415 175 1545 225
rect 1415 125 1455 175
rect 1505 125 1545 175
rect 1415 95 1545 125
rect 1605 625 1735 655
rect 1605 575 1645 625
rect 1695 575 1735 625
rect 1605 475 1735 575
rect 1605 425 1645 475
rect 1695 425 1735 475
rect 1605 375 1735 425
rect 1605 325 1645 375
rect 1695 325 1735 375
rect 1605 275 1735 325
rect 1605 225 1645 275
rect 1695 225 1735 275
rect 1605 175 1735 225
rect 1605 125 1645 175
rect 1695 125 1735 175
rect 1605 95 1735 125
rect 1795 625 1915 655
rect 1795 575 1835 625
rect 1885 575 1915 625
rect 1795 475 1915 575
rect 1795 425 1835 475
rect 1885 425 1915 475
rect 1795 375 1915 425
rect 1795 325 1835 375
rect 1885 325 1915 375
rect 1795 275 1915 325
rect 1795 225 1835 275
rect 1885 225 1915 275
rect 1795 175 1915 225
rect 1795 125 1835 175
rect 1885 125 1915 175
rect 1795 95 1915 125
<< pdiffusion >>
rect 1045 2275 1165 2305
rect 1045 2225 1075 2275
rect 1125 2225 1165 2275
rect 1045 2135 1165 2225
rect 1045 2085 1075 2135
rect 1125 2085 1165 2135
rect 1045 2035 1165 2085
rect 1045 1985 1075 2035
rect 1125 1985 1165 2035
rect 1045 1935 1165 1985
rect 1045 1885 1075 1935
rect 1125 1885 1165 1935
rect 1045 1835 1165 1885
rect 1045 1785 1075 1835
rect 1125 1785 1165 1835
rect 1045 1735 1165 1785
rect 1045 1685 1075 1735
rect 1125 1685 1165 1735
rect 1045 1635 1165 1685
rect 1045 1585 1075 1635
rect 1125 1585 1165 1635
rect 1045 1535 1165 1585
rect 1045 1485 1075 1535
rect 1125 1485 1165 1535
rect 1045 1435 1165 1485
rect 1045 1385 1075 1435
rect 1125 1385 1165 1435
rect 1045 1335 1165 1385
rect 1045 1285 1075 1335
rect 1125 1285 1165 1335
rect 1045 1235 1165 1285
rect 1045 1185 1075 1235
rect 1125 1185 1165 1235
rect 1045 1135 1165 1185
rect 1045 1085 1075 1135
rect 1125 1085 1165 1135
rect 1045 955 1165 1085
rect 1225 955 1355 2305
rect 1415 2235 1545 2305
rect 1415 2185 1455 2235
rect 1505 2185 1545 2235
rect 1415 2135 1545 2185
rect 1415 2085 1455 2135
rect 1505 2085 1545 2135
rect 1415 2035 1545 2085
rect 1415 1985 1455 2035
rect 1505 1985 1545 2035
rect 1415 1935 1545 1985
rect 1415 1885 1455 1935
rect 1505 1885 1545 1935
rect 1415 1835 1545 1885
rect 1415 1785 1455 1835
rect 1505 1785 1545 1835
rect 1415 1735 1545 1785
rect 1415 1685 1455 1735
rect 1505 1685 1545 1735
rect 1415 1635 1545 1685
rect 1415 1585 1455 1635
rect 1505 1585 1545 1635
rect 1415 1535 1545 1585
rect 1415 1485 1455 1535
rect 1505 1485 1545 1535
rect 1415 1435 1545 1485
rect 1415 1385 1455 1435
rect 1505 1385 1545 1435
rect 1415 1245 1545 1385
rect 1415 1195 1455 1245
rect 1505 1195 1545 1245
rect 1415 1145 1545 1195
rect 1415 1095 1455 1145
rect 1505 1095 1545 1145
rect 1415 955 1545 1095
rect 1605 955 1735 2305
rect 1795 2275 1915 2305
rect 1795 2225 1835 2275
rect 1885 2225 1915 2275
rect 1795 2135 1915 2225
rect 1795 2085 1835 2135
rect 1885 2085 1915 2135
rect 1795 2035 1915 2085
rect 1795 1985 1835 2035
rect 1885 1985 1915 2035
rect 1795 1935 1915 1985
rect 1795 1885 1835 1935
rect 1885 1885 1915 1935
rect 1795 1835 1915 1885
rect 1795 1785 1835 1835
rect 1885 1785 1915 1835
rect 1795 1735 1915 1785
rect 1795 1685 1835 1735
rect 1885 1685 1915 1735
rect 1795 1635 1915 1685
rect 1795 1585 1835 1635
rect 1885 1585 1915 1635
rect 1795 1535 1915 1585
rect 1795 1485 1835 1535
rect 1885 1485 1915 1535
rect 1795 1435 1915 1485
rect 1795 1385 1835 1435
rect 1885 1385 1915 1435
rect 1795 1335 1915 1385
rect 1795 1285 1835 1335
rect 1885 1285 1915 1335
rect 1795 1235 1915 1285
rect 1795 1185 1835 1235
rect 1885 1185 1915 1235
rect 1795 1135 1915 1185
rect 1795 1085 1835 1135
rect 1885 1085 1915 1135
rect 1795 1035 1915 1085
rect 1795 985 1835 1035
rect 1885 985 1915 1035
rect 1795 955 1915 985
<< ndcontact >>
rect 1075 575 1125 625
rect 1075 425 1125 475
rect 1075 325 1125 375
rect 1075 225 1125 275
rect 1075 125 1125 175
rect 1265 575 1315 625
rect 1265 425 1315 475
rect 1265 325 1315 375
rect 1265 225 1315 275
rect 1265 125 1315 175
rect 1455 575 1505 625
rect 1455 425 1505 475
rect 1455 325 1505 375
rect 1455 225 1505 275
rect 1455 125 1505 175
rect 1645 575 1695 625
rect 1645 425 1695 475
rect 1645 325 1695 375
rect 1645 225 1695 275
rect 1645 125 1695 175
rect 1835 575 1885 625
rect 1835 425 1885 475
rect 1835 325 1885 375
rect 1835 225 1885 275
rect 1835 125 1885 175
<< pdcontact >>
rect 1075 2225 1125 2275
rect 1075 2085 1125 2135
rect 1075 1985 1125 2035
rect 1075 1885 1125 1935
rect 1075 1785 1125 1835
rect 1075 1685 1125 1735
rect 1075 1585 1125 1635
rect 1075 1485 1125 1535
rect 1075 1385 1125 1435
rect 1075 1285 1125 1335
rect 1075 1185 1125 1235
rect 1075 1085 1125 1135
rect 1455 2185 1505 2235
rect 1455 2085 1505 2135
rect 1455 1985 1505 2035
rect 1455 1885 1505 1935
rect 1455 1785 1505 1835
rect 1455 1685 1505 1735
rect 1455 1585 1505 1635
rect 1455 1485 1505 1535
rect 1455 1385 1505 1435
rect 1455 1195 1505 1245
rect 1455 1095 1505 1145
rect 1835 2225 1885 2275
rect 1835 2085 1885 2135
rect 1835 1985 1885 2035
rect 1835 1885 1885 1935
rect 1835 1785 1885 1835
rect 1835 1685 1885 1735
rect 1835 1585 1885 1635
rect 1835 1485 1885 1535
rect 1835 1385 1885 1435
rect 1835 1285 1885 1335
rect 1835 1185 1885 1235
rect 1835 1085 1885 1135
rect 1835 985 1885 1035
<< polysilicon >>
rect 1165 2305 1225 2370
rect 1355 2305 1415 2370
rect 1545 2305 1605 2370
rect 1735 2305 1795 2370
rect 1165 845 1225 955
rect 1055 825 1225 845
rect 1055 775 1075 825
rect 1125 775 1225 825
rect 1055 755 1225 775
rect 1165 655 1225 755
rect 1355 930 1415 955
rect 1545 930 1605 955
rect 1355 825 1605 930
rect 1355 775 1455 825
rect 1505 775 1605 825
rect 1355 695 1605 775
rect 1355 655 1415 695
rect 1545 655 1605 695
rect 1735 845 1795 955
rect 1735 825 1905 845
rect 1735 775 1835 825
rect 1885 775 1905 825
rect 1735 755 1905 775
rect 1735 655 1795 755
rect 1165 30 1225 95
rect 1355 30 1415 95
rect 1545 30 1605 95
rect 1735 30 1795 95
<< polycontact >>
rect 1075 775 1125 825
rect 1455 775 1505 825
rect 1835 775 1885 825
<< metal1 >>
rect 1000 2355 1960 2445
rect 1055 2275 1145 2355
rect 1055 2225 1075 2275
rect 1125 2225 1145 2275
rect 1815 2275 1905 2355
rect 1055 2135 1145 2225
rect 1055 2085 1075 2135
rect 1125 2085 1145 2135
rect 1055 2035 1145 2085
rect 1055 1985 1075 2035
rect 1125 1985 1145 2035
rect 1055 1935 1145 1985
rect 1055 1885 1075 1935
rect 1125 1885 1145 1935
rect 1055 1835 1145 1885
rect 1055 1785 1075 1835
rect 1125 1785 1145 1835
rect 1055 1735 1145 1785
rect 1055 1685 1075 1735
rect 1125 1685 1145 1735
rect 1055 1635 1145 1685
rect 1055 1585 1075 1635
rect 1125 1585 1145 1635
rect 1055 1535 1145 1585
rect 1055 1485 1075 1535
rect 1125 1485 1145 1535
rect 1055 1435 1145 1485
rect 1055 1385 1075 1435
rect 1125 1385 1145 1435
rect 1055 1335 1145 1385
rect 1055 1285 1075 1335
rect 1125 1285 1145 1335
rect 1055 1235 1145 1285
rect 1435 2235 1525 2255
rect 1435 2185 1455 2235
rect 1505 2185 1525 2235
rect 1435 2135 1525 2185
rect 1435 2085 1455 2135
rect 1505 2085 1525 2135
rect 1435 2035 1525 2085
rect 1435 1985 1455 2035
rect 1505 1985 1525 2035
rect 1435 1935 1525 1985
rect 1435 1885 1455 1935
rect 1505 1885 1525 1935
rect 1435 1835 1525 1885
rect 1435 1785 1455 1835
rect 1505 1785 1525 1835
rect 1435 1735 1525 1785
rect 1435 1685 1455 1735
rect 1505 1685 1525 1735
rect 1435 1635 1525 1685
rect 1435 1585 1455 1635
rect 1505 1585 1525 1635
rect 1435 1535 1525 1585
rect 1435 1485 1455 1535
rect 1505 1485 1525 1535
rect 1435 1435 1525 1485
rect 1435 1385 1455 1435
rect 1505 1385 1525 1435
rect 1435 1275 1525 1385
rect 1815 2225 1835 2275
rect 1885 2225 1905 2275
rect 1815 2135 1905 2225
rect 1815 2085 1835 2135
rect 1885 2085 1905 2135
rect 1815 2035 1905 2085
rect 1815 1985 1835 2035
rect 1885 1985 1905 2035
rect 1815 1935 1905 1985
rect 1815 1885 1835 1935
rect 1885 1885 1905 1935
rect 1815 1835 1905 1885
rect 1815 1785 1835 1835
rect 1885 1785 1905 1835
rect 1815 1735 1905 1785
rect 1815 1685 1835 1735
rect 1885 1685 1905 1735
rect 1815 1635 1905 1685
rect 1815 1585 1835 1635
rect 1885 1585 1905 1635
rect 1815 1535 1905 1585
rect 1815 1485 1835 1535
rect 1885 1485 1905 1535
rect 1815 1435 1905 1485
rect 1815 1385 1835 1435
rect 1885 1385 1905 1435
rect 1815 1335 1905 1385
rect 1815 1285 1835 1335
rect 1885 1285 1905 1335
rect 1055 1185 1075 1235
rect 1125 1185 1145 1235
rect 1055 1135 1145 1185
rect 1055 1085 1075 1135
rect 1125 1085 1145 1135
rect 1055 975 1145 1085
rect 1245 1245 1715 1275
rect 1245 1195 1455 1245
rect 1505 1195 1715 1245
rect 1245 1145 1715 1195
rect 1245 1095 1455 1145
rect 1505 1095 1715 1145
rect 1245 1075 1715 1095
rect 1055 825 1145 915
rect 1055 775 1075 825
rect 1125 775 1145 825
rect 1055 705 1145 775
rect 1055 625 1145 645
rect 1055 575 1075 625
rect 1125 575 1145 625
rect 1055 475 1145 575
rect 1055 425 1075 475
rect 1125 425 1145 475
rect 1055 375 1145 425
rect 1055 325 1075 375
rect 1125 325 1145 375
rect 1055 275 1145 325
rect 1055 225 1075 275
rect 1125 225 1145 275
rect 1055 175 1145 225
rect 1055 125 1075 175
rect 1125 125 1145 175
rect 1055 45 1145 125
rect 1245 625 1335 1075
rect 1435 825 1525 1005
rect 1435 775 1455 825
rect 1505 775 1525 825
rect 1435 755 1525 775
rect 1245 575 1265 625
rect 1315 575 1335 625
rect 1245 475 1335 575
rect 1245 425 1265 475
rect 1315 425 1335 475
rect 1245 375 1335 425
rect 1245 325 1265 375
rect 1315 325 1335 375
rect 1245 275 1335 325
rect 1245 225 1265 275
rect 1315 225 1335 275
rect 1245 175 1335 225
rect 1245 125 1265 175
rect 1315 125 1335 175
rect 1245 105 1335 125
rect 1435 625 1525 645
rect 1435 575 1455 625
rect 1505 575 1525 625
rect 1435 475 1525 575
rect 1435 425 1455 475
rect 1505 425 1525 475
rect 1435 375 1525 425
rect 1435 325 1455 375
rect 1505 325 1525 375
rect 1435 275 1525 325
rect 1435 225 1455 275
rect 1505 225 1525 275
rect 1435 175 1525 225
rect 1435 125 1455 175
rect 1505 125 1525 175
rect 1435 45 1525 125
rect 1625 625 1715 1075
rect 1815 1235 1905 1285
rect 1815 1185 1835 1235
rect 1885 1185 1905 1235
rect 1815 1135 1905 1185
rect 1815 1085 1835 1135
rect 1885 1085 1905 1135
rect 1815 1035 1905 1085
rect 1815 985 1835 1035
rect 1885 985 1905 1035
rect 1815 965 1905 985
rect 1815 825 1905 845
rect 1815 775 1835 825
rect 1885 775 1905 825
rect 1815 755 1905 775
rect 1625 575 1645 625
rect 1695 575 1715 625
rect 1625 475 1715 575
rect 1625 425 1645 475
rect 1695 425 1715 475
rect 1625 375 1715 425
rect 1625 325 1645 375
rect 1695 325 1715 375
rect 1625 275 1715 325
rect 1625 225 1645 275
rect 1695 225 1715 275
rect 1625 175 1715 225
rect 1625 125 1645 175
rect 1695 125 1715 175
rect 1625 105 1715 125
rect 1815 625 1905 645
rect 1815 575 1835 625
rect 1885 575 1905 625
rect 1815 475 1905 575
rect 1815 425 1835 475
rect 1885 425 1905 475
rect 1815 375 1905 425
rect 1815 325 1835 375
rect 1885 325 1905 375
rect 1815 275 1905 325
rect 1815 225 1835 275
rect 1885 225 1905 275
rect 1815 175 1905 225
rect 1815 125 1835 175
rect 1885 125 1905 175
rect 1815 45 1905 125
rect 1000 -45 1960 45
<< via1 >>
rect 1075 775 1125 825
rect 1835 775 1885 825
<< metal2 >>
rect 1055 825 1145 845
rect 1055 775 1075 825
rect 1125 775 1145 825
rect 1055 685 1145 775
rect 1815 825 1905 845
rect 1815 775 1835 825
rect 1885 775 1905 825
rect 1815 685 1905 775
rect 1055 595 1905 685
<< labels >>
flabel metal1 s 1075 765 1075 765 2 FreeSans 400 0 0 0 a
port 2 ne
flabel metal1 s 1065 2375 1065 2375 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 1075 -25 1075 -25 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 1275 725 1275 725 2 FreeSans 400 0 0 0 z
port 1 ne
flabel nwell 1020 915 1020 915 8 FreeSans 400 180 0 0 vdd
flabel ndiffusion s 1245 1510 1245 1510 2 FreeSans 400 0 0 0 x1
flabel ndiffusion s 1645 1495 1645 1495 2 FreeSans 400 0 0 0 x2
flabel metal1 s 1445 770 1445 770 2 FreeSans 400 0 0 0 b
port 3 ne
<< end >>
