magic
tech amic5n
timestamp 1608317707
<< poly2 >>
rect 73830 21270 74970 22410
<< poly2cap >>
rect 16740 13500 17880 14640
rect 37650 7800 38790 8940
rect 180 210 570 570
rect 17820 390 18960 1530
<< poly2capcontact >>
rect 16895 13655 16945 13705
<< poly2capcontact >>
rect 17975 545 18025 595
<< poly2capcontact >>
rect 335 365 385 415
<< polysilicon >>
rect 58140 20610 59640 22110
rect 16560 14640 18060 14790
rect 16560 13500 16740 14640
rect 17880 13500 18060 14640
rect 16560 13290 18060 13500
rect -2940 8400 -1440 9900
rect 37470 8940 38970 9090
rect 37470 7800 37650 8940
rect 38790 7800 38970 8940
rect 37470 7590 38970 7800
rect 17640 1530 19140 1680
rect 0 570 1500 1500
rect 0 210 180 570
rect 570 210 1500 570
rect 0 0 1500 210
rect 17640 390 17820 1530
rect 18960 390 19140 1530
rect 17640 180 19140 390
<< metal1 >>
rect 58440 20940 59370 21870
rect 73950 21390 74880 22320
rect 45690 19890 46620 20820
rect 16860 13620 17790 14550
rect 37770 7920 38700 8850
rect 17940 510 18060 630
rect 300 330 420 450
<< labels >>
flabel polysilicon s 30 30 30 30 2 FreeSans 400 0 0 0 a
flabel metal1 s 330 360 330 360 2 FreeSans 400 0 0 0 b
flabel polysilicon s -2790 8550 -2790 8550 2 FreeSans 400 0 0 0 c
flabel polysilicon s 17670 210 17670 210 2 FreeSans 400 0 0 0 a1
flabel metal1 s 17970 540 17970 540 2 FreeSans 400 0 0 0 b1
flabel polysilicon s 16590 13320 16590 13320 2 FreeSans 400 0 0 0 a2
flabel electrode s 16890 13650 16890 13650 2 FreeSans 400 0 0 0 b2
flabel polysilicon s 37500 7620 37500 7620 2 FreeSans 400 0 0 0 a3
flabel metal1 s 37800 7950 37800 7950 2 FreeSans 400 0 0 0 c3
flabel electrode s 37710 7860 37710 7860 2 FreeSans 400 0 0 0 b3
flabel metal1 s 45720 19920 45720 19920 2 FreeSans 400 0 0 0 n1
flabel polysilicon s 58170 20640 58170 20640 2 FreeSans 400 0 0 0 p2
flabel metal1 s 58470 20970 58470 20970 2 FreeSans 400 0 0 0 n2
flabel metal1 s 73980 21420 73980 21420 2 FreeSans 400 0 0 0 c4
flabel electrode s 73890 21330 73890 21330 2 FreeSans 400 0 0 0 b4
<< checkpaint >>
rect -2950 -10 74980 22420
<< end >>
