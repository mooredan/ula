magic
tech amic5n
timestamp 1607100556
<< metal1 >>
rect 0 0 46350 46350
<< end >>
