# LEF 

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.050 ;

USEMINSPACING OBS ON ;
CLEARANCEMEASURE EUCLIDEAN ;

# LAYER nwell
#   TYPE	MASTERSLICE ;
# END nwell
# 
# LAYER nactive
#   TYPE	MASTERSLICE ;
# END nactive
# 
# LAYER pactive
#   TYPE	MASTERSLICE ;
# END pactive

# LAYER poly
#   TYPE	MASTERSLICE ;
# END poly
# 
# LAYER cc
#   TYPE	CUT ;
#   SPACING	0.9 ;
# END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.5  ;
  OFFSET	1.5 ;
  WIDTH		0.9 ;
  SPACING	0.6 ;
  RESISTANCE	RPERSQ 0.085 ;
  CAPACITANCE	CPERSQDIST 3.2e-05 ;
END metal1

LAYER via1
  TYPE	CUT ;
  WIDTH 0.5 ;
  SPACING 0.6 ;
  ENCLOSURE BELOW 0.2 0.2 ;
  ENCLOSURE ABOVE 0.2 0.2 ;
  RESISTANCE 1.0 ;
#  SPACING	1.1
#    CENTERTOCENTER ;
#  PROPERTY contactResistance 1.0 ;
END via1

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		1.6 ;
  OFFSET	0.0 ;
  WIDTH		0.9 ;
  SPACING	0.7 ;
  RESISTANCE	RPERSQ 0.085 ;
  CAPACITANCE	CPERSQDIST 1.6e-05 ;
END metal2

LAYER via2
  TYPE	CUT ;
  WIDTH 0.5 ;
  SPACING 0.8 ;
  ENCLOSURE BELOW 0.2 0.2 ;
  ENCLOSURE ABOVE 0.2 0.2 ;
  RESISTANCE 1.0 ;
#  SPACING	1.3 
#    CENTERTOCENTER ;
#  PROPERTY contactResistance 1.0 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.6 ;
  OFFSET	1.5 ;
  WIDTH		0.9 ;
  SPACING	0.7 ;
  RESISTANCE	RPERSQ 0.040 ;
  CAPACITANCE	CPERSQDIST 1e-05 ;
END metal3

# SPACING
#   SAMENET cc  via	0.150 ;
#   SAMENET via  via2	0.150 ;
# END SPACING

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER via1 ;
    RECT -0.250 -0.250 0.250 0.250 ;
  LAYER metal2 ;
    RECT -0.450 -0.450 0.450 0.450 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER via2 ;
    RECT -0.250 -0.250 0.250 0.250 ;
  LAYER metal3 ;
    RECT -0.450 -0.450 0.450 0.450 ;
END M3_M2

VIARULE viagen21 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER metal2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via1 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1.1 BY 1.1 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER metal3 ;
    ENCLOSURE 0.2 0.2 ;
  LAYER via2 ;
    RECT -0.25 -0.25 0.25 0.25 ;
    SPACING 1.3 BY 1.3 ;
END viagen32

# VIARULE viagen21 GENERATE
#   LAYER metal1 ;
#     WIDTH 1.2 TO 120 ;
#     DIRECTION VERTICAL ;
#     OVERHANG 0.2 ;
#   LAYER metal2 ;
#     WIDTH 1.2 TO 120 ;
#     DIRECTION HORIZONTAL ;
#     OVERHANG 0.2 ;
#   LAYER via1 ;
#     RECT -0.25 -0.25 0.25 0.25 ;
#     SPACING 1.1 BY 1.1 ;
# END viagen21
# 
# VIARULE viagen32 GENERATE
#   LAYER metal3 ;
#     WIDTH 1.8 TO 180 ;
#     DIRECTION VERTICAL ;
#     OVERHANG 0.2 ;
#   LAYER metal2 ;
#     WIDTH 1.2 TO 120 ;
#     DIRECTION HORIZONTAL ;
#     OVERHANG 0.2 ;
#   LAYER via2 ;
#     RECT -0.25 -0.25 0.25 0.25 ;
#     SPACING 1.3 BY 1.3 ;
# END viagen32

# VIARULE TURN1 GENERATE
#   LAYER metal1 ;
#     DIRECTION VERTICAL ;
#   LAYER metal1 ;
#     DIRECTION HORIZONTAL ;
# END TURN1
# 
# VIARULE TURN2 GENERATE
#   LAYER metal2 ;
#     DIRECTION HORIZONTAL ;
#   LAYER metal2 ;
#     DIRECTION VERTICAL ;
# END TURN2
# 
# VIARULE TURN3 GENERATE
#   LAYER metal3 ;
#     DIRECTION VERTICAL ;
#   LAYER metal3 ;
#     DIRECTION HORIZONTAL ;
# END TURN3

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	1.500 BY 14.400 ;
END  core

END LIBRARY
