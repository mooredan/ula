module decap5 ();
endmodule
