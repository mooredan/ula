magic
tech amic5n
timestamp 1625245169
<< nwell >>
rect -130 550 1330 1495
rect 105 150 1095 550
<< polysilicon >>
rect 105 1240 1095 1290
rect 105 1220 225 1240
rect 105 1170 125 1220
rect 175 1170 225 1220
rect 975 1220 1095 1240
rect 105 1120 225 1170
rect 975 1170 1025 1220
rect 1075 1170 1095 1220
rect 105 1070 125 1120
rect 175 1070 225 1120
rect 975 1120 1095 1170
rect 975 1070 1025 1120
rect 1075 1070 1095 1120
rect 105 1020 225 1070
rect 975 1020 1095 1070
rect 105 970 125 1020
rect 175 970 225 1020
rect 105 920 225 970
rect 975 970 1025 1020
rect 1075 970 1095 1020
rect 105 870 125 920
rect 175 870 225 920
rect 975 920 1095 970
rect 105 820 225 870
rect 975 870 1025 920
rect 1075 870 1095 920
rect 105 770 125 820
rect 175 770 225 820
rect 975 820 1095 870
rect 105 720 225 770
rect 975 770 1025 820
rect 1075 770 1095 820
rect 105 670 125 720
rect 175 670 225 720
rect 975 720 1095 770
rect 105 620 225 670
rect 975 670 1025 720
rect 1075 670 1095 720
rect 105 570 125 620
rect 175 570 225 620
rect 975 620 1095 670
rect 105 520 225 570
rect 975 570 1025 620
rect 1075 570 1095 620
rect 975 520 1095 570
rect 105 470 125 520
rect 175 470 225 520
rect 975 470 1025 520
rect 1075 470 1095 520
rect 105 420 225 470
rect 105 370 125 420
rect 175 370 225 420
rect 975 420 1095 470
rect 105 320 225 370
rect 975 370 1025 420
rect 1075 370 1095 420
rect 105 270 125 320
rect 175 270 225 320
rect 975 320 1095 370
rect 105 220 225 270
rect 975 270 1025 320
rect 1075 270 1095 320
rect 105 170 125 220
rect 175 200 225 220
rect 975 220 1095 270
rect 975 200 1025 220
rect 175 170 1025 200
rect 1075 170 1095 220
rect 105 150 1095 170
<< polycontact >>
rect 125 1170 175 1220
rect 1025 1170 1075 1220
rect 125 1070 175 1120
rect 1025 1070 1075 1120
rect 125 970 175 1020
rect 1025 970 1075 1020
rect 125 870 175 920
rect 1025 870 1075 920
rect 125 770 175 820
rect 1025 770 1075 820
rect 125 670 175 720
rect 1025 670 1075 720
rect 125 570 175 620
rect 1025 570 1075 620
rect 125 470 175 520
rect 1025 470 1075 520
rect 125 370 175 420
rect 1025 370 1075 420
rect 125 270 175 320
rect 1025 270 1075 320
rect 125 170 175 220
rect 1025 170 1075 220
<< poly2cap >>
rect 225 1180 975 1240
rect 225 1130 275 1180
rect 325 1130 400 1180
rect 450 1130 515 1180
rect 565 1130 640 1180
rect 690 1130 755 1180
rect 805 1130 875 1180
rect 925 1130 975 1180
rect 225 1070 975 1130
rect 225 1020 275 1070
rect 325 1020 400 1070
rect 450 1020 515 1070
rect 565 1020 640 1070
rect 690 1020 755 1070
rect 805 1020 875 1070
rect 925 1020 975 1070
rect 225 960 975 1020
rect 225 910 275 960
rect 325 910 400 960
rect 450 910 515 960
rect 565 910 640 960
rect 690 910 755 960
rect 805 910 875 960
rect 925 910 975 960
rect 225 850 975 910
rect 225 800 275 850
rect 325 800 400 850
rect 450 800 515 850
rect 565 800 640 850
rect 690 800 755 850
rect 805 800 875 850
rect 925 800 975 850
rect 225 740 975 800
rect 225 690 275 740
rect 325 690 400 740
rect 450 690 515 740
rect 565 690 640 740
rect 690 690 755 740
rect 805 690 875 740
rect 925 690 975 740
rect 225 630 975 690
rect 225 580 275 630
rect 325 580 400 630
rect 450 580 515 630
rect 565 580 640 630
rect 690 580 755 630
rect 805 580 875 630
rect 925 580 975 630
rect 225 520 975 580
rect 225 470 275 520
rect 325 470 400 520
rect 450 470 515 520
rect 565 470 640 520
rect 690 470 755 520
rect 805 470 875 520
rect 925 470 975 520
rect 225 410 975 470
rect 225 360 275 410
rect 325 360 400 410
rect 450 360 515 410
rect 565 360 640 410
rect 690 360 755 410
rect 805 360 875 410
rect 925 360 975 410
rect 225 300 975 360
rect 225 250 275 300
rect 325 250 400 300
rect 450 250 515 300
rect 565 250 640 300
rect 690 250 755 300
rect 805 250 875 300
rect 925 250 975 300
rect 225 200 975 250
<< poly2capcontact >>
rect 275 1130 325 1180
rect 400 1130 450 1180
rect 515 1130 565 1180
rect 640 1130 690 1180
rect 755 1130 805 1180
rect 875 1130 925 1180
rect 275 1020 325 1070
rect 400 1020 450 1070
rect 515 1020 565 1070
rect 640 1020 690 1070
rect 755 1020 805 1070
rect 875 1020 925 1070
rect 275 910 325 960
rect 400 910 450 960
rect 515 910 565 960
rect 640 910 690 960
rect 755 910 805 960
rect 875 910 925 960
rect 275 800 325 850
rect 400 800 450 850
rect 515 800 565 850
rect 640 800 690 850
rect 755 800 805 850
rect 875 800 925 850
rect 275 690 325 740
rect 400 690 450 740
rect 515 690 565 740
rect 640 690 690 740
rect 755 690 805 740
rect 875 690 925 740
rect 275 580 325 630
rect 400 580 450 630
rect 515 580 565 630
rect 640 580 690 630
rect 755 580 805 630
rect 875 580 925 630
rect 275 470 325 520
rect 400 470 450 520
rect 515 470 565 520
rect 640 470 690 520
rect 755 470 805 520
rect 875 470 925 520
rect 275 360 325 410
rect 400 360 450 410
rect 515 360 565 410
rect 640 360 690 410
rect 755 360 805 410
rect 875 360 925 410
rect 275 250 325 300
rect 400 250 450 300
rect 515 250 565 300
rect 640 250 690 300
rect 755 250 805 300
rect 875 250 925 300
<< metal1 >>
rect 0 1395 1200 1485
rect 165 1305 1035 1395
rect 105 1220 195 1240
rect 105 1170 125 1220
rect 175 1170 195 1220
rect 105 1120 195 1170
rect 105 1070 125 1120
rect 175 1070 195 1120
rect 105 1020 195 1070
rect 105 970 125 1020
rect 175 970 195 1020
rect 105 920 195 970
rect 105 870 125 920
rect 175 870 195 920
rect 105 820 195 870
rect 105 770 125 820
rect 175 770 195 820
rect 105 720 195 770
rect 105 670 125 720
rect 175 670 195 720
rect 105 620 195 670
rect 105 570 125 620
rect 175 570 195 620
rect 105 520 195 570
rect 105 470 125 520
rect 175 470 195 520
rect 105 420 195 470
rect 105 370 125 420
rect 175 370 195 420
rect 105 320 195 370
rect 105 270 125 320
rect 175 270 195 320
rect 105 220 195 270
rect 255 1180 945 1305
rect 255 1130 275 1180
rect 325 1130 400 1180
rect 450 1130 515 1180
rect 565 1130 640 1180
rect 690 1130 755 1180
rect 805 1130 875 1180
rect 925 1130 945 1180
rect 255 1070 945 1130
rect 255 1020 275 1070
rect 325 1020 400 1070
rect 450 1020 515 1070
rect 565 1020 640 1070
rect 690 1020 755 1070
rect 805 1020 875 1070
rect 925 1020 945 1070
rect 255 960 945 1020
rect 255 910 275 960
rect 325 910 400 960
rect 450 910 515 960
rect 565 910 640 960
rect 690 910 755 960
rect 805 910 875 960
rect 925 910 945 960
rect 255 850 945 910
rect 255 800 275 850
rect 325 800 400 850
rect 450 800 515 850
rect 565 800 640 850
rect 690 800 755 850
rect 805 800 875 850
rect 925 800 945 850
rect 255 740 945 800
rect 255 690 275 740
rect 325 690 400 740
rect 450 690 515 740
rect 565 690 640 740
rect 690 690 755 740
rect 805 690 875 740
rect 925 690 945 740
rect 255 630 945 690
rect 255 580 275 630
rect 325 580 400 630
rect 450 580 515 630
rect 565 580 640 630
rect 690 580 755 630
rect 805 580 875 630
rect 925 580 945 630
rect 255 520 945 580
rect 255 470 275 520
rect 325 470 400 520
rect 450 470 515 520
rect 565 470 640 520
rect 690 470 755 520
rect 805 470 875 520
rect 925 470 945 520
rect 255 410 945 470
rect 255 360 275 410
rect 325 360 400 410
rect 450 360 515 410
rect 565 360 640 410
rect 690 360 755 410
rect 805 360 875 410
rect 925 360 945 410
rect 255 300 945 360
rect 255 250 275 300
rect 325 250 400 300
rect 450 250 515 300
rect 565 250 640 300
rect 690 250 755 300
rect 805 250 875 300
rect 925 250 945 300
rect 255 230 945 250
rect 1005 1220 1095 1240
rect 1005 1170 1025 1220
rect 1075 1170 1095 1220
rect 1005 1120 1095 1170
rect 1005 1070 1025 1120
rect 1075 1070 1095 1120
rect 1005 1020 1095 1070
rect 1005 970 1025 1020
rect 1075 970 1095 1020
rect 1005 920 1095 970
rect 1005 870 1025 920
rect 1075 870 1095 920
rect 1005 820 1095 870
rect 1005 770 1025 820
rect 1075 770 1095 820
rect 1005 720 1095 770
rect 1005 670 1025 720
rect 1075 670 1095 720
rect 1005 620 1095 670
rect 1005 570 1025 620
rect 1075 570 1095 620
rect 1005 520 1095 570
rect 1005 470 1025 520
rect 1075 470 1095 520
rect 1005 420 1095 470
rect 1005 370 1025 420
rect 1075 370 1095 420
rect 1005 320 1095 370
rect 1005 270 1025 320
rect 1075 270 1095 320
rect 105 170 125 220
rect 175 170 195 220
rect 105 150 195 170
rect 1005 220 1095 270
rect 1005 170 1025 220
rect 1075 170 1095 220
rect 1005 150 1095 170
rect 105 45 1095 150
rect 0 -45 1200 45
<< labels >>
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 0 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 1 ne
flabel nwell 5 580 5 580 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFsite core
string LEFclass CORE
string FIXED_BBOX 0 0 1200 1440
string LEFsymmetry X Y
<< end >>
