`celldefine
module decap7 ();
endmodule
`endcelldefine
