magic
tech amic5n
timestamp 1608317707
<< poly2 >>
rect -600 -330 510 480
<< poly2contact >>
rect -175 5 -125 115
<< metal1 >>
rect -450 -210 420 390
<< checkpaint >>
rect -610 -340 520 490
<< end >>
