magic
tech amic5n
timestamp 1624142612
<< nwell >>
rect -130 550 1180 1495
<< ntransistor >>
rect 165 95 225 400
rect 800 95 860 400
<< ptransistor >>
rect 165 700 225 1345
rect 355 700 415 1345
rect 610 700 670 1345
rect 800 700 860 1345
<< nselect >>
rect -10 295 1060 430
rect -10 100 400 295
rect 630 100 1060 295
rect -10 0 1060 100
<< pselect >>
rect -10 670 1060 1440
rect 400 100 630 295
<< ndiffusion >>
rect 45 370 165 400
rect 45 320 75 370
rect 125 320 165 370
rect 45 175 165 320
rect 45 125 75 175
rect 125 125 165 175
rect 45 95 165 125
rect 225 370 345 400
rect 225 320 265 370
rect 315 320 345 370
rect 225 175 345 320
rect 680 370 800 400
rect 680 320 710 370
rect 760 320 800 370
rect 225 125 265 175
rect 315 125 345 175
rect 680 175 800 320
rect 225 95 345 125
rect 680 125 710 175
rect 760 125 800 175
rect 680 95 800 125
rect 860 355 980 400
rect 860 305 900 355
rect 950 305 980 355
rect 860 175 980 305
rect 860 125 900 175
rect 950 125 980 175
rect 860 95 980 125
<< pdiffusion >>
rect 45 1315 165 1345
rect 45 1265 75 1315
rect 125 1265 165 1315
rect 45 1200 165 1265
rect 45 1150 75 1200
rect 125 1150 165 1200
rect 45 1065 165 1150
rect 45 1015 75 1065
rect 125 1015 165 1065
rect 45 945 165 1015
rect 45 895 75 945
rect 125 895 165 945
rect 45 825 165 895
rect 45 775 75 825
rect 125 775 165 825
rect 45 700 165 775
rect 225 1315 355 1345
rect 225 1265 265 1315
rect 315 1265 355 1315
rect 225 1215 355 1265
rect 225 1165 265 1215
rect 315 1165 355 1215
rect 225 1115 355 1165
rect 225 1065 265 1115
rect 315 1065 355 1115
rect 225 985 355 1065
rect 225 935 265 985
rect 315 935 355 985
rect 225 700 355 935
rect 415 1315 610 1345
rect 415 1265 475 1315
rect 525 1265 610 1315
rect 415 1200 610 1265
rect 415 1150 475 1200
rect 525 1150 610 1200
rect 415 1065 610 1150
rect 415 1015 475 1065
rect 525 1015 610 1065
rect 415 945 610 1015
rect 415 895 475 945
rect 525 895 610 945
rect 415 825 610 895
rect 415 775 475 825
rect 525 775 610 825
rect 415 700 610 775
rect 670 1155 800 1345
rect 670 1105 710 1155
rect 760 1105 800 1155
rect 670 1015 800 1105
rect 670 965 710 1015
rect 760 965 800 1015
rect 670 915 800 965
rect 670 865 710 915
rect 760 865 800 915
rect 670 815 800 865
rect 670 765 710 815
rect 760 765 800 815
rect 670 700 800 765
rect 860 1315 980 1345
rect 860 1265 900 1315
rect 950 1265 980 1315
rect 860 1180 980 1265
rect 860 1130 900 1180
rect 950 1130 980 1180
rect 860 1080 980 1130
rect 860 1030 900 1080
rect 950 1030 980 1080
rect 860 980 980 1030
rect 860 930 900 980
rect 950 930 980 980
rect 860 880 980 930
rect 860 830 900 880
rect 950 830 980 880
rect 860 780 980 830
rect 860 730 900 780
rect 950 730 980 780
rect 860 700 980 730
<< psubstratepdiff >>
rect 455 220 565 250
rect 455 170 485 220
rect 535 170 565 220
rect 455 140 565 170
<< psubstratepcontact >>
rect 485 170 535 220
<< ndcontact >>
rect 75 320 125 370
rect 75 125 125 175
rect 265 320 315 370
rect 710 320 760 370
rect 265 125 315 175
rect 710 125 760 175
rect 900 305 950 355
rect 900 125 950 175
<< pdcontact >>
rect 75 1265 125 1315
rect 75 1150 125 1200
rect 75 1015 125 1065
rect 75 895 125 945
rect 75 775 125 825
rect 265 1265 315 1315
rect 265 1165 315 1215
rect 265 1065 315 1115
rect 265 935 315 985
rect 475 1265 525 1315
rect 475 1150 525 1200
rect 475 1015 525 1065
rect 475 895 525 945
rect 475 775 525 825
rect 710 1105 760 1155
rect 710 965 760 1015
rect 710 865 760 915
rect 710 765 760 815
rect 900 1265 950 1315
rect 900 1130 950 1180
rect 900 1030 950 1080
rect 900 930 950 980
rect 900 830 950 880
rect 900 730 950 780
<< polysilicon >>
rect 165 1345 225 1410
rect 355 1345 415 1410
rect 610 1345 670 1410
rect 800 1345 860 1410
rect 165 630 225 700
rect 355 630 415 700
rect 165 610 415 630
rect 165 560 225 610
rect 275 560 415 610
rect 165 540 415 560
rect 610 560 670 700
rect 800 560 860 700
rect 610 540 1020 560
rect 165 400 225 540
rect 610 490 950 540
rect 1000 490 1020 540
rect 610 470 1020 490
rect 800 400 860 470
rect 165 30 225 95
rect 800 30 860 95
<< polycontact >>
rect 225 560 275 610
rect 950 490 1000 540
<< metal1 >>
rect 0 1395 1050 1485
rect 55 1315 145 1335
rect 55 1265 75 1315
rect 125 1265 145 1315
rect 55 1200 145 1265
rect 55 1150 75 1200
rect 125 1150 145 1200
rect 55 1065 145 1150
rect 55 1015 75 1065
rect 125 1015 145 1065
rect 55 945 145 1015
rect 55 895 75 945
rect 125 895 145 945
rect 245 1315 335 1395
rect 245 1265 265 1315
rect 315 1265 335 1315
rect 245 1215 335 1265
rect 245 1165 265 1215
rect 315 1165 335 1215
rect 245 1115 335 1165
rect 245 1065 265 1115
rect 315 1065 335 1115
rect 245 985 335 1065
rect 245 935 265 985
rect 315 935 335 985
rect 245 915 335 935
rect 455 1325 545 1335
rect 880 1325 970 1335
rect 455 1315 970 1325
rect 455 1265 475 1315
rect 525 1265 900 1315
rect 950 1265 970 1315
rect 455 1235 970 1265
rect 455 1200 545 1235
rect 455 1150 475 1200
rect 525 1150 545 1200
rect 880 1180 970 1235
rect 455 1065 545 1150
rect 455 1015 475 1065
rect 525 1015 545 1065
rect 455 945 545 1015
rect 55 845 145 895
rect 455 895 475 945
rect 525 895 545 945
rect 455 845 545 895
rect 55 825 545 845
rect 55 775 75 825
rect 125 775 475 825
rect 525 775 545 825
rect 55 755 545 775
rect 690 1155 780 1175
rect 690 1105 710 1155
rect 760 1105 780 1155
rect 690 1015 780 1105
rect 690 965 710 1015
rect 760 965 780 1015
rect 690 915 780 965
rect 690 865 710 915
rect 760 865 780 915
rect 690 815 780 865
rect 690 765 710 815
rect 760 765 780 815
rect 205 610 295 685
rect 205 560 225 610
rect 275 560 295 610
rect 205 540 295 560
rect 690 390 780 765
rect 880 1130 900 1180
rect 950 1130 970 1180
rect 880 1080 970 1130
rect 880 1030 900 1080
rect 950 1030 970 1080
rect 880 980 970 1030
rect 880 930 900 980
rect 950 930 970 980
rect 880 880 970 930
rect 880 830 900 880
rect 950 830 970 880
rect 880 780 970 830
rect 880 730 900 780
rect 950 730 970 780
rect 880 710 970 730
rect 930 540 1020 560
rect 930 490 950 540
rect 1000 490 1020 540
rect 930 435 1020 490
rect 55 370 145 390
rect 55 320 75 370
rect 125 320 145 370
rect 55 175 145 320
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 245 370 780 390
rect 245 320 265 370
rect 315 320 710 370
rect 760 320 780 370
rect 245 300 780 320
rect 245 175 335 300
rect 245 125 265 175
rect 315 125 335 175
rect 245 105 335 125
rect 465 220 555 240
rect 465 170 485 220
rect 535 170 555 220
rect 465 45 555 170
rect 690 175 780 300
rect 690 125 710 175
rect 760 125 780 175
rect 690 105 780 125
rect 880 355 970 375
rect 880 305 900 355
rect 950 305 970 355
rect 880 175 970 305
rect 880 125 900 175
rect 950 125 970 175
rect 880 45 970 125
rect 0 -45 1050 45
<< labels >>
flabel metal1 s 720 1045 720 1045 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 950 480 950 480 2 FreeSans 400 0 0 0 b
port 2 ne
flabel metal1 s 120 1415 120 1415 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel nwell 55 600 55 600 8 FreeSans 400 180 0 0 vdd
flabel metal1 s 225 550 225 550 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 4 ne
<< end >>
