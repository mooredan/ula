magic
tech scmos
timestamp 1511590936
<< nwell >>
rect 26 24 42 65
<< nselect >>
rect 30 24 38 61
<< pselect >>
rect 30 2 38 24
<< psubstratepdiff >>
rect 32 4 36 21
<< nsubstratendiff >>
rect 32 27 36 59
<< genericcontact >>
rect 33 56 35 58
rect 33 51 35 53
rect 33 46 35 48
rect 33 41 35 43
rect 33 36 35 38
rect 33 31 35 33
rect 33 18 35 20
rect 33 13 35 15
rect 33 8 35 10
<< metal1 >>
rect 32 30 36 63
rect 32 0 36 21
<< bb >>
rect 27 0 41 63
use INV_B  INV_B_0
timestamp 1511585079
transform 1 0 1 0 1 0
box -1 0 27 65
use INV_B  INV_B_1
timestamp 1511585079
transform 1 0 41 0 1 0
box -1 0 27 65
<< end >>
