magic
tech scmos
timestamp 1591761821
<< nwell >>
rect -1 24 34 65
rect 43 29 75 81
<< nselect >>
rect 6 46 30 61
rect 6 2 27 19
rect 47 2 71 25
<< pselect >>
rect 6 30 30 46
rect 47 33 71 77
rect 54 32 56 33
<< ntransistor >>
rect 13 4 15 17
rect 18 4 20 17
rect 54 4 56 23
rect 62 4 64 23
<< ptransistor >>
rect 13 32 15 43
rect 21 32 23 43
rect 54 35 56 75
rect 62 35 64 75
<< ndiffusion >>
rect 8 4 13 17
rect 15 4 18 17
rect 20 4 25 17
rect 49 4 54 23
rect 56 4 62 23
rect 64 4 69 23
<< pdiffusion >>
rect 8 32 13 43
rect 15 32 21 43
rect 23 32 28 43
rect 49 35 54 75
rect 56 35 62 75
rect 64 35 69 75
<< nsubstratendiff >>
rect 15 53 21 58
<< polysilicon >>
rect 54 75 56 77
rect 62 75 64 77
rect 13 43 15 45
rect 21 43 23 45
rect 54 32 56 35
rect 13 24 15 32
rect 8 18 15 24
rect 21 24 23 32
rect 49 26 56 32
rect 21 20 28 24
rect 54 23 56 26
rect 62 32 64 35
rect 62 26 69 32
rect 62 23 64 26
rect 13 17 15 18
rect 18 18 28 20
rect 18 17 20 18
rect 13 2 15 4
rect 18 2 20 4
rect 54 2 56 4
rect 62 2 64 4
<< genericcontact >>
rect 50 72 52 74
rect 58 70 60 72
rect 66 70 68 72
rect 50 66 52 68
rect 58 65 60 67
rect 66 65 68 67
rect 50 61 52 63
rect 58 59 60 61
rect 66 59 68 61
rect 17 55 19 57
rect 50 56 52 58
rect 50 51 52 53
rect 58 52 60 54
rect 66 53 68 55
rect 50 46 52 48
rect 58 46 60 48
rect 66 47 68 49
rect 9 39 11 41
rect 17 40 19 42
rect 50 41 52 43
rect 58 41 60 43
rect 66 41 68 43
rect 25 39 27 41
rect 50 36 52 38
rect 58 36 60 38
rect 66 36 68 38
rect 9 34 11 36
rect 17 34 19 36
rect 25 34 27 36
rect 51 28 53 30
rect 65 28 67 30
rect 10 20 12 22
rect 24 20 26 22
rect 50 20 52 22
rect 66 20 68 22
rect 50 15 52 17
rect 9 13 11 15
rect 22 13 24 15
rect 66 14 68 16
rect 50 10 52 12
rect 9 6 11 8
rect 22 7 24 9
rect 66 7 68 9
rect 50 5 52 7
<< metal1 >>
rect 47 76 71 79
rect 5 60 28 63
rect 8 33 12 60
rect 16 54 20 60
rect 9 19 13 23
rect 16 16 20 43
rect 24 33 28 60
rect 49 35 53 76
rect 50 27 54 31
rect 57 23 61 73
rect 65 35 69 76
rect 64 27 68 31
rect 23 19 27 23
rect 8 3 12 16
rect 16 12 25 16
rect 21 6 25 12
rect 49 3 53 23
rect 57 19 69 23
rect 65 6 69 19
rect 5 0 28 3
rect 47 0 71 3
<< bb >>
rect 0 0 33 63
<< labels >>
rlabel metal1 16 12 20 43 0 z
port 1 new
rlabel metal1 21 6 25 16 0 z
port 1 e
rlabel metal1 9 19 13 23 0 a
port 2 nw
rlabel metal1 23 19 27 23 0 b
port 3 ne
rlabel metal1 5 60 28 63 0 Vdd
port 4 new
rlabel metal1 5 0 28 3 0 Gnd
port 5 sew
rlabel ndiffusion 16 8 16 8 2 x1
rlabel nwell 3 25 3 25 2 Vdd
rlabel nwell 47 31 47 31 2 vdd
rlabel metal1 s 48 1 48 1 2 vss
port 5 ne
rlabel metal1 s 48 77 48 77 2 vdd
port 4 ne
rlabel metal1 s 52 29 52 29 2 a
port 2 ne
rlabel metal1 s 59 26 59 26 2 z
port 1 ne
rlabel ndiffusion s 59 11 59 11 2 x1
rlabel metal1 s 66 29 66 29 2 b
port 3 ne
<< end >>
