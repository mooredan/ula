`celldefine
module or2_b (z, a, b);
  output z;
  input  a;
  input  b;

  or G1 (z, a, b);
endmodule
`endcelldefine
