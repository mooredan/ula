`celldefine
module inv_b (z, a);
  output z;
  input  a;

  not G1 (z, a);
endmodule
`endcelldefine
