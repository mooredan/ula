magic
tech scmos
timestamp 1606089699
<< error_p >>
rect -101 -3 -100 9
<< nselect >>
rect -14 -30 29 -14
<< electrode >>
rect -96 -3 -85 9
rect -82 -3 -72 9
rect -14 -42 4 -29
rect 70 -40 81 52
<< electrodecap >>
rect -96 19 -85 31
rect -82 19 -69 31
rect -18 8 -5 19
rect -28 1 -5 8
rect -18 -9 -5 1
rect -2 -9 8 19
<< genericpoly2contact >>
rect -1 16 1 18
rect -16 14 -14 16
rect -1 11 1 13
rect -16 9 -14 11
rect -13 -41 -11 -39
rect 1 -41 3 -39
<< ntransistor >>
rect -12 -23 27 -21
<< ndiffusion >>
rect -12 -21 27 -16
rect -12 -28 27 -23
<< ndcontact >>
rect 62 39 69 45
<< pdcontact >>
rect 62 21 69 27
<< psubstratepdiff >>
rect 65 -40 69 -36
<< psubstratepcontact >>
rect 62 5 69 11
<< nsubstratencontact >>
rect 62 -11 69 -5
<< polysilicon >>
rect -98 31 -67 33
rect -98 19 -96 31
rect -85 19 -82 31
rect -69 19 -67 31
rect -98 17 -67 19
rect -20 19 13 21
rect -20 10 -18 19
rect -111 -3 -100 9
rect -30 8 -18 10
rect -30 1 -28 8
rect -30 -1 -18 1
rect -20 -9 -18 -1
rect -5 -9 -2 19
rect 8 -9 13 19
rect -20 -11 13 -9
rect 30 -21 34 -20
rect -14 -23 -12 -21
rect 27 -23 34 -21
rect 30 -24 34 -23
<< polycontact >>
rect 58 -22 65 -16
<< genericcontact >>
rect 10 16 12 18
rect 10 11 12 13
rect 10 6 12 8
rect -11 -19 -9 -17
rect -6 -19 -4 -17
rect -1 -19 1 -17
rect 4 -19 6 -17
rect 9 -19 11 -17
rect 14 -19 16 -17
rect 19 -19 21 -17
rect 24 -19 26 -17
rect 31 -23 33 -21
rect 14 -27 16 -25
rect 19 -27 21 -25
rect 24 -27 26 -25
rect 66 -39 68 -37
<< metal1 >>
rect -17 8 -13 17
rect -2 9 2 19
rect 9 5 13 19
rect -12 -20 27 -16
rect 30 -24 34 -20
rect 13 -28 27 -24
rect -14 -42 -10 -38
rect 0 -42 4 -38
rect 65 -40 69 -36
<< end >>
