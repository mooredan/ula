magic
tech scmos
timestamp 1591541005
<< nwell >>
rect -1 29 15 81
<< metal1 >>
rect 5 76 9 79
rect 5 69 8 73
rect 5 62 8 66
rect 5 55 8 59
rect 5 48 8 52
rect 5 41 8 45
rect 5 34 8 38
rect 5 27 8 31
rect 5 20 8 24
rect 5 13 8 17
rect 5 6 8 10
rect 5 0 9 3
rect -2 -10 2 -3
rect 5 -10 9 -3
rect 12 -10 16 -3
<< bb >>
rect 0 0 14 79
<< labels >>
rlabel metal1 5 0 5 0 2 Gnd
port 3 ne
rlabel nwell 5 30 5 30 2 Vdd
rlabel metal1 5 76 5 76 2 Vdd
port 2 ne
<< end >>
