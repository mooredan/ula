magic
tech amic5n
timestamp 1606481034
<< error_p >>
rect 10730 -10 11320 100
<< nwell >>
rect 6670 1890 7560 2500
rect 2880 80 3500 570
rect 5340 30 6110 930
rect 6900 -2200 8130 -1700
rect 8720 -1890 8970 -1640
rect 9370 -1810 10140 -1240
<< nselect >>
rect 4900 1890 5200 2170
rect 5300 1980 5390 2070
rect 6820 2050 7120 2330
rect 7220 2140 7310 2230
rect 7470 1110 7840 1470
rect 5790 580 5990 810
rect 4410 330 4760 560
rect 4410 -100 4960 330
rect 8600 -140 8900 140
rect 9000 -50 9090 40
rect 3620 -620 3990 -260
rect 4670 -510 4940 -180
rect 5500 -530 5670 -170
rect 3760 -1080 4210 -790
rect 6900 -1580 7870 -1180
rect 7870 -2080 8110 -1740
rect 9340 -1840 9510 -1670
<< pselect >>
rect 5200 2070 5500 2170
rect 5200 1980 5300 2070
rect 5390 1980 5500 2070
rect 7120 2230 7420 2330
rect 7120 2140 7220 2230
rect 7310 2140 7420 2230
rect 7120 2050 7420 2140
rect 5200 1890 5500 1980
rect 5440 580 5790 810
rect 3000 240 3380 440
rect 4760 330 4960 560
rect 5440 150 5990 580
rect 8900 40 9200 140
rect 8900 -50 9000 40
rect 9090 -50 9200 40
rect 8900 -140 9200 -50
rect 4670 -580 4940 -510
rect 7870 -1580 8110 -1180
rect 7020 -2080 7870 -1740
rect 9350 -2310 9520 -2140
<< poly2 >>
rect 9040 740 9240 940
rect 10770 110 11130 310
rect 7330 -330 8170 -100
rect 10930 -10 11130 110
rect 8250 -330 9290 -130
rect 10930 -210 11130 -100
rect 10770 -430 11130 -210
<< poly2cap >>
rect 6910 630 7200 910
rect 7280 630 7720 910
<< ntransistor >>
rect 7500 1260 7810 1320
rect 4460 150 4930 210
rect 4700 -390 4910 -330
rect 5530 -380 5640 -320
rect 3650 -470 3960 -410
rect 3790 -980 4180 -910
<< ptransistor >>
rect 3160 280 3220 390
rect 5490 400 5960 460
<< ndiffusion >>
rect 4930 1920 5200 2140
rect 5300 1980 5390 2070
rect 7500 1320 7810 1440
rect 7500 1140 7810 1260
rect 4460 330 4760 530
rect 4460 210 4930 330
rect 4460 -70 4930 150
rect 3650 -410 3960 -290
rect 4700 -330 4910 -210
rect 5530 -320 5640 -200
rect 8630 -110 8900 110
rect 9000 -50 9090 40
rect 3650 -590 3960 -470
rect 4700 -510 4910 -390
rect 5530 -500 5640 -380
rect 3790 -910 4180 -820
rect 3790 -1050 4180 -980
rect 7060 -1550 7290 -1330
rect 7380 -1550 7810 -1330
<< pdiffusion >>
rect 7120 2080 7390 2300
rect 5490 580 5790 780
rect 3090 380 3160 390
rect 3030 290 3160 380
rect 3090 280 3160 290
rect 3220 280 3350 390
rect 5490 460 5960 580
rect 5490 180 5960 400
rect 7050 -2050 7290 -1850
rect 7380 -2050 7800 -1850
<< psubstratepdiff >>
rect 5200 2070 5470 2140
rect 5200 1980 5300 2070
rect 5390 1980 5470 2070
rect 5200 1920 5470 1980
rect 4760 330 4930 530
rect 8900 40 9170 110
rect 8900 -50 9000 40
rect 9090 -50 9170 40
rect 8900 -110 9170 -50
rect 4700 -570 4910 -510
rect 7930 -1550 8080 -1330
rect 9380 -2280 9490 -2170
<< nsubstratendiff >>
rect 6850 2080 7120 2300
rect 5790 580 5960 780
rect 9370 -1810 9480 -1700
rect 7920 -2050 8080 -1850
<< polysilicon >>
rect 7350 1320 7440 1350
rect 7350 1260 7500 1320
rect 7810 1260 7880 1320
rect 6860 910 7930 960
rect 6860 630 6910 910
rect 7200 630 7280 910
rect 7720 630 7930 910
rect 6860 580 7930 630
rect 3160 390 3220 510
rect 8280 550 8750 970
rect 5410 400 5490 460
rect 5960 400 6030 460
rect 3160 200 3220 280
rect 4380 150 4460 210
rect 4930 150 5000 210
rect -40 -40 50 50
rect 3500 -410 3590 -380
rect 4550 -330 4640 -300
rect 5380 -320 5470 -290
rect 4550 -390 4700 -330
rect 4910 -390 4980 -330
rect 5380 -380 5530 -320
rect 5640 -380 5710 -320
rect 3500 -470 3650 -410
rect 3960 -470 4030 -410
rect 2830 -850 2890 -820
rect 2830 -910 3170 -850
rect 3720 -980 3790 -910
rect 4180 -980 4250 -910
<< genericcontact >>
rect 6940 2160 6990 2210
rect 7240 2160 7290 2210
rect 5020 2000 5070 2050
rect 5320 2000 5370 2050
rect 7530 1360 7580 1410
rect 7630 1360 7680 1410
rect 7730 1360 7780 1410
rect 7370 1280 7420 1330
rect 7530 1170 7580 1220
rect 7630 1170 7680 1220
rect 7730 1170 7780 1220
rect 7390 740 7440 790
rect 7490 740 7540 790
rect 7770 750 7820 800
rect 3260 310 3310 360
rect -20 -20 30 30
rect 8720 -30 8770 20
rect 9020 -30 9070 20
rect 7350 -170 7400 -120
rect 8100 -170 8150 -120
rect 4730 -290 4780 -240
rect 4830 -290 4880 -240
rect 5560 -280 5610 -230
rect 7350 -310 7400 -260
rect 8100 -310 8150 -260
rect 3680 -370 3730 -320
rect 3780 -370 3830 -320
rect 3880 -370 3930 -320
rect 4570 -370 4620 -320
rect 5400 -360 5450 -310
rect 3520 -450 3570 -400
rect 4730 -480 4780 -430
rect 4830 -480 4880 -430
rect 5560 -470 5610 -420
rect 3680 -560 3730 -510
rect 3780 -560 3830 -510
rect 3880 -560 3930 -510
rect 9400 -1780 9450 -1730
rect 9410 -2250 9460 -2200
<< metal1 >>
rect 6830 2140 7010 2230
rect 7220 2140 7410 2230
rect 4910 1980 5090 2070
rect 5300 1980 5490 2070
rect 7350 1260 7440 1350
rect 7510 1340 7800 1430
rect 7510 1150 7800 1240
rect 7370 720 7570 810
rect 7650 630 7840 880
rect 3190 240 3340 420
rect -70 -70 90 70
rect 1230 30 1320 45
rect 250 -30 2170 30
rect 1230 -45 1320 -30
rect 8610 -50 8790 40
rect 9000 -50 9190 40
rect 1390 -110 1480 -95
rect 1180 -170 1660 -110
rect 1390 -185 1480 -170
rect 3500 -470 3590 -380
rect 3660 -390 3950 -300
rect 4550 -390 4640 -300
rect 4710 -310 4900 -220
rect 5380 -380 5470 -290
rect 5540 -300 5630 -210
rect 7330 -330 7420 -100
rect 8080 -330 8170 -100
rect 3660 -580 3950 -490
rect 4710 -500 4900 -410
rect 5540 -490 5630 -400
rect 9380 -1800 9470 -1710
rect 9390 -2270 9480 -2180
<< metal2 >>
rect 2100 -12580 4160 -4760
rect 4280 -12580 6330 -4760
<< high_resist >>
rect 10730 -100 10930 -10
rect 11130 -100 11320 -10
<< poly2_high_resist >>
rect 10930 -100 11130 -10
<< end >>
