magic
tech amic5n
timestamp 1608317708
<< ntransistor >>
rect 2250 1830 4800 1920
<< ndiffusion >>
rect 2250 1920 4800 2580
rect 2250 1440 4800 1830
<< psubstratepdiff >>
rect 2250 1020 4800 1440
<< nsubstratendiff >>
rect 3900 660 4140 840
<< polysilicon >>
rect 1710 1920 1980 2010
rect 1710 1830 2250 1920
rect 4800 1830 4860 1920
rect 1710 1740 1980 1830
<< ndcontact >>
rect 2375 2435 2425 2485
<< ndcontact >>
rect 2525 2435 2575 2485
<< ndcontact >>
rect 2675 2435 2725 2485
<< ndcontact >>
rect 2825 2435 2875 2485
<< ndcontact >>
rect 2975 2435 3025 2485
<< ndcontact >>
rect 3125 2435 3175 2485
<< ndcontact >>
rect 3275 2435 3325 2485
<< ndcontact >>
rect 3425 2435 3475 2485
<< ndcontact >>
rect 3575 2435 3625 2485
<< ndcontact >>
rect 3725 2435 3775 2485
<< ndcontact >>
rect 3875 2435 3925 2485
<< ndcontact >>
rect 4025 2435 4075 2485
<< ndcontact >>
rect 4175 2435 4225 2485
<< polycontact >>
rect 1805 1835 1855 1885
<< ndcontact >>
rect 2525 1625 2575 1675
<< ndcontact >>
rect 2675 1625 2725 1675
<< ndcontact >>
rect 2825 1625 2875 1675
<< ndcontact >>
rect 2975 1625 3025 1675
<< ndcontact >>
rect 3125 1625 3175 1675
<< ndcontact >>
rect 3275 1625 3325 1675
<< ndcontact >>
rect 3425 1625 3475 1675
<< ndcontact >>
rect 3575 1625 3625 1675
<< ndcontact >>
rect 3725 1625 3775 1675
<< ndcontact >>
rect 3875 1625 3925 1675
<< ndcontact >>
rect 4025 1625 4075 1675
<< ndcontact >>
rect 4175 1625 4225 1675
<< ndcontact >>
rect 4325 1625 4375 1675
<< ndcontact >>
rect 4475 1625 4525 1675
<< psubstratepcontact >>
rect 2615 1145 2665 1195
<< psubstratepcontact >>
rect 2915 1145 2965 1195
<< psubstratepcontact >>
rect 3215 1145 3265 1195
<< psubstratepcontact >>
rect 3515 1145 3565 1195
<< psubstratepcontact >>
rect 3815 1145 3865 1195
<< psubstratepcontact >>
rect 4115 1145 4165 1195
<< psubstratepcontact >>
rect 4415 1145 4465 1195
<< nsubstratencontact >>
rect 3995 755 4045 805
<< metal1 >>
rect 2340 2160 4740 2580
rect 1740 1770 1920 1950
rect 2460 1020 4620 1740
rect 3960 720 4110 1020
<< labels >>
flabel space  2400 840 2400 840 1 FreeSans 400 0 0 0 vss
<< checkpaint >>
rect -10 -10 4870 2590
<< end >>
