magic
tech amic5n
timestamp 1621899855
<< error_p >>
rect 45 985 75 1005
rect 125 985 155 1005
rect 45 955 155 985
rect 245 985 275 1005
rect 325 985 365 1005
rect 245 955 365 985
rect 425 985 465 1005
rect 425 955 505 985
<< nwell >>
rect -105 805 695 2455
<< ntransistor >>
rect 365 95 425 655
<< ptransistor >>
rect 365 955 425 2305
<< nselect >>
rect 0 925 200 2400
rect 200 0 590 685
<< pselect >>
rect 200 925 590 2400
rect 0 0 200 690
<< ndiffusion >>
rect 245 625 365 655
rect 245 575 275 625
rect 325 575 365 625
rect 245 475 365 575
rect 245 425 275 475
rect 325 425 365 475
rect 245 375 365 425
rect 245 325 275 375
rect 325 325 365 375
rect 245 275 365 325
rect 245 225 275 275
rect 325 225 365 275
rect 245 175 365 225
rect 245 125 275 175
rect 325 125 365 175
rect 245 95 365 125
rect 425 625 545 655
rect 425 575 465 625
rect 515 575 545 625
rect 425 475 545 575
rect 425 425 465 475
rect 515 425 545 475
rect 425 375 545 425
rect 425 325 465 375
rect 515 325 545 375
rect 425 275 545 325
rect 425 225 465 275
rect 515 225 545 275
rect 425 175 545 225
rect 425 125 465 175
rect 515 125 545 175
rect 425 95 545 125
<< pdiffusion >>
rect 245 2275 365 2305
rect 245 2225 275 2275
rect 325 2225 365 2275
rect 245 2135 365 2225
rect 245 2085 275 2135
rect 325 2085 365 2135
rect 245 2035 365 2085
rect 245 1985 275 2035
rect 325 1985 365 2035
rect 245 1935 365 1985
rect 245 1885 275 1935
rect 325 1885 365 1935
rect 245 1835 365 1885
rect 245 1785 275 1835
rect 325 1785 365 1835
rect 245 1735 365 1785
rect 245 1685 275 1735
rect 325 1685 365 1735
rect 245 1635 365 1685
rect 245 1585 275 1635
rect 325 1585 365 1635
rect 245 1535 365 1585
rect 245 1485 275 1535
rect 325 1485 365 1535
rect 245 1435 365 1485
rect 245 1385 275 1435
rect 325 1385 365 1435
rect 245 1335 365 1385
rect 245 1285 275 1335
rect 325 1285 365 1335
rect 245 1235 365 1285
rect 245 1185 275 1235
rect 325 1185 365 1235
rect 245 1135 365 1185
rect 245 1085 275 1135
rect 325 1085 365 1135
rect 245 1035 365 1085
rect 245 985 275 1035
rect 325 985 365 1035
rect 245 955 365 985
rect 425 2275 545 2305
rect 425 2225 465 2275
rect 515 2225 545 2275
rect 425 2135 545 2225
rect 425 2085 465 2135
rect 515 2085 545 2135
rect 425 2035 545 2085
rect 425 1985 465 2035
rect 515 1985 545 2035
rect 425 1935 545 1985
rect 425 1885 465 1935
rect 515 1885 545 1935
rect 425 1835 545 1885
rect 425 1785 465 1835
rect 515 1785 545 1835
rect 425 1735 545 1785
rect 425 1685 465 1735
rect 515 1685 545 1735
rect 425 1635 545 1685
rect 425 1585 465 1635
rect 515 1585 545 1635
rect 425 1535 545 1585
rect 425 1485 465 1535
rect 515 1485 545 1535
rect 425 1435 545 1485
rect 425 1385 465 1435
rect 515 1385 545 1435
rect 425 1335 545 1385
rect 425 1285 465 1335
rect 515 1285 545 1335
rect 425 1235 545 1285
rect 425 1185 465 1235
rect 515 1185 545 1235
rect 425 1135 545 1185
rect 425 1085 465 1135
rect 515 1085 545 1135
rect 425 1035 545 1085
rect 425 985 465 1035
rect 515 985 545 1035
rect 425 955 545 985
<< psubstratepdiff >>
rect 45 575 155 655
rect 45 525 75 575
rect 125 525 155 575
rect 45 475 155 525
rect 45 425 75 475
rect 125 425 155 475
rect 45 375 155 425
rect 45 325 75 375
rect 125 325 155 375
rect 45 275 155 325
rect 45 225 75 275
rect 125 225 155 275
rect 45 175 155 225
rect 45 125 75 175
rect 125 125 155 175
rect 45 95 155 125
<< nsubstratendiff >>
rect 45 2235 155 2305
rect 45 2185 75 2235
rect 125 2185 155 2235
rect 45 2135 155 2185
rect 45 2085 75 2135
rect 125 2085 155 2135
rect 45 2035 155 2085
rect 45 1985 75 2035
rect 125 1985 155 2035
rect 45 1935 155 1985
rect 45 1885 75 1935
rect 125 1885 155 1935
rect 45 1835 155 1885
rect 45 1785 75 1835
rect 125 1785 155 1835
rect 45 1735 155 1785
rect 45 1685 75 1735
rect 125 1685 155 1735
rect 45 1635 155 1685
rect 45 1585 75 1635
rect 125 1585 155 1635
rect 45 1535 155 1585
rect 45 1485 75 1535
rect 125 1485 155 1535
rect 45 1435 155 1485
rect 45 1385 75 1435
rect 125 1385 155 1435
rect 45 1335 155 1385
rect 45 1285 75 1335
rect 125 1285 155 1335
rect 45 1235 155 1285
rect 45 1185 75 1235
rect 125 1185 155 1235
rect 45 1135 155 1185
rect 45 1085 75 1135
rect 125 1085 155 1135
rect 45 1035 155 1085
rect 45 985 75 1035
rect 125 985 155 1035
rect 45 955 155 985
<< nsubstratencontact >>
rect 75 2185 125 2235
rect 75 2085 125 2135
rect 75 1985 125 2035
rect 75 1885 125 1935
rect 75 1785 125 1835
rect 75 1685 125 1735
rect 75 1585 125 1635
rect 75 1485 125 1535
rect 75 1385 125 1435
rect 75 1285 125 1335
rect 75 1185 125 1235
rect 75 1085 125 1135
rect 75 985 125 1035
<< psubstratepcontact >>
rect 75 525 125 575
rect 75 425 125 475
rect 75 325 125 375
rect 75 225 125 275
rect 75 125 125 175
<< ndcontact >>
rect 275 575 325 625
rect 275 425 325 475
rect 275 325 325 375
rect 275 225 325 275
rect 275 125 325 175
rect 465 575 515 625
rect 465 425 515 475
rect 465 325 515 375
rect 465 225 515 275
rect 465 125 515 175
<< pdcontact >>
rect 275 2225 325 2275
rect 275 2085 325 2135
rect 275 1985 325 2035
rect 275 1885 325 1935
rect 275 1785 325 1835
rect 275 1685 325 1735
rect 275 1585 325 1635
rect 275 1485 325 1535
rect 275 1385 325 1435
rect 275 1285 325 1335
rect 275 1185 325 1235
rect 275 1085 325 1135
rect 275 985 325 1035
rect 465 2225 515 2275
rect 465 2085 515 2135
rect 465 1985 515 2035
rect 465 1885 515 1935
rect 465 1785 515 1835
rect 465 1685 515 1735
rect 465 1585 515 1635
rect 465 1485 515 1535
rect 465 1385 515 1435
rect 465 1285 515 1335
rect 465 1185 515 1235
rect 465 1085 515 1135
rect 465 985 515 1035
<< polysilicon >>
rect 365 2305 425 2370
rect 365 845 425 955
rect 255 825 425 845
rect 255 775 275 825
rect 325 775 425 825
rect 255 755 425 775
rect 365 655 425 755
rect 365 30 425 95
<< polycontact >>
rect 275 775 325 825
<< metal1 >>
rect 0 2355 590 2445
rect 55 2235 145 2355
rect 55 2185 75 2235
rect 125 2185 145 2235
rect 55 2135 145 2185
rect 55 2085 75 2135
rect 125 2085 145 2135
rect 55 2035 145 2085
rect 55 1985 75 2035
rect 125 1985 145 2035
rect 55 1935 145 1985
rect 55 1885 75 1935
rect 125 1885 145 1935
rect 55 1835 145 1885
rect 55 1785 75 1835
rect 125 1785 145 1835
rect 55 1735 145 1785
rect 55 1685 75 1735
rect 125 1685 145 1735
rect 55 1635 145 1685
rect 55 1585 75 1635
rect 125 1585 145 1635
rect 55 1535 145 1585
rect 55 1485 75 1535
rect 125 1485 145 1535
rect 55 1435 145 1485
rect 55 1385 75 1435
rect 125 1385 145 1435
rect 55 1335 145 1385
rect 55 1285 75 1335
rect 125 1285 145 1335
rect 55 1235 145 1285
rect 55 1185 75 1235
rect 125 1185 145 1235
rect 55 1135 145 1185
rect 55 1085 75 1135
rect 125 1085 145 1135
rect 55 1035 145 1085
rect 55 985 75 1035
rect 125 985 145 1035
rect 55 965 145 985
rect 255 2275 345 2355
rect 255 2225 275 2275
rect 325 2225 345 2275
rect 255 2135 345 2225
rect 255 2085 275 2135
rect 325 2085 345 2135
rect 255 2035 345 2085
rect 255 1985 275 2035
rect 325 1985 345 2035
rect 255 1935 345 1985
rect 255 1885 275 1935
rect 325 1885 345 1935
rect 255 1835 345 1885
rect 255 1785 275 1835
rect 325 1785 345 1835
rect 255 1735 345 1785
rect 255 1685 275 1735
rect 325 1685 345 1735
rect 255 1635 345 1685
rect 255 1585 275 1635
rect 325 1585 345 1635
rect 255 1535 345 1585
rect 255 1485 275 1535
rect 325 1485 345 1535
rect 255 1435 345 1485
rect 255 1385 275 1435
rect 325 1385 345 1435
rect 255 1335 345 1385
rect 255 1285 275 1335
rect 325 1285 345 1335
rect 255 1235 345 1285
rect 255 1185 275 1235
rect 325 1185 345 1235
rect 255 1135 345 1185
rect 255 1085 275 1135
rect 325 1085 345 1135
rect 255 1035 345 1085
rect 255 985 275 1035
rect 325 985 345 1035
rect 255 965 345 985
rect 445 2275 535 2295
rect 445 2225 465 2275
rect 515 2225 535 2275
rect 445 2135 535 2225
rect 445 2085 465 2135
rect 515 2085 535 2135
rect 445 2035 535 2085
rect 445 1985 465 2035
rect 515 1985 535 2035
rect 445 1935 535 1985
rect 445 1885 465 1935
rect 515 1885 535 1935
rect 445 1835 535 1885
rect 445 1785 465 1835
rect 515 1785 535 1835
rect 445 1735 535 1785
rect 445 1685 465 1735
rect 515 1685 535 1735
rect 445 1635 535 1685
rect 445 1585 465 1635
rect 515 1585 535 1635
rect 445 1535 535 1585
rect 445 1485 465 1535
rect 515 1485 535 1535
rect 445 1435 535 1485
rect 445 1385 465 1435
rect 515 1385 535 1435
rect 445 1335 535 1385
rect 445 1285 465 1335
rect 515 1285 535 1335
rect 445 1235 535 1285
rect 445 1185 465 1235
rect 515 1185 535 1235
rect 445 1135 535 1185
rect 445 1085 465 1135
rect 515 1085 535 1135
rect 445 1035 535 1085
rect 445 985 465 1035
rect 515 985 535 1035
rect 255 825 345 845
rect 255 775 275 825
rect 325 775 345 825
rect 255 755 345 775
rect 55 575 145 645
rect 55 525 75 575
rect 125 525 145 575
rect 55 475 145 525
rect 55 425 75 475
rect 125 425 145 475
rect 55 375 145 425
rect 55 325 75 375
rect 125 325 145 375
rect 55 275 145 325
rect 55 225 75 275
rect 125 225 145 275
rect 55 175 145 225
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 255 625 345 645
rect 255 575 275 625
rect 325 575 345 625
rect 255 475 345 575
rect 255 425 275 475
rect 325 425 345 475
rect 255 375 345 425
rect 255 325 275 375
rect 325 325 345 375
rect 255 275 345 325
rect 255 225 275 275
rect 325 225 345 275
rect 255 175 345 225
rect 255 125 275 175
rect 325 125 345 175
rect 255 45 345 125
rect 445 625 535 985
rect 445 575 465 625
rect 515 575 535 625
rect 445 475 535 575
rect 445 425 465 475
rect 515 425 535 475
rect 445 375 535 425
rect 445 325 465 375
rect 515 325 535 375
rect 445 275 535 325
rect 445 225 465 275
rect 515 225 535 275
rect 445 175 535 225
rect 445 125 465 175
rect 515 125 535 175
rect 445 105 535 125
rect 0 -45 590 45
<< labels >>
flabel metal1 s 75 -25 75 -25 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 65 2375 65 2375 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel nwell 215 855 215 855 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 475 725 475 725 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 275 -25 275 -25 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 265 2375 265 2375 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 275 765 275 765 2 FreeSans 400 0 0 0 a
port 2 ne
flabel nwell 565 855 565 855 2 FreeSans 400 0 0 0 vdd
<< end >>
