magic
tech scmos
magscale 1 2
timestamp 1570494029
<< error_p >>
rect 20 1320 22 1322
rect 18 1318 20 1320
rect 74 1290 76 1292
rect 104 1290 106 1292
rect 134 1290 136 1292
rect 164 1290 166 1292
rect 194 1290 196 1292
rect 224 1290 226 1292
rect 254 1290 256 1292
rect 284 1290 286 1292
rect 314 1290 316 1292
rect 344 1290 346 1292
rect 374 1290 376 1292
rect 404 1290 406 1292
rect 434 1290 436 1292
rect 464 1290 466 1292
rect 494 1290 496 1292
rect 524 1290 526 1292
rect 76 1288 78 1290
rect 82 1288 84 1290
rect 106 1288 108 1290
rect 112 1288 114 1290
rect 136 1288 138 1290
rect 142 1288 144 1290
rect 166 1288 168 1290
rect 172 1288 174 1290
rect 196 1288 198 1290
rect 202 1288 204 1290
rect 226 1288 228 1290
rect 232 1288 234 1290
rect 256 1288 258 1290
rect 262 1288 264 1290
rect 286 1288 288 1290
rect 292 1288 294 1290
rect 316 1288 318 1290
rect 322 1288 324 1290
rect 346 1288 348 1290
rect 352 1288 354 1290
rect 376 1288 378 1290
rect 382 1288 384 1290
rect 406 1288 408 1290
rect 412 1288 414 1290
rect 436 1288 438 1290
rect 442 1288 444 1290
rect 466 1288 468 1290
rect 472 1288 474 1290
rect 496 1288 498 1290
rect 502 1288 504 1290
rect 526 1288 528 1290
rect 532 1288 534 1290
rect 84 1286 86 1288
rect 114 1286 116 1288
rect 144 1286 146 1288
rect 174 1286 176 1288
rect 204 1286 206 1288
rect 234 1286 236 1288
rect 264 1286 266 1288
rect 294 1286 296 1288
rect 324 1286 326 1288
rect 354 1286 356 1288
rect 384 1286 386 1288
rect 414 1286 416 1288
rect 444 1286 446 1288
rect 474 1286 476 1288
rect 504 1286 506 1288
rect 534 1286 536 1288
rect 84 1280 86 1282
rect 114 1280 116 1282
rect 144 1280 146 1282
rect 174 1280 176 1282
rect 204 1280 206 1282
rect 234 1280 236 1282
rect 264 1280 266 1282
rect 294 1280 296 1282
rect 324 1280 326 1282
rect 354 1280 356 1282
rect 384 1280 386 1282
rect 414 1280 416 1282
rect 444 1280 446 1282
rect 474 1280 476 1282
rect 504 1280 506 1282
rect 534 1280 536 1282
rect 76 1278 78 1280
rect 82 1278 84 1280
rect 106 1278 108 1280
rect 112 1278 114 1280
rect 136 1278 138 1280
rect 142 1278 144 1280
rect 166 1278 168 1280
rect 172 1278 174 1280
rect 196 1278 198 1280
rect 202 1278 204 1280
rect 226 1278 228 1280
rect 232 1278 234 1280
rect 256 1278 258 1280
rect 262 1278 264 1280
rect 286 1278 288 1280
rect 292 1278 294 1280
rect 316 1278 318 1280
rect 322 1278 324 1280
rect 346 1278 348 1280
rect 352 1278 354 1280
rect 376 1278 378 1280
rect 382 1278 384 1280
rect 406 1278 408 1280
rect 412 1278 414 1280
rect 436 1278 438 1280
rect 442 1278 444 1280
rect 466 1278 468 1280
rect 472 1278 474 1280
rect 496 1278 498 1280
rect 502 1278 504 1280
rect 526 1278 528 1280
rect 532 1278 534 1280
rect 74 1276 76 1278
rect 104 1276 106 1278
rect 134 1276 136 1278
rect 164 1276 166 1278
rect 194 1276 196 1278
rect 224 1276 226 1278
rect 254 1276 256 1278
rect 284 1276 286 1278
rect 314 1276 316 1278
rect 344 1276 346 1278
rect 374 1276 376 1278
rect 404 1276 406 1278
rect 434 1276 436 1278
rect 464 1276 466 1278
rect 494 1276 496 1278
rect 524 1276 526 1278
rect 74 1270 76 1272
rect 104 1270 106 1272
rect 134 1270 136 1272
rect 164 1270 166 1272
rect 194 1270 196 1272
rect 224 1270 226 1272
rect 254 1270 256 1272
rect 284 1270 286 1272
rect 314 1270 316 1272
rect 344 1270 346 1272
rect 374 1270 376 1272
rect 404 1270 406 1272
rect 434 1270 436 1272
rect 464 1270 466 1272
rect 494 1270 496 1272
rect 524 1270 526 1272
rect 76 1268 78 1270
rect 82 1268 84 1270
rect 106 1268 108 1270
rect 112 1268 114 1270
rect 136 1268 138 1270
rect 142 1268 144 1270
rect 166 1268 168 1270
rect 172 1268 174 1270
rect 196 1268 198 1270
rect 202 1268 204 1270
rect 226 1268 228 1270
rect 232 1268 234 1270
rect 256 1268 258 1270
rect 262 1268 264 1270
rect 286 1268 288 1270
rect 292 1268 294 1270
rect 316 1268 318 1270
rect 322 1268 324 1270
rect 346 1268 348 1270
rect 352 1268 354 1270
rect 376 1268 378 1270
rect 382 1268 384 1270
rect 406 1268 408 1270
rect 412 1268 414 1270
rect 436 1268 438 1270
rect 442 1268 444 1270
rect 466 1268 468 1270
rect 472 1268 474 1270
rect 496 1268 498 1270
rect 502 1268 504 1270
rect 526 1268 528 1270
rect 532 1268 534 1270
rect 84 1266 86 1268
rect 114 1266 116 1268
rect 144 1266 146 1268
rect 174 1266 176 1268
rect 204 1266 206 1268
rect 234 1266 236 1268
rect 264 1266 266 1268
rect 294 1266 296 1268
rect 324 1266 326 1268
rect 354 1266 356 1268
rect 384 1266 386 1268
rect 414 1266 416 1268
rect 444 1266 446 1268
rect 474 1266 476 1268
rect 504 1266 506 1268
rect 534 1266 536 1268
rect 84 1260 86 1262
rect 114 1260 116 1262
rect 144 1260 146 1262
rect 174 1260 176 1262
rect 204 1260 206 1262
rect 234 1260 236 1262
rect 264 1260 266 1262
rect 294 1260 296 1262
rect 324 1260 326 1262
rect 354 1260 356 1262
rect 384 1260 386 1262
rect 414 1260 416 1262
rect 444 1260 446 1262
rect 474 1260 476 1262
rect 504 1260 506 1262
rect 534 1260 536 1262
rect 76 1258 78 1260
rect 82 1258 84 1260
rect 106 1258 108 1260
rect 112 1258 114 1260
rect 136 1258 138 1260
rect 142 1258 144 1260
rect 166 1258 168 1260
rect 172 1258 174 1260
rect 196 1258 198 1260
rect 202 1258 204 1260
rect 226 1258 228 1260
rect 232 1258 234 1260
rect 256 1258 258 1260
rect 262 1258 264 1260
rect 286 1258 288 1260
rect 292 1258 294 1260
rect 316 1258 318 1260
rect 322 1258 324 1260
rect 346 1258 348 1260
rect 352 1258 354 1260
rect 376 1258 378 1260
rect 382 1258 384 1260
rect 406 1258 408 1260
rect 412 1258 414 1260
rect 436 1258 438 1260
rect 442 1258 444 1260
rect 466 1258 468 1260
rect 472 1258 474 1260
rect 496 1258 498 1260
rect 502 1258 504 1260
rect 526 1258 528 1260
rect 532 1258 534 1260
rect 74 1256 76 1258
rect 104 1256 106 1258
rect 134 1256 136 1258
rect 164 1256 166 1258
rect 194 1256 196 1258
rect 224 1256 226 1258
rect 254 1256 256 1258
rect 284 1256 286 1258
rect 314 1256 316 1258
rect 344 1256 346 1258
rect 374 1256 376 1258
rect 404 1256 406 1258
rect 434 1256 436 1258
rect 464 1256 466 1258
rect 494 1256 496 1258
rect 524 1256 526 1258
rect 74 1250 76 1252
rect 104 1250 106 1252
rect 134 1250 136 1252
rect 164 1250 166 1252
rect 194 1250 196 1252
rect 224 1250 226 1252
rect 254 1250 256 1252
rect 284 1250 286 1252
rect 314 1250 316 1252
rect 344 1250 346 1252
rect 374 1250 376 1252
rect 404 1250 406 1252
rect 434 1250 436 1252
rect 464 1250 466 1252
rect 494 1250 496 1252
rect 524 1250 526 1252
rect 76 1248 78 1250
rect 82 1248 84 1250
rect 106 1248 108 1250
rect 112 1248 114 1250
rect 136 1248 138 1250
rect 142 1248 144 1250
rect 166 1248 168 1250
rect 172 1248 174 1250
rect 196 1248 198 1250
rect 202 1248 204 1250
rect 226 1248 228 1250
rect 232 1248 234 1250
rect 256 1248 258 1250
rect 262 1248 264 1250
rect 286 1248 288 1250
rect 292 1248 294 1250
rect 316 1248 318 1250
rect 322 1248 324 1250
rect 346 1248 348 1250
rect 352 1248 354 1250
rect 376 1248 378 1250
rect 382 1248 384 1250
rect 406 1248 408 1250
rect 412 1248 414 1250
rect 436 1248 438 1250
rect 442 1248 444 1250
rect 466 1248 468 1250
rect 472 1248 474 1250
rect 496 1248 498 1250
rect 502 1248 504 1250
rect 526 1248 528 1250
rect 532 1248 534 1250
rect 84 1246 86 1248
rect 114 1246 116 1248
rect 144 1246 146 1248
rect 174 1246 176 1248
rect 204 1246 206 1248
rect 234 1246 236 1248
rect 264 1246 266 1248
rect 294 1246 296 1248
rect 324 1246 326 1248
rect 354 1246 356 1248
rect 384 1246 386 1248
rect 414 1246 416 1248
rect 444 1246 446 1248
rect 474 1246 476 1248
rect 504 1246 506 1248
rect 534 1246 536 1248
rect 84 1240 86 1242
rect 114 1240 116 1242
rect 144 1240 146 1242
rect 174 1240 176 1242
rect 204 1240 206 1242
rect 234 1240 236 1242
rect 264 1240 266 1242
rect 294 1240 296 1242
rect 324 1240 326 1242
rect 354 1240 356 1242
rect 384 1240 386 1242
rect 414 1240 416 1242
rect 444 1240 446 1242
rect 474 1240 476 1242
rect 504 1240 506 1242
rect 534 1240 536 1242
rect 76 1238 78 1240
rect 82 1238 84 1240
rect 106 1238 108 1240
rect 112 1238 114 1240
rect 136 1238 138 1240
rect 142 1238 144 1240
rect 166 1238 168 1240
rect 172 1238 174 1240
rect 196 1238 198 1240
rect 202 1238 204 1240
rect 226 1238 228 1240
rect 232 1238 234 1240
rect 256 1238 258 1240
rect 262 1238 264 1240
rect 286 1238 288 1240
rect 292 1238 294 1240
rect 316 1238 318 1240
rect 322 1238 324 1240
rect 346 1238 348 1240
rect 352 1238 354 1240
rect 376 1238 378 1240
rect 382 1238 384 1240
rect 406 1238 408 1240
rect 412 1238 414 1240
rect 436 1238 438 1240
rect 442 1238 444 1240
rect 466 1238 468 1240
rect 472 1238 474 1240
rect 496 1238 498 1240
rect 502 1238 504 1240
rect 526 1238 528 1240
rect 532 1238 534 1240
rect 74 1236 76 1238
rect 104 1236 106 1238
rect 134 1236 136 1238
rect 164 1236 166 1238
rect 194 1236 196 1238
rect 224 1236 226 1238
rect 254 1236 256 1238
rect 284 1236 286 1238
rect 314 1236 316 1238
rect 344 1236 346 1238
rect 374 1236 376 1238
rect 404 1236 406 1238
rect 434 1236 436 1238
rect 464 1236 466 1238
rect 494 1236 496 1238
rect 524 1236 526 1238
rect 74 1230 76 1232
rect 104 1230 106 1232
rect 134 1230 136 1232
rect 164 1230 166 1232
rect 194 1230 196 1232
rect 224 1230 226 1232
rect 254 1230 256 1232
rect 284 1230 286 1232
rect 314 1230 316 1232
rect 344 1230 346 1232
rect 374 1230 376 1232
rect 404 1230 406 1232
rect 434 1230 436 1232
rect 464 1230 466 1232
rect 494 1230 496 1232
rect 524 1230 526 1232
rect 76 1228 78 1230
rect 82 1228 84 1230
rect 106 1228 108 1230
rect 112 1228 114 1230
rect 136 1228 138 1230
rect 142 1228 144 1230
rect 166 1228 168 1230
rect 172 1228 174 1230
rect 196 1228 198 1230
rect 202 1228 204 1230
rect 226 1228 228 1230
rect 232 1228 234 1230
rect 256 1228 258 1230
rect 262 1228 264 1230
rect 286 1228 288 1230
rect 292 1228 294 1230
rect 316 1228 318 1230
rect 322 1228 324 1230
rect 346 1228 348 1230
rect 352 1228 354 1230
rect 376 1228 378 1230
rect 382 1228 384 1230
rect 406 1228 408 1230
rect 412 1228 414 1230
rect 436 1228 438 1230
rect 442 1228 444 1230
rect 466 1228 468 1230
rect 472 1228 474 1230
rect 496 1228 498 1230
rect 502 1228 504 1230
rect 526 1228 528 1230
rect 532 1228 534 1230
rect 84 1226 86 1228
rect 114 1226 116 1228
rect 144 1226 146 1228
rect 174 1226 176 1228
rect 204 1226 206 1228
rect 234 1226 236 1228
rect 264 1226 266 1228
rect 294 1226 296 1228
rect 324 1226 326 1228
rect 354 1226 356 1228
rect 384 1226 386 1228
rect 414 1226 416 1228
rect 444 1226 446 1228
rect 474 1226 476 1228
rect 504 1226 506 1228
rect 534 1226 536 1228
rect 84 1220 86 1222
rect 114 1220 116 1222
rect 144 1220 146 1222
rect 174 1220 176 1222
rect 204 1220 206 1222
rect 234 1220 236 1222
rect 264 1220 266 1222
rect 294 1220 296 1222
rect 324 1220 326 1222
rect 354 1220 356 1222
rect 384 1220 386 1222
rect 414 1220 416 1222
rect 444 1220 446 1222
rect 474 1220 476 1222
rect 504 1220 506 1222
rect 534 1220 536 1222
rect 76 1218 78 1220
rect 82 1218 84 1220
rect 106 1218 108 1220
rect 112 1218 114 1220
rect 136 1218 138 1220
rect 142 1218 144 1220
rect 166 1218 168 1220
rect 172 1218 174 1220
rect 196 1218 198 1220
rect 202 1218 204 1220
rect 226 1218 228 1220
rect 232 1218 234 1220
rect 256 1218 258 1220
rect 262 1218 264 1220
rect 286 1218 288 1220
rect 292 1218 294 1220
rect 316 1218 318 1220
rect 322 1218 324 1220
rect 346 1218 348 1220
rect 352 1218 354 1220
rect 376 1218 378 1220
rect 382 1218 384 1220
rect 406 1218 408 1220
rect 412 1218 414 1220
rect 436 1218 438 1220
rect 442 1218 444 1220
rect 466 1218 468 1220
rect 472 1218 474 1220
rect 496 1218 498 1220
rect 502 1218 504 1220
rect 526 1218 528 1220
rect 532 1218 534 1220
rect 74 1216 76 1218
rect 104 1216 106 1218
rect 134 1216 136 1218
rect 164 1216 166 1218
rect 194 1216 196 1218
rect 224 1216 226 1218
rect 254 1216 256 1218
rect 284 1216 286 1218
rect 314 1216 316 1218
rect 344 1216 346 1218
rect 374 1216 376 1218
rect 404 1216 406 1218
rect 434 1216 436 1218
rect 464 1216 466 1218
rect 494 1216 496 1218
rect 524 1216 526 1218
rect 74 1210 76 1212
rect 104 1210 106 1212
rect 134 1210 136 1212
rect 164 1210 166 1212
rect 194 1210 196 1212
rect 224 1210 226 1212
rect 254 1210 256 1212
rect 284 1210 286 1212
rect 314 1210 316 1212
rect 344 1210 346 1212
rect 374 1210 376 1212
rect 404 1210 406 1212
rect 434 1210 436 1212
rect 464 1210 466 1212
rect 494 1210 496 1212
rect 524 1210 526 1212
rect 76 1208 78 1210
rect 82 1208 84 1210
rect 106 1208 108 1210
rect 112 1208 114 1210
rect 136 1208 138 1210
rect 142 1208 144 1210
rect 166 1208 168 1210
rect 172 1208 174 1210
rect 196 1208 198 1210
rect 202 1208 204 1210
rect 226 1208 228 1210
rect 232 1208 234 1210
rect 256 1208 258 1210
rect 262 1208 264 1210
rect 286 1208 288 1210
rect 292 1208 294 1210
rect 316 1208 318 1210
rect 322 1208 324 1210
rect 346 1208 348 1210
rect 352 1208 354 1210
rect 376 1208 378 1210
rect 382 1208 384 1210
rect 406 1208 408 1210
rect 412 1208 414 1210
rect 436 1208 438 1210
rect 442 1208 444 1210
rect 466 1208 468 1210
rect 472 1208 474 1210
rect 496 1208 498 1210
rect 502 1208 504 1210
rect 526 1208 528 1210
rect 532 1208 534 1210
rect 84 1206 86 1208
rect 114 1206 116 1208
rect 144 1206 146 1208
rect 174 1206 176 1208
rect 204 1206 206 1208
rect 234 1206 236 1208
rect 264 1206 266 1208
rect 294 1206 296 1208
rect 324 1206 326 1208
rect 354 1206 356 1208
rect 384 1206 386 1208
rect 414 1206 416 1208
rect 444 1206 446 1208
rect 474 1206 476 1208
rect 504 1206 506 1208
rect 534 1206 536 1208
rect 84 1200 86 1202
rect 114 1200 116 1202
rect 144 1200 146 1202
rect 174 1200 176 1202
rect 204 1200 206 1202
rect 234 1200 236 1202
rect 264 1200 266 1202
rect 294 1200 296 1202
rect 324 1200 326 1202
rect 354 1200 356 1202
rect 384 1200 386 1202
rect 414 1200 416 1202
rect 444 1200 446 1202
rect 474 1200 476 1202
rect 504 1200 506 1202
rect 534 1200 536 1202
rect 76 1198 78 1200
rect 82 1198 84 1200
rect 106 1198 108 1200
rect 112 1198 114 1200
rect 136 1198 138 1200
rect 142 1198 144 1200
rect 166 1198 168 1200
rect 172 1198 174 1200
rect 196 1198 198 1200
rect 202 1198 204 1200
rect 226 1198 228 1200
rect 232 1198 234 1200
rect 256 1198 258 1200
rect 262 1198 264 1200
rect 286 1198 288 1200
rect 292 1198 294 1200
rect 316 1198 318 1200
rect 322 1198 324 1200
rect 346 1198 348 1200
rect 352 1198 354 1200
rect 376 1198 378 1200
rect 382 1198 384 1200
rect 406 1198 408 1200
rect 412 1198 414 1200
rect 436 1198 438 1200
rect 442 1198 444 1200
rect 466 1198 468 1200
rect 472 1198 474 1200
rect 496 1198 498 1200
rect 502 1198 504 1200
rect 526 1198 528 1200
rect 532 1198 534 1200
rect 74 1196 76 1198
rect 104 1196 106 1198
rect 134 1196 136 1198
rect 164 1196 166 1198
rect 194 1196 196 1198
rect 224 1196 226 1198
rect 254 1196 256 1198
rect 284 1196 286 1198
rect 314 1196 316 1198
rect 344 1196 346 1198
rect 374 1196 376 1198
rect 404 1196 406 1198
rect 434 1196 436 1198
rect 464 1196 466 1198
rect 494 1196 496 1198
rect 524 1196 526 1198
rect 74 1190 76 1192
rect 524 1190 526 1192
rect 76 1188 78 1190
rect 82 1188 84 1190
rect 526 1188 528 1190
rect 532 1188 534 1190
rect 84 1186 86 1188
rect 534 1186 536 1188
rect 84 1180 86 1182
rect 534 1180 536 1182
rect 76 1178 78 1180
rect 82 1178 84 1180
rect 526 1178 528 1180
rect 532 1178 534 1180
rect 74 1176 76 1178
rect 524 1176 526 1178
rect 74 1170 76 1172
rect 104 1170 106 1172
rect 134 1170 136 1172
rect 164 1170 166 1172
rect 194 1170 196 1172
rect 224 1170 226 1172
rect 254 1170 256 1172
rect 284 1170 286 1172
rect 314 1170 316 1172
rect 344 1170 346 1172
rect 374 1170 376 1172
rect 404 1170 406 1172
rect 434 1170 436 1172
rect 464 1170 466 1172
rect 494 1170 496 1172
rect 524 1170 526 1172
rect 76 1168 78 1170
rect 82 1168 84 1170
rect 106 1168 108 1170
rect 112 1168 114 1170
rect 136 1168 138 1170
rect 142 1168 144 1170
rect 166 1168 168 1170
rect 172 1168 174 1170
rect 196 1168 198 1170
rect 202 1168 204 1170
rect 226 1168 228 1170
rect 232 1168 234 1170
rect 256 1168 258 1170
rect 262 1168 264 1170
rect 286 1168 288 1170
rect 292 1168 294 1170
rect 316 1168 318 1170
rect 322 1168 324 1170
rect 346 1168 348 1170
rect 352 1168 354 1170
rect 376 1168 378 1170
rect 382 1168 384 1170
rect 406 1168 408 1170
rect 412 1168 414 1170
rect 436 1168 438 1170
rect 442 1168 444 1170
rect 466 1168 468 1170
rect 472 1168 474 1170
rect 496 1168 498 1170
rect 502 1168 504 1170
rect 526 1168 528 1170
rect 532 1168 534 1170
rect 84 1166 86 1168
rect 114 1166 116 1168
rect 144 1166 146 1168
rect 174 1166 176 1168
rect 204 1166 206 1168
rect 234 1166 236 1168
rect 264 1166 266 1168
rect 294 1166 296 1168
rect 324 1166 326 1168
rect 354 1166 356 1168
rect 384 1166 386 1168
rect 414 1166 416 1168
rect 444 1166 446 1168
rect 474 1166 476 1168
rect 504 1166 506 1168
rect 534 1166 536 1168
rect 84 1160 86 1162
rect 114 1160 116 1162
rect 144 1160 146 1162
rect 174 1160 176 1162
rect 204 1160 206 1162
rect 234 1160 236 1162
rect 264 1160 266 1162
rect 294 1160 296 1162
rect 324 1160 326 1162
rect 354 1160 356 1162
rect 384 1160 386 1162
rect 414 1160 416 1162
rect 444 1160 446 1162
rect 474 1160 476 1162
rect 504 1160 506 1162
rect 534 1160 536 1162
rect 76 1158 78 1160
rect 82 1158 84 1160
rect 106 1158 108 1160
rect 112 1158 114 1160
rect 136 1158 138 1160
rect 142 1158 144 1160
rect 166 1158 168 1160
rect 172 1158 174 1160
rect 196 1158 198 1160
rect 202 1158 204 1160
rect 226 1158 228 1160
rect 232 1158 234 1160
rect 256 1158 258 1160
rect 262 1158 264 1160
rect 286 1158 288 1160
rect 292 1158 294 1160
rect 316 1158 318 1160
rect 322 1158 324 1160
rect 346 1158 348 1160
rect 352 1158 354 1160
rect 376 1158 378 1160
rect 382 1158 384 1160
rect 406 1158 408 1160
rect 412 1158 414 1160
rect 436 1158 438 1160
rect 442 1158 444 1160
rect 466 1158 468 1160
rect 472 1158 474 1160
rect 496 1158 498 1160
rect 502 1158 504 1160
rect 526 1158 528 1160
rect 532 1158 534 1160
rect 74 1156 76 1158
rect 104 1156 106 1158
rect 134 1156 136 1158
rect 164 1156 166 1158
rect 194 1156 196 1158
rect 224 1156 226 1158
rect 254 1156 256 1158
rect 284 1156 286 1158
rect 314 1156 316 1158
rect 344 1156 346 1158
rect 374 1156 376 1158
rect 404 1156 406 1158
rect 434 1156 436 1158
rect 464 1156 466 1158
rect 494 1156 496 1158
rect 524 1156 526 1158
rect 74 1150 76 1152
rect 104 1150 106 1152
rect 134 1150 136 1152
rect 164 1150 166 1152
rect 194 1150 196 1152
rect 224 1150 226 1152
rect 254 1150 256 1152
rect 284 1150 286 1152
rect 314 1150 316 1152
rect 344 1150 346 1152
rect 374 1150 376 1152
rect 404 1150 406 1152
rect 434 1150 436 1152
rect 464 1150 466 1152
rect 494 1150 496 1152
rect 524 1150 526 1152
rect 76 1148 78 1150
rect 82 1148 84 1150
rect 106 1148 108 1150
rect 112 1148 114 1150
rect 136 1148 138 1150
rect 142 1148 144 1150
rect 166 1148 168 1150
rect 172 1148 174 1150
rect 196 1148 198 1150
rect 202 1148 204 1150
rect 226 1148 228 1150
rect 232 1148 234 1150
rect 256 1148 258 1150
rect 262 1148 264 1150
rect 286 1148 288 1150
rect 292 1148 294 1150
rect 316 1148 318 1150
rect 322 1148 324 1150
rect 346 1148 348 1150
rect 352 1148 354 1150
rect 376 1148 378 1150
rect 382 1148 384 1150
rect 406 1148 408 1150
rect 412 1148 414 1150
rect 436 1148 438 1150
rect 442 1148 444 1150
rect 466 1148 468 1150
rect 472 1148 474 1150
rect 496 1148 498 1150
rect 502 1148 504 1150
rect 526 1148 528 1150
rect 532 1148 534 1150
rect 84 1146 86 1148
rect 114 1146 116 1148
rect 144 1146 146 1148
rect 174 1146 176 1148
rect 204 1146 206 1148
rect 234 1146 236 1148
rect 264 1146 266 1148
rect 294 1146 296 1148
rect 324 1146 326 1148
rect 354 1146 356 1148
rect 384 1146 386 1148
rect 414 1146 416 1148
rect 444 1146 446 1148
rect 474 1146 476 1148
rect 504 1146 506 1148
rect 534 1146 536 1148
rect 84 1140 86 1142
rect 114 1140 116 1142
rect 144 1140 146 1142
rect 174 1140 176 1142
rect 204 1140 206 1142
rect 234 1140 236 1142
rect 264 1140 266 1142
rect 294 1140 296 1142
rect 324 1140 326 1142
rect 354 1140 356 1142
rect 384 1140 386 1142
rect 414 1140 416 1142
rect 444 1140 446 1142
rect 474 1140 476 1142
rect 504 1140 506 1142
rect 534 1140 536 1142
rect 76 1138 78 1140
rect 82 1138 84 1140
rect 106 1138 108 1140
rect 112 1138 114 1140
rect 136 1138 138 1140
rect 142 1138 144 1140
rect 166 1138 168 1140
rect 172 1138 174 1140
rect 196 1138 198 1140
rect 202 1138 204 1140
rect 226 1138 228 1140
rect 232 1138 234 1140
rect 256 1138 258 1140
rect 262 1138 264 1140
rect 286 1138 288 1140
rect 292 1138 294 1140
rect 316 1138 318 1140
rect 322 1138 324 1140
rect 346 1138 348 1140
rect 352 1138 354 1140
rect 376 1138 378 1140
rect 382 1138 384 1140
rect 406 1138 408 1140
rect 412 1138 414 1140
rect 436 1138 438 1140
rect 442 1138 444 1140
rect 466 1138 468 1140
rect 472 1138 474 1140
rect 496 1138 498 1140
rect 502 1138 504 1140
rect 526 1138 528 1140
rect 532 1138 534 1140
rect 74 1136 76 1138
rect 104 1136 106 1138
rect 134 1136 136 1138
rect 164 1136 166 1138
rect 194 1136 196 1138
rect 224 1136 226 1138
rect 254 1136 256 1138
rect 284 1136 286 1138
rect 314 1136 316 1138
rect 344 1136 346 1138
rect 374 1136 376 1138
rect 404 1136 406 1138
rect 434 1136 436 1138
rect 464 1136 466 1138
rect 494 1136 496 1138
rect 524 1136 526 1138
rect 74 1130 76 1132
rect 104 1130 106 1132
rect 134 1130 136 1132
rect 164 1130 166 1132
rect 194 1130 196 1132
rect 224 1130 226 1132
rect 254 1130 256 1132
rect 284 1130 286 1132
rect 314 1130 316 1132
rect 344 1130 346 1132
rect 374 1130 376 1132
rect 404 1130 406 1132
rect 434 1130 436 1132
rect 464 1130 466 1132
rect 494 1130 496 1132
rect 524 1130 526 1132
rect 76 1128 78 1130
rect 82 1128 84 1130
rect 106 1128 108 1130
rect 112 1128 114 1130
rect 136 1128 138 1130
rect 142 1128 144 1130
rect 166 1128 168 1130
rect 172 1128 174 1130
rect 196 1128 198 1130
rect 202 1128 204 1130
rect 226 1128 228 1130
rect 232 1128 234 1130
rect 256 1128 258 1130
rect 262 1128 264 1130
rect 286 1128 288 1130
rect 292 1128 294 1130
rect 316 1128 318 1130
rect 322 1128 324 1130
rect 346 1128 348 1130
rect 352 1128 354 1130
rect 376 1128 378 1130
rect 382 1128 384 1130
rect 406 1128 408 1130
rect 412 1128 414 1130
rect 436 1128 438 1130
rect 442 1128 444 1130
rect 466 1128 468 1130
rect 472 1128 474 1130
rect 496 1128 498 1130
rect 502 1128 504 1130
rect 526 1128 528 1130
rect 532 1128 534 1130
rect 84 1126 86 1128
rect 114 1126 116 1128
rect 144 1126 146 1128
rect 174 1126 176 1128
rect 204 1126 206 1128
rect 234 1126 236 1128
rect 264 1126 266 1128
rect 294 1126 296 1128
rect 324 1126 326 1128
rect 354 1126 356 1128
rect 384 1126 386 1128
rect 414 1126 416 1128
rect 444 1126 446 1128
rect 474 1126 476 1128
rect 504 1126 506 1128
rect 534 1126 536 1128
rect 84 1120 86 1122
rect 504 1120 506 1122
rect 534 1120 536 1122
rect 86 1118 88 1120
rect 506 1118 508 1120
rect 532 1118 534 1120
rect 86 1108 88 1110
rect 506 1108 508 1110
rect 532 1108 534 1110
rect 84 1106 86 1108
rect 504 1106 506 1108
rect 534 1106 536 1108
rect 84 1100 86 1102
rect 114 1100 116 1102
rect 144 1100 146 1102
rect 174 1100 176 1102
rect 204 1100 206 1102
rect 234 1100 236 1102
rect 264 1100 266 1102
rect 294 1100 296 1102
rect 324 1100 326 1102
rect 354 1100 356 1102
rect 384 1100 386 1102
rect 414 1100 416 1102
rect 444 1100 446 1102
rect 474 1100 476 1102
rect 504 1100 506 1102
rect 534 1100 536 1102
rect 76 1098 78 1100
rect 82 1098 84 1100
rect 106 1098 108 1100
rect 112 1098 114 1100
rect 136 1098 138 1100
rect 142 1098 144 1100
rect 166 1098 168 1100
rect 172 1098 174 1100
rect 196 1098 198 1100
rect 202 1098 204 1100
rect 226 1098 228 1100
rect 232 1098 234 1100
rect 256 1098 258 1100
rect 262 1098 264 1100
rect 286 1098 288 1100
rect 292 1098 294 1100
rect 316 1098 318 1100
rect 322 1098 324 1100
rect 346 1098 348 1100
rect 352 1098 354 1100
rect 376 1098 378 1100
rect 382 1098 384 1100
rect 406 1098 408 1100
rect 412 1098 414 1100
rect 436 1098 438 1100
rect 442 1098 444 1100
rect 466 1098 468 1100
rect 472 1098 474 1100
rect 496 1098 498 1100
rect 502 1098 504 1100
rect 526 1098 528 1100
rect 532 1098 534 1100
rect 74 1096 76 1098
rect 104 1096 106 1098
rect 134 1096 136 1098
rect 164 1096 166 1098
rect 194 1096 196 1098
rect 224 1096 226 1098
rect 254 1096 256 1098
rect 284 1096 286 1098
rect 314 1096 316 1098
rect 344 1096 346 1098
rect 374 1096 376 1098
rect 404 1096 406 1098
rect 434 1096 436 1098
rect 464 1096 466 1098
rect 494 1096 496 1098
rect 524 1096 526 1098
rect 74 1090 76 1092
rect 104 1090 106 1092
rect 134 1090 136 1092
rect 164 1090 166 1092
rect 194 1090 196 1092
rect 224 1090 226 1092
rect 254 1090 256 1092
rect 284 1090 286 1092
rect 314 1090 316 1092
rect 344 1090 346 1092
rect 374 1090 376 1092
rect 404 1090 406 1092
rect 434 1090 436 1092
rect 464 1090 466 1092
rect 494 1090 496 1092
rect 524 1090 526 1092
rect 76 1088 78 1090
rect 82 1088 84 1090
rect 106 1088 108 1090
rect 112 1088 114 1090
rect 136 1088 138 1090
rect 142 1088 144 1090
rect 166 1088 168 1090
rect 172 1088 174 1090
rect 196 1088 198 1090
rect 202 1088 204 1090
rect 226 1088 228 1090
rect 232 1088 234 1090
rect 256 1088 258 1090
rect 262 1088 264 1090
rect 286 1088 288 1090
rect 292 1088 294 1090
rect 316 1088 318 1090
rect 322 1088 324 1090
rect 346 1088 348 1090
rect 352 1088 354 1090
rect 376 1088 378 1090
rect 382 1088 384 1090
rect 406 1088 408 1090
rect 412 1088 414 1090
rect 436 1088 438 1090
rect 442 1088 444 1090
rect 466 1088 468 1090
rect 472 1088 474 1090
rect 496 1088 498 1090
rect 502 1088 504 1090
rect 526 1088 528 1090
rect 532 1088 534 1090
rect 84 1086 86 1088
rect 114 1086 116 1088
rect 144 1086 146 1088
rect 174 1086 176 1088
rect 204 1086 206 1088
rect 234 1086 236 1088
rect 264 1086 266 1088
rect 294 1086 296 1088
rect 324 1086 326 1088
rect 354 1086 356 1088
rect 384 1086 386 1088
rect 414 1086 416 1088
rect 444 1086 446 1088
rect 474 1086 476 1088
rect 504 1086 506 1088
rect 534 1086 536 1088
rect 84 1080 86 1082
rect 114 1080 116 1082
rect 144 1080 146 1082
rect 174 1080 176 1082
rect 204 1080 206 1082
rect 234 1080 236 1082
rect 264 1080 266 1082
rect 294 1080 296 1082
rect 324 1080 326 1082
rect 354 1080 356 1082
rect 384 1080 386 1082
rect 414 1080 416 1082
rect 444 1080 446 1082
rect 474 1080 476 1082
rect 504 1080 506 1082
rect 534 1080 536 1082
rect 76 1078 78 1080
rect 82 1078 84 1080
rect 106 1078 108 1080
rect 112 1078 114 1080
rect 136 1078 138 1080
rect 142 1078 144 1080
rect 166 1078 168 1080
rect 172 1078 174 1080
rect 196 1078 198 1080
rect 202 1078 204 1080
rect 226 1078 228 1080
rect 232 1078 234 1080
rect 256 1078 258 1080
rect 262 1078 264 1080
rect 286 1078 288 1080
rect 292 1078 294 1080
rect 316 1078 318 1080
rect 322 1078 324 1080
rect 346 1078 348 1080
rect 352 1078 354 1080
rect 376 1078 378 1080
rect 382 1078 384 1080
rect 406 1078 408 1080
rect 412 1078 414 1080
rect 436 1078 438 1080
rect 442 1078 444 1080
rect 466 1078 468 1080
rect 472 1078 474 1080
rect 496 1078 498 1080
rect 502 1078 504 1080
rect 526 1078 528 1080
rect 532 1078 534 1080
rect 74 1076 76 1078
rect 104 1076 106 1078
rect 134 1076 136 1078
rect 164 1076 166 1078
rect 194 1076 196 1078
rect 224 1076 226 1078
rect 254 1076 256 1078
rect 284 1076 286 1078
rect 314 1076 316 1078
rect 344 1076 346 1078
rect 374 1076 376 1078
rect 404 1076 406 1078
rect 434 1076 436 1078
rect 464 1076 466 1078
rect 494 1076 496 1078
rect 524 1076 526 1078
rect 74 1070 76 1072
rect 104 1070 106 1072
rect 134 1070 136 1072
rect 164 1070 166 1072
rect 194 1070 196 1072
rect 224 1070 226 1072
rect 254 1070 256 1072
rect 284 1070 286 1072
rect 314 1070 316 1072
rect 344 1070 346 1072
rect 374 1070 376 1072
rect 404 1070 406 1072
rect 434 1070 436 1072
rect 464 1070 466 1072
rect 494 1070 496 1072
rect 524 1070 526 1072
rect 76 1068 78 1070
rect 82 1068 84 1070
rect 106 1068 108 1070
rect 112 1068 114 1070
rect 136 1068 138 1070
rect 142 1068 144 1070
rect 166 1068 168 1070
rect 172 1068 174 1070
rect 196 1068 198 1070
rect 202 1068 204 1070
rect 226 1068 228 1070
rect 232 1068 234 1070
rect 256 1068 258 1070
rect 262 1068 264 1070
rect 286 1068 288 1070
rect 292 1068 294 1070
rect 316 1068 318 1070
rect 322 1068 324 1070
rect 346 1068 348 1070
rect 352 1068 354 1070
rect 376 1068 378 1070
rect 382 1068 384 1070
rect 406 1068 408 1070
rect 412 1068 414 1070
rect 436 1068 438 1070
rect 442 1068 444 1070
rect 466 1068 468 1070
rect 472 1068 474 1070
rect 496 1068 498 1070
rect 502 1068 504 1070
rect 526 1068 528 1070
rect 532 1068 534 1070
rect 84 1066 86 1068
rect 114 1066 116 1068
rect 144 1066 146 1068
rect 174 1066 176 1068
rect 204 1066 206 1068
rect 234 1066 236 1068
rect 264 1066 266 1068
rect 294 1066 296 1068
rect 324 1066 326 1068
rect 354 1066 356 1068
rect 384 1066 386 1068
rect 414 1066 416 1068
rect 444 1066 446 1068
rect 474 1066 476 1068
rect 504 1066 506 1068
rect 534 1066 536 1068
rect 84 1060 86 1062
rect 114 1060 116 1062
rect 144 1060 146 1062
rect 174 1060 176 1062
rect 204 1060 206 1062
rect 234 1060 236 1062
rect 264 1060 266 1062
rect 294 1060 296 1062
rect 324 1060 326 1062
rect 354 1060 356 1062
rect 384 1060 386 1062
rect 414 1060 416 1062
rect 444 1060 446 1062
rect 474 1060 476 1062
rect 504 1060 506 1062
rect 534 1060 536 1062
rect 76 1058 78 1060
rect 82 1058 84 1060
rect 106 1058 108 1060
rect 112 1058 114 1060
rect 136 1058 138 1060
rect 142 1058 144 1060
rect 166 1058 168 1060
rect 172 1058 174 1060
rect 196 1058 198 1060
rect 202 1058 204 1060
rect 226 1058 228 1060
rect 232 1058 234 1060
rect 256 1058 258 1060
rect 262 1058 264 1060
rect 286 1058 288 1060
rect 292 1058 294 1060
rect 316 1058 318 1060
rect 322 1058 324 1060
rect 346 1058 348 1060
rect 352 1058 354 1060
rect 376 1058 378 1060
rect 382 1058 384 1060
rect 406 1058 408 1060
rect 412 1058 414 1060
rect 436 1058 438 1060
rect 442 1058 444 1060
rect 466 1058 468 1060
rect 472 1058 474 1060
rect 496 1058 498 1060
rect 502 1058 504 1060
rect 526 1058 528 1060
rect 532 1058 534 1060
rect 74 1056 76 1058
rect 104 1056 106 1058
rect 134 1056 136 1058
rect 164 1056 166 1058
rect 194 1056 196 1058
rect 224 1056 226 1058
rect 254 1056 256 1058
rect 284 1056 286 1058
rect 314 1056 316 1058
rect 344 1056 346 1058
rect 374 1056 376 1058
rect 404 1056 406 1058
rect 434 1056 436 1058
rect 464 1056 466 1058
rect 494 1056 496 1058
rect 524 1056 526 1058
rect 74 1050 76 1052
rect 104 1050 106 1052
rect 134 1050 136 1052
rect 164 1050 166 1052
rect 194 1050 196 1052
rect 224 1050 226 1052
rect 254 1050 256 1052
rect 284 1050 286 1052
rect 314 1050 316 1052
rect 344 1050 346 1052
rect 374 1050 376 1052
rect 404 1050 406 1052
rect 434 1050 436 1052
rect 464 1050 466 1052
rect 494 1050 496 1052
rect 524 1050 526 1052
rect 76 1048 78 1050
rect 82 1048 84 1050
rect 106 1048 108 1050
rect 112 1048 114 1050
rect 136 1048 138 1050
rect 142 1048 144 1050
rect 166 1048 168 1050
rect 172 1048 174 1050
rect 196 1048 198 1050
rect 202 1048 204 1050
rect 226 1048 228 1050
rect 232 1048 234 1050
rect 256 1048 258 1050
rect 262 1048 264 1050
rect 286 1048 288 1050
rect 292 1048 294 1050
rect 316 1048 318 1050
rect 322 1048 324 1050
rect 346 1048 348 1050
rect 352 1048 354 1050
rect 376 1048 378 1050
rect 382 1048 384 1050
rect 406 1048 408 1050
rect 412 1048 414 1050
rect 436 1048 438 1050
rect 442 1048 444 1050
rect 466 1048 468 1050
rect 472 1048 474 1050
rect 496 1048 498 1050
rect 502 1048 504 1050
rect 526 1048 528 1050
rect 532 1048 534 1050
rect 84 1046 86 1048
rect 114 1046 116 1048
rect 144 1046 146 1048
rect 174 1046 176 1048
rect 204 1046 206 1048
rect 234 1046 236 1048
rect 264 1046 266 1048
rect 294 1046 296 1048
rect 324 1046 326 1048
rect 354 1046 356 1048
rect 384 1046 386 1048
rect 414 1046 416 1048
rect 444 1046 446 1048
rect 474 1046 476 1048
rect 504 1046 506 1048
rect 534 1046 536 1048
rect 84 1040 86 1042
rect 504 1040 506 1042
rect 534 1040 536 1042
rect 76 1038 78 1040
rect 82 1038 84 1040
rect 506 1038 508 1040
rect 532 1038 534 1040
rect 74 1036 76 1038
rect 74 1030 76 1032
rect 76 1028 78 1030
rect 82 1028 84 1030
rect 506 1028 508 1030
rect 532 1028 534 1030
rect 84 1026 86 1028
rect 504 1026 506 1028
rect 534 1026 536 1028
rect 84 1020 86 1022
rect 114 1020 116 1022
rect 144 1020 146 1022
rect 174 1020 176 1022
rect 204 1020 206 1022
rect 234 1020 236 1022
rect 264 1020 266 1022
rect 294 1020 296 1022
rect 324 1020 326 1022
rect 354 1020 356 1022
rect 384 1020 386 1022
rect 414 1020 416 1022
rect 444 1020 446 1022
rect 474 1020 476 1022
rect 504 1020 506 1022
rect 534 1020 536 1022
rect 76 1018 78 1020
rect 82 1018 84 1020
rect 106 1018 108 1020
rect 112 1018 114 1020
rect 136 1018 138 1020
rect 142 1018 144 1020
rect 166 1018 168 1020
rect 172 1018 174 1020
rect 196 1018 198 1020
rect 202 1018 204 1020
rect 226 1018 228 1020
rect 232 1018 234 1020
rect 256 1018 258 1020
rect 262 1018 264 1020
rect 286 1018 288 1020
rect 292 1018 294 1020
rect 316 1018 318 1020
rect 322 1018 324 1020
rect 346 1018 348 1020
rect 352 1018 354 1020
rect 376 1018 378 1020
rect 382 1018 384 1020
rect 406 1018 408 1020
rect 412 1018 414 1020
rect 436 1018 438 1020
rect 442 1018 444 1020
rect 466 1018 468 1020
rect 472 1018 474 1020
rect 496 1018 498 1020
rect 502 1018 504 1020
rect 526 1018 528 1020
rect 532 1018 534 1020
rect 74 1016 76 1018
rect 104 1016 106 1018
rect 134 1016 136 1018
rect 164 1016 166 1018
rect 194 1016 196 1018
rect 224 1016 226 1018
rect 254 1016 256 1018
rect 284 1016 286 1018
rect 314 1016 316 1018
rect 344 1016 346 1018
rect 374 1016 376 1018
rect 404 1016 406 1018
rect 434 1016 436 1018
rect 464 1016 466 1018
rect 494 1016 496 1018
rect 524 1016 526 1018
rect 74 1010 76 1012
rect 104 1010 106 1012
rect 134 1010 136 1012
rect 164 1010 166 1012
rect 194 1010 196 1012
rect 224 1010 226 1012
rect 254 1010 256 1012
rect 284 1010 286 1012
rect 314 1010 316 1012
rect 344 1010 346 1012
rect 374 1010 376 1012
rect 404 1010 406 1012
rect 434 1010 436 1012
rect 464 1010 466 1012
rect 494 1010 496 1012
rect 524 1010 526 1012
rect 76 1008 78 1010
rect 82 1008 84 1010
rect 106 1008 108 1010
rect 112 1008 114 1010
rect 136 1008 138 1010
rect 142 1008 144 1010
rect 166 1008 168 1010
rect 172 1008 174 1010
rect 196 1008 198 1010
rect 202 1008 204 1010
rect 226 1008 228 1010
rect 232 1008 234 1010
rect 256 1008 258 1010
rect 262 1008 264 1010
rect 286 1008 288 1010
rect 292 1008 294 1010
rect 316 1008 318 1010
rect 322 1008 324 1010
rect 346 1008 348 1010
rect 352 1008 354 1010
rect 376 1008 378 1010
rect 382 1008 384 1010
rect 406 1008 408 1010
rect 412 1008 414 1010
rect 436 1008 438 1010
rect 442 1008 444 1010
rect 466 1008 468 1010
rect 472 1008 474 1010
rect 496 1008 498 1010
rect 502 1008 504 1010
rect 526 1008 528 1010
rect 532 1008 534 1010
rect 84 1006 86 1008
rect 114 1006 116 1008
rect 144 1006 146 1008
rect 174 1006 176 1008
rect 204 1006 206 1008
rect 234 1006 236 1008
rect 264 1006 266 1008
rect 294 1006 296 1008
rect 324 1006 326 1008
rect 354 1006 356 1008
rect 384 1006 386 1008
rect 414 1006 416 1008
rect 444 1006 446 1008
rect 474 1006 476 1008
rect 504 1006 506 1008
rect 534 1006 536 1008
rect 84 1000 86 1002
rect 114 1000 116 1002
rect 144 1000 146 1002
rect 174 1000 176 1002
rect 204 1000 206 1002
rect 234 1000 236 1002
rect 264 1000 266 1002
rect 294 1000 296 1002
rect 324 1000 326 1002
rect 354 1000 356 1002
rect 384 1000 386 1002
rect 414 1000 416 1002
rect 444 1000 446 1002
rect 474 1000 476 1002
rect 504 1000 506 1002
rect 534 1000 536 1002
rect 76 998 78 1000
rect 82 998 84 1000
rect 106 998 108 1000
rect 112 998 114 1000
rect 136 998 138 1000
rect 142 998 144 1000
rect 166 998 168 1000
rect 172 998 174 1000
rect 196 998 198 1000
rect 202 998 204 1000
rect 226 998 228 1000
rect 232 998 234 1000
rect 256 998 258 1000
rect 262 998 264 1000
rect 286 998 288 1000
rect 292 998 294 1000
rect 316 998 318 1000
rect 322 998 324 1000
rect 346 998 348 1000
rect 352 998 354 1000
rect 376 998 378 1000
rect 382 998 384 1000
rect 406 998 408 1000
rect 412 998 414 1000
rect 436 998 438 1000
rect 442 998 444 1000
rect 466 998 468 1000
rect 472 998 474 1000
rect 496 998 498 1000
rect 502 998 504 1000
rect 526 998 528 1000
rect 532 998 534 1000
rect 74 996 76 998
rect 104 996 106 998
rect 134 996 136 998
rect 164 996 166 998
rect 194 996 196 998
rect 224 996 226 998
rect 254 996 256 998
rect 284 996 286 998
rect 314 996 316 998
rect 344 996 346 998
rect 374 996 376 998
rect 404 996 406 998
rect 434 996 436 998
rect 464 996 466 998
rect 494 996 496 998
rect 524 996 526 998
rect 74 990 76 992
rect 104 990 106 992
rect 134 990 136 992
rect 164 990 166 992
rect 194 990 196 992
rect 224 990 226 992
rect 254 990 256 992
rect 284 990 286 992
rect 314 990 316 992
rect 344 990 346 992
rect 374 990 376 992
rect 404 990 406 992
rect 434 990 436 992
rect 464 990 466 992
rect 494 990 496 992
rect 524 990 526 992
rect 76 988 78 990
rect 82 988 84 990
rect 106 988 108 990
rect 112 988 114 990
rect 136 988 138 990
rect 142 988 144 990
rect 166 988 168 990
rect 172 988 174 990
rect 196 988 198 990
rect 202 988 204 990
rect 226 988 228 990
rect 232 988 234 990
rect 256 988 258 990
rect 262 988 264 990
rect 286 988 288 990
rect 292 988 294 990
rect 316 988 318 990
rect 322 988 324 990
rect 346 988 348 990
rect 352 988 354 990
rect 376 988 378 990
rect 382 988 384 990
rect 406 988 408 990
rect 412 988 414 990
rect 436 988 438 990
rect 442 988 444 990
rect 466 988 468 990
rect 472 988 474 990
rect 496 988 498 990
rect 502 988 504 990
rect 526 988 528 990
rect 532 988 534 990
rect 84 986 86 988
rect 114 986 116 988
rect 144 986 146 988
rect 174 986 176 988
rect 204 986 206 988
rect 234 986 236 988
rect 264 986 266 988
rect 294 986 296 988
rect 324 986 326 988
rect 354 986 356 988
rect 384 986 386 988
rect 414 986 416 988
rect 444 986 446 988
rect 474 986 476 988
rect 504 986 506 988
rect 534 986 536 988
rect 84 980 86 982
rect 114 980 116 982
rect 144 980 146 982
rect 174 980 176 982
rect 204 980 206 982
rect 234 980 236 982
rect 264 980 266 982
rect 294 980 296 982
rect 324 980 326 982
rect 354 980 356 982
rect 384 980 386 982
rect 414 980 416 982
rect 444 980 446 982
rect 474 980 476 982
rect 504 980 506 982
rect 534 980 536 982
rect 76 978 78 980
rect 82 978 84 980
rect 106 978 108 980
rect 112 978 114 980
rect 136 978 138 980
rect 142 978 144 980
rect 166 978 168 980
rect 172 978 174 980
rect 196 978 198 980
rect 202 978 204 980
rect 226 978 228 980
rect 232 978 234 980
rect 256 978 258 980
rect 262 978 264 980
rect 286 978 288 980
rect 292 978 294 980
rect 316 978 318 980
rect 322 978 324 980
rect 346 978 348 980
rect 352 978 354 980
rect 376 978 378 980
rect 382 978 384 980
rect 406 978 408 980
rect 412 978 414 980
rect 436 978 438 980
rect 442 978 444 980
rect 466 978 468 980
rect 472 978 474 980
rect 496 978 498 980
rect 502 978 504 980
rect 526 978 528 980
rect 532 978 534 980
rect 74 976 76 978
rect 104 976 106 978
rect 134 976 136 978
rect 164 976 166 978
rect 194 976 196 978
rect 224 976 226 978
rect 254 976 256 978
rect 284 976 286 978
rect 314 976 316 978
rect 344 976 346 978
rect 374 976 376 978
rect 404 976 406 978
rect 434 976 436 978
rect 464 976 466 978
rect 494 976 496 978
rect 524 976 526 978
rect 74 950 76 952
rect 104 950 106 952
rect 134 950 136 952
rect 164 950 166 952
rect 194 950 196 952
rect 224 950 226 952
rect 254 950 256 952
rect 284 950 286 952
rect 314 950 316 952
rect 344 950 346 952
rect 374 950 376 952
rect 404 950 406 952
rect 434 950 436 952
rect 464 950 466 952
rect 494 950 496 952
rect 524 950 526 952
rect 76 948 78 950
rect 82 948 84 950
rect 106 948 108 950
rect 112 948 114 950
rect 136 948 138 950
rect 142 948 144 950
rect 166 948 168 950
rect 172 948 174 950
rect 196 948 198 950
rect 202 948 204 950
rect 226 948 228 950
rect 232 948 234 950
rect 256 948 258 950
rect 262 948 264 950
rect 286 948 288 950
rect 292 948 294 950
rect 316 948 318 950
rect 322 948 324 950
rect 346 948 348 950
rect 352 948 354 950
rect 376 948 378 950
rect 382 948 384 950
rect 406 948 408 950
rect 412 948 414 950
rect 436 948 438 950
rect 442 948 444 950
rect 466 948 468 950
rect 472 948 474 950
rect 496 948 498 950
rect 502 948 504 950
rect 526 948 528 950
rect 532 948 534 950
rect 84 946 86 948
rect 114 946 116 948
rect 144 946 146 948
rect 174 946 176 948
rect 204 946 206 948
rect 234 946 236 948
rect 264 946 266 948
rect 294 946 296 948
rect 324 946 326 948
rect 354 946 356 948
rect 384 946 386 948
rect 414 946 416 948
rect 444 946 446 948
rect 474 946 476 948
rect 504 946 506 948
rect 534 946 536 948
rect 84 940 86 942
rect 114 940 116 942
rect 144 940 146 942
rect 174 940 176 942
rect 204 940 206 942
rect 234 940 236 942
rect 264 940 266 942
rect 294 940 296 942
rect 324 940 326 942
rect 354 940 356 942
rect 384 940 386 942
rect 414 940 416 942
rect 444 940 446 942
rect 474 940 476 942
rect 504 940 506 942
rect 534 940 536 942
rect 76 938 78 940
rect 82 938 84 940
rect 106 938 108 940
rect 112 938 114 940
rect 136 938 138 940
rect 142 938 144 940
rect 166 938 168 940
rect 172 938 174 940
rect 196 938 198 940
rect 202 938 204 940
rect 226 938 228 940
rect 232 938 234 940
rect 256 938 258 940
rect 262 938 264 940
rect 286 938 288 940
rect 292 938 294 940
rect 316 938 318 940
rect 322 938 324 940
rect 346 938 348 940
rect 352 938 354 940
rect 376 938 378 940
rect 382 938 384 940
rect 406 938 408 940
rect 412 938 414 940
rect 436 938 438 940
rect 442 938 444 940
rect 466 938 468 940
rect 472 938 474 940
rect 496 938 498 940
rect 502 938 504 940
rect 526 938 528 940
rect 532 938 534 940
rect 74 936 76 938
rect 104 936 106 938
rect 134 936 136 938
rect 164 936 166 938
rect 194 936 196 938
rect 224 936 226 938
rect 254 936 256 938
rect 284 936 286 938
rect 314 936 316 938
rect 344 936 346 938
rect 374 936 376 938
rect 404 936 406 938
rect 434 936 436 938
rect 464 936 466 938
rect 494 936 496 938
rect 524 936 526 938
rect 74 930 76 932
rect 104 930 106 932
rect 134 930 136 932
rect 164 930 166 932
rect 194 930 196 932
rect 224 930 226 932
rect 254 930 256 932
rect 284 930 286 932
rect 314 930 316 932
rect 344 930 346 932
rect 374 930 376 932
rect 404 930 406 932
rect 434 930 436 932
rect 464 930 466 932
rect 494 930 496 932
rect 524 930 526 932
rect 76 928 78 930
rect 82 928 84 930
rect 106 928 108 930
rect 112 928 114 930
rect 136 928 138 930
rect 142 928 144 930
rect 166 928 168 930
rect 172 928 174 930
rect 196 928 198 930
rect 202 928 204 930
rect 226 928 228 930
rect 232 928 234 930
rect 256 928 258 930
rect 262 928 264 930
rect 286 928 288 930
rect 292 928 294 930
rect 316 928 318 930
rect 322 928 324 930
rect 346 928 348 930
rect 352 928 354 930
rect 376 928 378 930
rect 382 928 384 930
rect 406 928 408 930
rect 412 928 414 930
rect 436 928 438 930
rect 442 928 444 930
rect 466 928 468 930
rect 472 928 474 930
rect 496 928 498 930
rect 502 928 504 930
rect 526 928 528 930
rect 532 928 534 930
rect 84 926 86 928
rect 114 926 116 928
rect 144 926 146 928
rect 174 926 176 928
rect 204 926 206 928
rect 234 926 236 928
rect 264 926 266 928
rect 294 926 296 928
rect 324 926 326 928
rect 354 926 356 928
rect 384 926 386 928
rect 414 926 416 928
rect 444 926 446 928
rect 474 926 476 928
rect 504 926 506 928
rect 534 926 536 928
rect 84 920 86 922
rect 114 920 116 922
rect 144 920 146 922
rect 174 920 176 922
rect 204 920 206 922
rect 234 920 236 922
rect 264 920 266 922
rect 294 920 296 922
rect 324 920 326 922
rect 354 920 356 922
rect 384 920 386 922
rect 414 920 416 922
rect 444 920 446 922
rect 474 920 476 922
rect 504 920 506 922
rect 534 920 536 922
rect 76 918 78 920
rect 82 918 84 920
rect 106 918 108 920
rect 112 918 114 920
rect 136 918 138 920
rect 142 918 144 920
rect 166 918 168 920
rect 172 918 174 920
rect 196 918 198 920
rect 202 918 204 920
rect 226 918 228 920
rect 232 918 234 920
rect 256 918 258 920
rect 262 918 264 920
rect 286 918 288 920
rect 292 918 294 920
rect 316 918 318 920
rect 322 918 324 920
rect 346 918 348 920
rect 352 918 354 920
rect 376 918 378 920
rect 382 918 384 920
rect 406 918 408 920
rect 412 918 414 920
rect 436 918 438 920
rect 442 918 444 920
rect 466 918 468 920
rect 472 918 474 920
rect 496 918 498 920
rect 502 918 504 920
rect 526 918 528 920
rect 532 918 534 920
rect 74 916 76 918
rect 104 916 106 918
rect 134 916 136 918
rect 164 916 166 918
rect 194 916 196 918
rect 224 916 226 918
rect 254 916 256 918
rect 284 916 286 918
rect 314 916 316 918
rect 344 916 346 918
rect 374 916 376 918
rect 404 916 406 918
rect 434 916 436 918
rect 464 916 466 918
rect 494 916 496 918
rect 524 916 526 918
rect 74 910 76 912
rect 104 910 106 912
rect 134 910 136 912
rect 164 910 166 912
rect 194 910 196 912
rect 224 910 226 912
rect 254 910 256 912
rect 284 910 286 912
rect 314 910 316 912
rect 344 910 346 912
rect 374 910 376 912
rect 404 910 406 912
rect 434 910 436 912
rect 464 910 466 912
rect 494 910 496 912
rect 524 910 526 912
rect 76 908 78 910
rect 82 908 84 910
rect 106 908 108 910
rect 112 908 114 910
rect 136 908 138 910
rect 142 908 144 910
rect 166 908 168 910
rect 172 908 174 910
rect 196 908 198 910
rect 202 908 204 910
rect 226 908 228 910
rect 232 908 234 910
rect 256 908 258 910
rect 262 908 264 910
rect 286 908 288 910
rect 292 908 294 910
rect 316 908 318 910
rect 322 908 324 910
rect 346 908 348 910
rect 352 908 354 910
rect 376 908 378 910
rect 382 908 384 910
rect 406 908 408 910
rect 412 908 414 910
rect 436 908 438 910
rect 442 908 444 910
rect 466 908 468 910
rect 472 908 474 910
rect 496 908 498 910
rect 502 908 504 910
rect 526 908 528 910
rect 532 908 534 910
rect 84 906 86 908
rect 114 906 116 908
rect 144 906 146 908
rect 174 906 176 908
rect 204 906 206 908
rect 234 906 236 908
rect 264 906 266 908
rect 294 906 296 908
rect 324 906 326 908
rect 354 906 356 908
rect 384 906 386 908
rect 414 906 416 908
rect 444 906 446 908
rect 474 906 476 908
rect 504 906 506 908
rect 534 906 536 908
rect 84 900 86 902
rect 114 900 116 902
rect 144 900 146 902
rect 174 900 176 902
rect 204 900 206 902
rect 234 900 236 902
rect 264 900 266 902
rect 294 900 296 902
rect 324 900 326 902
rect 354 900 356 902
rect 384 900 386 902
rect 414 900 416 902
rect 444 900 446 902
rect 474 900 476 902
rect 504 900 506 902
rect 534 900 536 902
rect 76 898 78 900
rect 82 898 84 900
rect 106 898 108 900
rect 112 898 114 900
rect 136 898 138 900
rect 142 898 144 900
rect 166 898 168 900
rect 172 898 174 900
rect 196 898 198 900
rect 202 898 204 900
rect 226 898 228 900
rect 232 898 234 900
rect 256 898 258 900
rect 262 898 264 900
rect 286 898 288 900
rect 292 898 294 900
rect 316 898 318 900
rect 322 898 324 900
rect 346 898 348 900
rect 352 898 354 900
rect 376 898 378 900
rect 382 898 384 900
rect 406 898 408 900
rect 412 898 414 900
rect 436 898 438 900
rect 442 898 444 900
rect 466 898 468 900
rect 472 898 474 900
rect 496 898 498 900
rect 502 898 504 900
rect 526 898 528 900
rect 532 898 534 900
rect 74 896 76 898
rect 104 896 106 898
rect 134 896 136 898
rect 164 896 166 898
rect 194 896 196 898
rect 224 896 226 898
rect 254 896 256 898
rect 284 896 286 898
rect 314 896 316 898
rect 344 896 346 898
rect 374 896 376 898
rect 404 896 406 898
rect 434 896 436 898
rect 464 896 466 898
rect 494 896 496 898
rect 524 896 526 898
rect 74 890 76 892
rect 104 890 106 892
rect 134 890 136 892
rect 164 890 166 892
rect 194 890 196 892
rect 224 890 226 892
rect 254 890 256 892
rect 284 890 286 892
rect 314 890 316 892
rect 344 890 346 892
rect 374 890 376 892
rect 404 890 406 892
rect 434 890 436 892
rect 464 890 466 892
rect 494 890 496 892
rect 524 890 526 892
rect 76 888 78 890
rect 82 888 84 890
rect 106 888 108 890
rect 112 888 114 890
rect 136 888 138 890
rect 142 888 144 890
rect 166 888 168 890
rect 172 888 174 890
rect 196 888 198 890
rect 202 888 204 890
rect 226 888 228 890
rect 232 888 234 890
rect 256 888 258 890
rect 262 888 264 890
rect 286 888 288 890
rect 292 888 294 890
rect 316 888 318 890
rect 322 888 324 890
rect 346 888 348 890
rect 352 888 354 890
rect 376 888 378 890
rect 382 888 384 890
rect 406 888 408 890
rect 412 888 414 890
rect 436 888 438 890
rect 442 888 444 890
rect 466 888 468 890
rect 472 888 474 890
rect 496 888 498 890
rect 502 888 504 890
rect 526 888 528 890
rect 532 888 534 890
rect 84 886 86 888
rect 114 886 116 888
rect 144 886 146 888
rect 174 886 176 888
rect 204 886 206 888
rect 234 886 236 888
rect 264 886 266 888
rect 294 886 296 888
rect 324 886 326 888
rect 354 886 356 888
rect 384 886 386 888
rect 414 886 416 888
rect 444 886 446 888
rect 474 886 476 888
rect 504 886 506 888
rect 534 886 536 888
rect 56 878 58 880
rect 62 878 64 880
rect 76 878 78 880
rect 92 878 94 880
rect 106 878 108 880
rect 122 878 124 880
rect 136 878 138 880
rect 152 878 154 880
rect 166 878 168 880
rect 182 878 184 880
rect 196 878 198 880
rect 212 878 214 880
rect 226 878 228 880
rect 242 878 244 880
rect 256 878 258 880
rect 272 878 274 880
rect 286 878 288 880
rect 302 878 304 880
rect 316 878 318 880
rect 332 878 334 880
rect 346 878 348 880
rect 362 878 364 880
rect 376 878 378 880
rect 392 878 394 880
rect 406 878 408 880
rect 422 878 424 880
rect 436 878 438 880
rect 452 878 454 880
rect 466 878 468 880
rect 482 878 484 880
rect 496 878 498 880
rect 512 878 514 880
rect 526 878 528 880
rect 542 878 544 880
rect 54 876 56 878
rect 64 876 66 878
rect 74 876 76 878
rect 94 876 96 878
rect 104 876 106 878
rect 124 876 126 878
rect 134 876 136 878
rect 154 876 156 878
rect 164 876 166 878
rect 184 876 186 878
rect 194 876 196 878
rect 214 876 216 878
rect 224 876 226 878
rect 244 876 246 878
rect 254 876 256 878
rect 274 876 276 878
rect 284 876 286 878
rect 304 876 306 878
rect 314 876 316 878
rect 334 876 336 878
rect 344 876 346 878
rect 364 876 366 878
rect 374 876 376 878
rect 394 876 396 878
rect 404 876 406 878
rect 424 876 426 878
rect 434 876 436 878
rect 454 876 456 878
rect 464 876 466 878
rect 484 876 486 878
rect 494 876 496 878
rect 514 876 516 878
rect 524 876 526 878
rect 544 876 546 878
rect 32 828 34 830
rect 62 828 64 830
rect 92 828 94 830
rect 122 828 124 830
rect 152 828 154 830
rect 446 828 448 830
rect 476 828 478 830
rect 506 828 508 830
rect 536 828 538 830
rect 566 828 568 830
rect 34 826 36 828
rect 40 826 42 828
rect 64 826 66 828
rect 70 826 72 828
rect 94 826 96 828
rect 100 826 102 828
rect 124 826 126 828
rect 130 826 132 828
rect 154 826 156 828
rect 160 826 162 828
rect 438 826 440 828
rect 444 826 446 828
rect 468 826 470 828
rect 474 826 476 828
rect 498 826 500 828
rect 504 826 506 828
rect 528 826 530 828
rect 534 826 536 828
rect 558 826 560 828
rect 564 826 566 828
rect 42 824 44 826
rect 72 824 74 826
rect 102 824 104 826
rect 132 824 134 826
rect 162 824 164 826
rect 436 824 438 826
rect 466 824 468 826
rect 496 824 498 826
rect 526 824 528 826
rect 556 824 558 826
rect 42 818 44 820
rect 72 818 74 820
rect 102 818 104 820
rect 132 818 134 820
rect 162 818 164 820
rect 436 818 438 820
rect 466 818 468 820
rect 496 818 498 820
rect 526 818 528 820
rect 556 818 558 820
rect 34 816 36 818
rect 40 816 42 818
rect 64 816 66 818
rect 70 816 72 818
rect 94 816 96 818
rect 100 816 102 818
rect 124 816 126 818
rect 130 816 132 818
rect 154 816 156 818
rect 160 816 162 818
rect 438 816 440 818
rect 444 816 446 818
rect 468 816 470 818
rect 474 816 476 818
rect 498 816 500 818
rect 504 816 506 818
rect 528 816 530 818
rect 534 816 536 818
rect 558 816 560 818
rect 564 816 566 818
rect 32 814 34 816
rect 62 814 64 816
rect 92 814 94 816
rect 122 814 124 816
rect 152 814 154 816
rect 446 814 448 816
rect 476 814 478 816
rect 506 814 508 816
rect 536 814 538 816
rect 566 814 568 816
rect 32 808 34 810
rect 62 808 64 810
rect 92 808 94 810
rect 122 808 124 810
rect 152 808 154 810
rect 446 808 448 810
rect 476 808 478 810
rect 506 808 508 810
rect 536 808 538 810
rect 566 808 568 810
rect 34 806 36 808
rect 40 806 42 808
rect 64 806 66 808
rect 70 806 72 808
rect 94 806 96 808
rect 100 806 102 808
rect 124 806 126 808
rect 130 806 132 808
rect 154 806 156 808
rect 160 806 162 808
rect 438 806 440 808
rect 444 806 446 808
rect 468 806 470 808
rect 474 806 476 808
rect 498 806 500 808
rect 504 806 506 808
rect 528 806 530 808
rect 534 806 536 808
rect 558 806 560 808
rect 564 806 566 808
rect 42 804 44 806
rect 72 804 74 806
rect 102 804 104 806
rect 132 804 134 806
rect 162 804 164 806
rect 436 804 438 806
rect 466 804 468 806
rect 496 804 498 806
rect 526 804 528 806
rect 556 804 558 806
rect 42 798 44 800
rect 72 798 74 800
rect 102 798 104 800
rect 132 798 134 800
rect 162 798 164 800
rect 436 798 438 800
rect 466 798 468 800
rect 496 798 498 800
rect 526 798 528 800
rect 556 798 558 800
rect 34 796 36 798
rect 40 796 42 798
rect 64 796 66 798
rect 70 796 72 798
rect 94 796 96 798
rect 100 796 102 798
rect 124 796 126 798
rect 130 796 132 798
rect 154 796 156 798
rect 160 796 162 798
rect 438 796 440 798
rect 444 796 446 798
rect 468 796 470 798
rect 474 796 476 798
rect 498 796 500 798
rect 504 796 506 798
rect 528 796 530 798
rect 534 796 536 798
rect 558 796 560 798
rect 564 796 566 798
rect 32 794 34 796
rect 62 794 64 796
rect 92 794 94 796
rect 122 794 124 796
rect 152 794 154 796
rect 446 794 448 796
rect 476 794 478 796
rect 506 794 508 796
rect 536 794 538 796
rect 566 794 568 796
rect 32 788 34 790
rect 62 788 64 790
rect 92 788 94 790
rect 122 788 124 790
rect 152 788 154 790
rect 446 788 448 790
rect 476 788 478 790
rect 506 788 508 790
rect 536 788 538 790
rect 566 788 568 790
rect 34 786 36 788
rect 40 786 42 788
rect 64 786 66 788
rect 70 786 72 788
rect 94 786 96 788
rect 100 786 102 788
rect 124 786 126 788
rect 130 786 132 788
rect 154 786 156 788
rect 160 786 162 788
rect 438 786 440 788
rect 444 786 446 788
rect 468 786 470 788
rect 474 786 476 788
rect 498 786 500 788
rect 504 786 506 788
rect 528 786 530 788
rect 534 786 536 788
rect 558 786 560 788
rect 564 786 566 788
rect 42 784 44 786
rect 72 784 74 786
rect 102 784 104 786
rect 132 784 134 786
rect 162 784 164 786
rect 436 784 438 786
rect 466 784 468 786
rect 496 784 498 786
rect 526 784 528 786
rect 556 784 558 786
rect 42 778 44 780
rect 72 778 74 780
rect 526 778 528 780
rect 556 778 558 780
rect 34 776 36 778
rect 40 776 42 778
rect 64 776 66 778
rect 70 776 72 778
rect 94 776 96 778
rect 110 776 112 778
rect 124 776 126 778
rect 140 776 142 778
rect 154 776 156 778
rect 170 776 172 778
rect 184 776 186 778
rect 292 776 294 778
rect 306 776 308 778
rect 414 776 416 778
rect 428 776 430 778
rect 444 776 446 778
rect 458 776 460 778
rect 474 776 476 778
rect 488 776 490 778
rect 504 776 506 778
rect 528 776 530 778
rect 534 776 536 778
rect 558 776 560 778
rect 564 776 566 778
rect 32 774 34 776
rect 62 774 64 776
rect 92 774 94 776
rect 112 774 114 776
rect 122 774 124 776
rect 142 774 144 776
rect 152 774 154 776
rect 172 774 174 776
rect 182 774 184 776
rect 294 774 296 776
rect 304 774 306 776
rect 416 774 418 776
rect 426 774 428 776
rect 446 774 448 776
rect 456 774 458 776
rect 476 774 478 776
rect 486 774 488 776
rect 506 774 508 776
rect 536 774 538 776
rect 566 774 568 776
rect 32 768 34 770
rect 62 768 64 770
rect 92 768 94 770
rect 112 768 114 770
rect 122 768 124 770
rect 142 768 144 770
rect 152 768 154 770
rect 172 768 174 770
rect 182 768 184 770
rect 294 768 296 770
rect 304 768 306 770
rect 416 768 418 770
rect 426 768 428 770
rect 446 768 448 770
rect 456 768 458 770
rect 476 768 478 770
rect 486 768 488 770
rect 506 768 508 770
rect 536 768 538 770
rect 566 768 568 770
rect 34 766 36 768
rect 40 766 42 768
rect 64 766 66 768
rect 70 766 72 768
rect 94 766 96 768
rect 110 766 112 768
rect 124 766 126 768
rect 140 766 142 768
rect 154 766 156 768
rect 170 766 172 768
rect 184 766 186 768
rect 296 766 298 768
rect 302 766 304 768
rect 414 766 416 768
rect 428 766 430 768
rect 444 766 446 768
rect 458 766 460 768
rect 474 766 476 768
rect 488 766 490 768
rect 504 766 506 768
rect 528 766 530 768
rect 534 766 536 768
rect 558 766 560 768
rect 564 766 566 768
rect 42 764 44 766
rect 72 764 74 766
rect 526 764 528 766
rect 556 764 558 766
rect 42 758 44 760
rect 72 758 74 760
rect 102 758 104 760
rect 132 758 134 760
rect 162 758 164 760
rect 436 758 438 760
rect 466 758 468 760
rect 496 758 498 760
rect 526 758 528 760
rect 556 758 558 760
rect 34 756 36 758
rect 40 756 42 758
rect 64 756 66 758
rect 70 756 72 758
rect 94 756 96 758
rect 100 756 102 758
rect 124 756 126 758
rect 130 756 132 758
rect 154 756 156 758
rect 160 756 162 758
rect 438 756 440 758
rect 444 756 446 758
rect 468 756 470 758
rect 474 756 476 758
rect 498 756 500 758
rect 504 756 506 758
rect 528 756 530 758
rect 534 756 536 758
rect 558 756 560 758
rect 564 756 566 758
rect 32 754 34 756
rect 62 754 64 756
rect 92 754 94 756
rect 122 754 124 756
rect 152 754 154 756
rect 446 754 448 756
rect 476 754 478 756
rect 506 754 508 756
rect 536 754 538 756
rect 566 754 568 756
rect 32 748 34 750
rect 62 748 64 750
rect 92 748 94 750
rect 122 748 124 750
rect 152 748 154 750
rect 446 748 448 750
rect 476 748 478 750
rect 506 748 508 750
rect 536 748 538 750
rect 566 748 568 750
rect 34 746 36 748
rect 40 746 42 748
rect 64 746 66 748
rect 70 746 72 748
rect 94 746 96 748
rect 100 746 102 748
rect 124 746 126 748
rect 130 746 132 748
rect 154 746 156 748
rect 160 746 162 748
rect 438 746 440 748
rect 444 746 446 748
rect 468 746 470 748
rect 474 746 476 748
rect 498 746 500 748
rect 504 746 506 748
rect 528 746 530 748
rect 534 746 536 748
rect 558 746 560 748
rect 564 746 566 748
rect 42 744 44 746
rect 72 744 74 746
rect 102 744 104 746
rect 132 744 134 746
rect 162 744 164 746
rect 436 744 438 746
rect 466 744 468 746
rect 496 744 498 746
rect 526 744 528 746
rect 556 744 558 746
rect 42 718 44 720
rect 72 718 74 720
rect 102 718 104 720
rect 132 718 134 720
rect 162 718 164 720
rect 436 718 438 720
rect 466 718 468 720
rect 496 718 498 720
rect 526 718 528 720
rect 556 718 558 720
rect 34 716 36 718
rect 40 716 42 718
rect 64 716 66 718
rect 70 716 72 718
rect 94 716 96 718
rect 100 716 102 718
rect 124 716 126 718
rect 130 716 132 718
rect 154 716 156 718
rect 160 716 162 718
rect 438 716 440 718
rect 444 716 446 718
rect 468 716 470 718
rect 474 716 476 718
rect 498 716 500 718
rect 504 716 506 718
rect 528 716 530 718
rect 534 716 536 718
rect 558 716 560 718
rect 564 716 566 718
rect 32 714 34 716
rect 62 714 64 716
rect 92 714 94 716
rect 122 714 124 716
rect 152 714 154 716
rect 446 714 448 716
rect 476 714 478 716
rect 506 714 508 716
rect 536 714 538 716
rect 566 714 568 716
rect 32 708 34 710
rect 62 708 64 710
rect 92 708 94 710
rect 122 708 124 710
rect 152 708 154 710
rect 446 708 448 710
rect 476 708 478 710
rect 506 708 508 710
rect 536 708 538 710
rect 566 708 568 710
rect 34 706 36 708
rect 40 706 42 708
rect 64 706 66 708
rect 70 706 72 708
rect 94 706 96 708
rect 100 706 102 708
rect 124 706 126 708
rect 130 706 132 708
rect 154 706 156 708
rect 160 706 162 708
rect 296 706 298 708
rect 302 706 304 708
rect 438 706 440 708
rect 444 706 446 708
rect 468 706 470 708
rect 474 706 476 708
rect 498 706 500 708
rect 504 706 506 708
rect 528 706 530 708
rect 534 706 536 708
rect 558 706 560 708
rect 564 706 566 708
rect 42 704 44 706
rect 72 704 74 706
rect 102 704 104 706
rect 132 704 134 706
rect 162 704 164 706
rect 294 704 296 706
rect 304 704 306 706
rect 436 704 438 706
rect 466 704 468 706
rect 496 704 498 706
rect 526 704 528 706
rect 556 704 558 706
rect 42 698 44 700
rect 72 698 74 700
rect 102 698 104 700
rect 132 698 134 700
rect 162 698 164 700
rect 436 698 438 700
rect 466 698 468 700
rect 496 698 498 700
rect 526 698 528 700
rect 556 698 558 700
rect 34 696 36 698
rect 40 696 42 698
rect 64 696 66 698
rect 70 696 72 698
rect 94 696 96 698
rect 100 696 102 698
rect 124 696 126 698
rect 130 696 132 698
rect 154 696 156 698
rect 160 696 162 698
rect 438 696 440 698
rect 444 696 446 698
rect 468 696 470 698
rect 474 696 476 698
rect 498 696 500 698
rect 504 696 506 698
rect 528 696 530 698
rect 534 696 536 698
rect 558 696 560 698
rect 564 696 566 698
rect 32 694 34 696
rect 62 694 64 696
rect 92 694 94 696
rect 122 694 124 696
rect 152 694 154 696
rect 446 694 448 696
rect 476 694 478 696
rect 506 694 508 696
rect 536 694 538 696
rect 566 694 568 696
rect 32 644 34 646
rect 62 644 64 646
rect 92 644 94 646
rect 122 644 124 646
rect 152 644 154 646
rect 182 644 184 646
rect 212 644 214 646
rect 284 644 286 646
rect 314 644 316 646
rect 386 644 388 646
rect 416 644 418 646
rect 446 644 448 646
rect 476 644 478 646
rect 506 644 508 646
rect 536 644 538 646
rect 566 644 568 646
rect 34 642 36 644
rect 40 642 42 644
rect 64 642 66 644
rect 70 642 72 644
rect 94 642 96 644
rect 100 642 102 644
rect 124 642 126 644
rect 130 642 132 644
rect 154 642 156 644
rect 160 642 162 644
rect 184 642 186 644
rect 190 642 192 644
rect 214 642 216 644
rect 220 642 222 644
rect 286 642 288 644
rect 292 642 294 644
rect 316 642 318 644
rect 322 642 324 644
rect 378 642 380 644
rect 384 642 386 644
rect 408 642 410 644
rect 414 642 416 644
rect 438 642 440 644
rect 444 642 446 644
rect 468 642 470 644
rect 474 642 476 644
rect 498 642 500 644
rect 504 642 506 644
rect 528 642 530 644
rect 534 642 536 644
rect 558 642 560 644
rect 564 642 566 644
rect 42 640 44 642
rect 72 640 74 642
rect 102 640 104 642
rect 132 640 134 642
rect 162 640 164 642
rect 192 640 194 642
rect 222 640 224 642
rect 294 640 296 642
rect 324 640 326 642
rect 376 640 378 642
rect 406 640 408 642
rect 436 640 438 642
rect 466 640 468 642
rect 496 640 498 642
rect 526 640 528 642
rect 556 640 558 642
rect 42 634 44 636
rect 72 634 74 636
rect 102 634 104 636
rect 132 634 134 636
rect 162 634 164 636
rect 192 634 194 636
rect 222 634 224 636
rect 294 634 296 636
rect 324 634 326 636
rect 376 634 378 636
rect 406 634 408 636
rect 436 634 438 636
rect 466 634 468 636
rect 496 634 498 636
rect 526 634 528 636
rect 556 634 558 636
rect 34 632 36 634
rect 40 632 42 634
rect 64 632 66 634
rect 70 632 72 634
rect 94 632 96 634
rect 100 632 102 634
rect 124 632 126 634
rect 130 632 132 634
rect 154 632 156 634
rect 160 632 162 634
rect 184 632 186 634
rect 190 632 192 634
rect 214 632 216 634
rect 220 632 222 634
rect 286 632 288 634
rect 292 632 294 634
rect 316 632 318 634
rect 322 632 324 634
rect 378 632 380 634
rect 384 632 386 634
rect 408 632 410 634
rect 414 632 416 634
rect 438 632 440 634
rect 444 632 446 634
rect 468 632 470 634
rect 474 632 476 634
rect 498 632 500 634
rect 504 632 506 634
rect 528 632 530 634
rect 534 632 536 634
rect 558 632 560 634
rect 564 632 566 634
rect 32 630 34 632
rect 62 630 64 632
rect 92 630 94 632
rect 122 630 124 632
rect 152 630 154 632
rect 182 630 184 632
rect 212 630 214 632
rect 284 630 286 632
rect 314 630 316 632
rect 386 630 388 632
rect 416 630 418 632
rect 446 630 448 632
rect 476 630 478 632
rect 506 630 508 632
rect 536 630 538 632
rect 566 630 568 632
rect 32 624 34 626
rect 62 624 64 626
rect 92 624 94 626
rect 122 624 124 626
rect 152 624 154 626
rect 182 624 184 626
rect 212 624 214 626
rect 284 624 286 626
rect 314 624 316 626
rect 386 624 388 626
rect 416 624 418 626
rect 446 624 448 626
rect 476 624 478 626
rect 506 624 508 626
rect 536 624 538 626
rect 566 624 568 626
rect 34 622 36 624
rect 40 622 42 624
rect 64 622 66 624
rect 70 622 72 624
rect 94 622 96 624
rect 100 622 102 624
rect 124 622 126 624
rect 130 622 132 624
rect 154 622 156 624
rect 160 622 162 624
rect 184 622 186 624
rect 190 622 192 624
rect 214 622 216 624
rect 220 622 222 624
rect 286 622 288 624
rect 292 622 294 624
rect 316 622 318 624
rect 322 622 324 624
rect 378 622 380 624
rect 384 622 386 624
rect 408 622 410 624
rect 414 622 416 624
rect 438 622 440 624
rect 444 622 446 624
rect 468 622 470 624
rect 474 622 476 624
rect 498 622 500 624
rect 504 622 506 624
rect 528 622 530 624
rect 534 622 536 624
rect 558 622 560 624
rect 564 622 566 624
rect 42 620 44 622
rect 72 620 74 622
rect 102 620 104 622
rect 132 620 134 622
rect 162 620 164 622
rect 192 620 194 622
rect 222 620 224 622
rect 294 620 296 622
rect 324 620 326 622
rect 376 620 378 622
rect 406 620 408 622
rect 436 620 438 622
rect 466 620 468 622
rect 496 620 498 622
rect 526 620 528 622
rect 556 620 558 622
rect 222 614 224 616
rect 294 614 296 616
rect 324 614 326 616
rect 376 614 378 616
rect 220 612 222 614
rect 286 612 288 614
rect 292 612 294 614
rect 316 612 318 614
rect 322 612 324 614
rect 378 612 380 614
rect 284 610 286 612
rect 314 610 316 612
rect 284 604 286 606
rect 314 604 316 606
rect 220 602 222 604
rect 286 602 288 604
rect 292 602 294 604
rect 316 602 318 604
rect 322 602 324 604
rect 378 602 380 604
rect 222 600 224 602
rect 294 600 296 602
rect 324 600 326 602
rect 376 600 378 602
rect 42 594 44 596
rect 72 594 74 596
rect 102 594 104 596
rect 132 594 134 596
rect 162 594 164 596
rect 192 594 194 596
rect 222 594 224 596
rect 376 594 378 596
rect 406 594 408 596
rect 436 594 438 596
rect 466 594 468 596
rect 496 594 498 596
rect 526 594 528 596
rect 556 594 558 596
rect 34 592 36 594
rect 40 592 42 594
rect 64 592 66 594
rect 70 592 72 594
rect 94 592 96 594
rect 100 592 102 594
rect 124 592 126 594
rect 130 592 132 594
rect 154 592 156 594
rect 160 592 162 594
rect 184 592 186 594
rect 190 592 192 594
rect 214 592 216 594
rect 220 592 222 594
rect 266 592 268 594
rect 272 592 274 594
rect 286 592 288 594
rect 302 592 304 594
rect 316 592 318 594
rect 332 592 334 594
rect 378 592 380 594
rect 384 592 386 594
rect 408 592 410 594
rect 414 592 416 594
rect 438 592 440 594
rect 444 592 446 594
rect 468 592 470 594
rect 474 592 476 594
rect 498 592 500 594
rect 504 592 506 594
rect 528 592 530 594
rect 534 592 536 594
rect 558 592 560 594
rect 564 592 566 594
rect 32 590 34 592
rect 62 590 64 592
rect 92 590 94 592
rect 122 590 124 592
rect 152 590 154 592
rect 182 590 184 592
rect 212 590 214 592
rect 264 590 266 592
rect 274 590 276 592
rect 284 590 286 592
rect 304 590 306 592
rect 314 590 316 592
rect 334 590 336 592
rect 386 590 388 592
rect 416 590 418 592
rect 446 590 448 592
rect 476 590 478 592
rect 506 590 508 592
rect 536 590 538 592
rect 566 590 568 592
rect 32 584 34 586
rect 62 584 64 586
rect 92 584 94 586
rect 506 584 508 586
rect 536 584 538 586
rect 566 584 568 586
rect 34 582 36 584
rect 40 582 42 584
rect 64 582 66 584
rect 70 582 72 584
rect 94 582 96 584
rect 100 582 102 584
rect 114 582 116 584
rect 130 582 132 584
rect 144 582 146 584
rect 160 582 162 584
rect 174 582 176 584
rect 190 582 192 584
rect 204 582 206 584
rect 220 582 222 584
rect 234 582 236 584
rect 240 582 242 584
rect 358 582 360 584
rect 364 582 366 584
rect 378 582 380 584
rect 394 582 396 584
rect 408 582 410 584
rect 424 582 426 584
rect 438 582 440 584
rect 454 582 456 584
rect 468 582 470 584
rect 484 582 486 584
rect 498 582 500 584
rect 504 582 506 584
rect 528 582 530 584
rect 534 582 536 584
rect 558 582 560 584
rect 564 582 566 584
rect 42 580 44 582
rect 72 580 74 582
rect 102 580 104 582
rect 112 580 114 582
rect 132 580 134 582
rect 142 580 144 582
rect 162 580 164 582
rect 172 580 174 582
rect 192 580 194 582
rect 202 580 204 582
rect 222 580 224 582
rect 232 580 234 582
rect 242 580 244 582
rect 356 580 358 582
rect 366 580 368 582
rect 376 580 378 582
rect 396 580 398 582
rect 406 580 408 582
rect 426 580 428 582
rect 436 580 438 582
rect 456 580 458 582
rect 466 580 468 582
rect 486 580 488 582
rect 496 580 498 582
rect 526 580 528 582
rect 556 580 558 582
rect 42 574 44 576
rect 72 574 74 576
rect 102 574 104 576
rect 112 574 114 576
rect 132 574 134 576
rect 142 574 144 576
rect 162 574 164 576
rect 172 574 174 576
rect 192 574 194 576
rect 202 574 204 576
rect 222 574 224 576
rect 232 574 234 576
rect 242 574 244 576
rect 264 574 266 576
rect 274 574 276 576
rect 294 574 296 576
rect 304 574 306 576
rect 324 574 326 576
rect 334 574 336 576
rect 356 574 358 576
rect 366 574 368 576
rect 376 574 378 576
rect 396 574 398 576
rect 406 574 408 576
rect 426 574 428 576
rect 436 574 438 576
rect 456 574 458 576
rect 466 574 468 576
rect 486 574 488 576
rect 496 574 498 576
rect 526 574 528 576
rect 556 574 558 576
rect 34 572 36 574
rect 40 572 42 574
rect 64 572 66 574
rect 70 572 72 574
rect 94 572 96 574
rect 100 572 102 574
rect 114 572 116 574
rect 130 572 132 574
rect 144 572 146 574
rect 160 572 162 574
rect 174 572 176 574
rect 190 572 192 574
rect 204 572 206 574
rect 220 572 222 574
rect 234 572 236 574
rect 240 572 242 574
rect 262 572 264 574
rect 276 572 278 574
rect 292 572 294 574
rect 306 572 308 574
rect 322 572 324 574
rect 336 572 338 574
rect 358 572 360 574
rect 364 572 366 574
rect 378 572 380 574
rect 394 572 396 574
rect 408 572 410 574
rect 424 572 426 574
rect 438 572 440 574
rect 454 572 456 574
rect 468 572 470 574
rect 484 572 486 574
rect 498 572 500 574
rect 504 572 506 574
rect 528 572 530 574
rect 534 572 536 574
rect 558 572 560 574
rect 564 572 566 574
rect 32 570 34 572
rect 62 570 64 572
rect 92 570 94 572
rect 506 570 508 572
rect 536 570 538 572
rect 566 570 568 572
rect 32 564 34 566
rect 62 564 64 566
rect 92 564 94 566
rect 122 564 124 566
rect 152 564 154 566
rect 182 564 184 566
rect 212 564 214 566
rect 284 564 286 566
rect 314 564 316 566
rect 386 564 388 566
rect 416 564 418 566
rect 446 564 448 566
rect 476 564 478 566
rect 506 564 508 566
rect 536 564 538 566
rect 566 564 568 566
rect 34 562 36 564
rect 40 562 42 564
rect 64 562 66 564
rect 70 562 72 564
rect 94 562 96 564
rect 100 562 102 564
rect 124 562 126 564
rect 130 562 132 564
rect 154 562 156 564
rect 160 562 162 564
rect 184 562 186 564
rect 190 562 192 564
rect 214 562 216 564
rect 220 562 222 564
rect 286 562 288 564
rect 292 562 294 564
rect 316 562 318 564
rect 322 562 324 564
rect 378 562 380 564
rect 384 562 386 564
rect 408 562 410 564
rect 414 562 416 564
rect 438 562 440 564
rect 444 562 446 564
rect 468 562 470 564
rect 474 562 476 564
rect 498 562 500 564
rect 504 562 506 564
rect 528 562 530 564
rect 534 562 536 564
rect 558 562 560 564
rect 564 562 566 564
rect 42 560 44 562
rect 72 560 74 562
rect 102 560 104 562
rect 132 560 134 562
rect 162 560 164 562
rect 192 560 194 562
rect 222 560 224 562
rect 294 560 296 562
rect 324 560 326 562
rect 376 560 378 562
rect 406 560 408 562
rect 436 560 438 562
rect 466 560 468 562
rect 496 560 498 562
rect 526 560 528 562
rect 556 560 558 562
rect 42 554 44 556
rect 72 554 74 556
rect 102 554 104 556
rect 132 554 134 556
rect 162 554 164 556
rect 192 554 194 556
rect 222 554 224 556
rect 294 554 296 556
rect 324 554 326 556
rect 376 554 378 556
rect 406 554 408 556
rect 436 554 438 556
rect 466 554 468 556
rect 496 554 498 556
rect 526 554 528 556
rect 556 554 558 556
rect 34 552 36 554
rect 40 552 42 554
rect 64 552 66 554
rect 70 552 72 554
rect 94 552 96 554
rect 100 552 102 554
rect 124 552 126 554
rect 130 552 132 554
rect 154 552 156 554
rect 160 552 162 554
rect 184 552 186 554
rect 190 552 192 554
rect 214 552 216 554
rect 220 552 222 554
rect 286 552 288 554
rect 292 552 294 554
rect 316 552 318 554
rect 322 552 324 554
rect 378 552 380 554
rect 384 552 386 554
rect 408 552 410 554
rect 414 552 416 554
rect 438 552 440 554
rect 444 552 446 554
rect 468 552 470 554
rect 474 552 476 554
rect 498 552 500 554
rect 504 552 506 554
rect 528 552 530 554
rect 534 552 536 554
rect 558 552 560 554
rect 564 552 566 554
rect 32 550 34 552
rect 62 550 64 552
rect 92 550 94 552
rect 122 550 124 552
rect 152 550 154 552
rect 182 550 184 552
rect 212 550 214 552
rect 284 550 286 552
rect 314 550 316 552
rect 386 550 388 552
rect 416 550 418 552
rect 446 550 448 552
rect 476 550 478 552
rect 506 550 508 552
rect 536 550 538 552
rect 566 550 568 552
rect 32 544 34 546
rect 62 544 64 546
rect 92 544 94 546
rect 122 544 124 546
rect 152 544 154 546
rect 182 544 184 546
rect 212 544 214 546
rect 284 544 286 546
rect 314 544 316 546
rect 386 544 388 546
rect 416 544 418 546
rect 446 544 448 546
rect 476 544 478 546
rect 506 544 508 546
rect 536 544 538 546
rect 566 544 568 546
rect 34 542 36 544
rect 40 542 42 544
rect 64 542 66 544
rect 70 542 72 544
rect 94 542 96 544
rect 100 542 102 544
rect 124 542 126 544
rect 130 542 132 544
rect 154 542 156 544
rect 160 542 162 544
rect 184 542 186 544
rect 190 542 192 544
rect 214 542 216 544
rect 220 542 222 544
rect 286 542 288 544
rect 292 542 294 544
rect 316 542 318 544
rect 322 542 324 544
rect 378 542 380 544
rect 384 542 386 544
rect 408 542 410 544
rect 414 542 416 544
rect 438 542 440 544
rect 444 542 446 544
rect 468 542 470 544
rect 474 542 476 544
rect 498 542 500 544
rect 504 542 506 544
rect 528 542 530 544
rect 534 542 536 544
rect 558 542 560 544
rect 564 542 566 544
rect 42 540 44 542
rect 72 540 74 542
rect 102 540 104 542
rect 132 540 134 542
rect 162 540 164 542
rect 192 540 194 542
rect 222 540 224 542
rect 294 540 296 542
rect 324 540 326 542
rect 376 540 378 542
rect 406 540 408 542
rect 436 540 438 542
rect 466 540 468 542
rect 496 540 498 542
rect 526 540 528 542
rect 556 540 558 542
rect 42 534 44 536
rect 72 534 74 536
rect 102 534 104 536
rect 132 534 134 536
rect 162 534 164 536
rect 192 534 194 536
rect 222 534 224 536
rect 294 534 296 536
rect 324 534 326 536
rect 376 534 378 536
rect 406 534 408 536
rect 436 534 438 536
rect 466 534 468 536
rect 496 534 498 536
rect 526 534 528 536
rect 556 534 558 536
rect 34 532 36 534
rect 40 532 42 534
rect 64 532 66 534
rect 70 532 72 534
rect 94 532 96 534
rect 100 532 102 534
rect 124 532 126 534
rect 130 532 132 534
rect 154 532 156 534
rect 160 532 162 534
rect 184 532 186 534
rect 190 532 192 534
rect 214 532 216 534
rect 220 532 222 534
rect 286 532 288 534
rect 292 532 294 534
rect 316 532 318 534
rect 322 532 324 534
rect 378 532 380 534
rect 384 532 386 534
rect 408 532 410 534
rect 414 532 416 534
rect 438 532 440 534
rect 444 532 446 534
rect 468 532 470 534
rect 474 532 476 534
rect 498 532 500 534
rect 504 532 506 534
rect 528 532 530 534
rect 534 532 536 534
rect 558 532 560 534
rect 564 532 566 534
rect 32 530 34 532
rect 62 530 64 532
rect 92 530 94 532
rect 122 530 124 532
rect 152 530 154 532
rect 182 530 184 532
rect 212 530 214 532
rect 284 530 286 532
rect 314 530 316 532
rect 386 530 388 532
rect 416 530 418 532
rect 446 530 448 532
rect 476 530 478 532
rect 506 530 508 532
rect 536 530 538 532
rect 566 530 568 532
rect 586 508 588 510
rect 588 506 590 508
rect 56 466 58 468
rect 76 466 78 468
rect 522 466 524 468
rect 542 466 544 468
rect 54 464 56 466
rect 78 464 80 466
rect 520 464 522 466
rect 544 464 546 466
rect 106 420 108 422
rect 492 420 494 422
rect 104 418 106 420
rect 494 418 496 420
rect 104 356 106 358
rect 494 356 496 358
rect 106 354 108 356
rect 492 354 494 356
rect 106 288 108 290
rect 492 288 494 290
rect 104 286 106 288
rect 494 286 496 288
rect 104 226 106 228
rect 494 226 496 228
rect 106 224 108 226
rect 492 224 494 226
rect 106 158 108 160
rect 492 158 494 160
rect 104 156 106 158
rect 494 156 496 158
rect 104 96 106 98
rect 494 96 496 98
rect 106 94 108 96
rect 492 94 494 96
rect 86 56 88 58
rect 96 56 98 58
rect 106 56 108 58
rect 116 56 118 58
rect 126 56 128 58
rect 136 56 138 58
rect 146 56 148 58
rect 156 56 158 58
rect 166 56 168 58
rect 176 56 178 58
rect 186 56 188 58
rect 412 56 414 58
rect 422 56 424 58
rect 432 56 434 58
rect 442 56 444 58
rect 452 56 454 58
rect 462 56 464 58
rect 472 56 474 58
rect 482 56 484 58
rect 492 56 494 58
rect 502 56 504 58
rect 512 56 514 58
rect 84 54 86 56
rect 98 54 100 56
rect 104 54 106 56
rect 118 54 120 56
rect 124 54 126 56
rect 138 54 140 56
rect 144 54 146 56
rect 158 54 160 56
rect 164 54 166 56
rect 178 54 180 56
rect 184 54 186 56
rect 414 54 416 56
rect 420 54 422 56
rect 434 54 436 56
rect 440 54 442 56
rect 454 54 456 56
rect 460 54 462 56
rect 474 54 476 56
rect 480 54 482 56
rect 494 54 496 56
rect 500 54 502 56
rect 514 54 516 56
rect 12 14 22 16
rect 10 12 22 14
rect 578 14 588 16
rect 578 12 590 14
rect 12 8 14 12
rect 586 8 588 12
rect 14 6 16 8
rect 584 6 586 8
<< error_s >>
rect 110 1598 118 1600
rect 134 1598 142 1600
rect 158 1598 166 1600
rect 182 1598 190 1600
rect 206 1598 214 1600
rect 230 1598 238 1600
rect 254 1598 262 1600
rect 278 1598 286 1600
rect 302 1598 310 1600
rect 326 1598 334 1600
rect 350 1598 358 1600
rect 374 1598 382 1600
rect 398 1598 406 1600
rect 422 1598 430 1600
rect 446 1598 454 1600
rect 470 1598 478 1600
rect 494 1598 502 1600
rect 98 1592 106 1594
rect 98 1588 100 1592
rect 104 1588 106 1592
rect 98 1586 106 1588
rect 122 1592 130 1594
rect 122 1588 124 1592
rect 128 1588 130 1592
rect 122 1586 130 1588
rect 146 1592 154 1594
rect 146 1588 148 1592
rect 152 1588 154 1592
rect 146 1586 154 1588
rect 170 1592 178 1594
rect 170 1588 172 1592
rect 176 1588 178 1592
rect 170 1586 178 1588
rect 194 1592 202 1594
rect 194 1588 196 1592
rect 200 1588 202 1592
rect 194 1586 202 1588
rect 218 1592 226 1594
rect 218 1588 220 1592
rect 224 1588 226 1592
rect 218 1586 226 1588
rect 242 1592 250 1594
rect 242 1588 244 1592
rect 248 1588 250 1592
rect 242 1586 250 1588
rect 266 1592 274 1594
rect 266 1588 268 1592
rect 272 1588 274 1592
rect 266 1586 274 1588
rect 290 1592 298 1594
rect 290 1588 292 1592
rect 296 1588 298 1592
rect 290 1586 298 1588
rect 314 1592 322 1594
rect 314 1588 316 1592
rect 320 1588 322 1592
rect 314 1586 322 1588
rect 338 1592 346 1594
rect 338 1588 340 1592
rect 344 1588 346 1592
rect 338 1586 346 1588
rect 362 1592 370 1594
rect 362 1588 364 1592
rect 368 1588 370 1592
rect 362 1586 370 1588
rect 386 1592 394 1594
rect 386 1588 388 1592
rect 392 1588 394 1592
rect 386 1586 394 1588
rect 410 1592 418 1594
rect 410 1588 412 1592
rect 416 1588 418 1592
rect 410 1586 418 1588
rect 434 1592 442 1594
rect 434 1588 436 1592
rect 440 1588 442 1592
rect 434 1586 442 1588
rect 458 1592 466 1594
rect 458 1588 460 1592
rect 464 1588 466 1592
rect 458 1586 466 1588
rect 482 1592 490 1594
rect 482 1588 484 1592
rect 488 1588 490 1592
rect 482 1586 490 1588
rect 110 1580 118 1582
rect 110 1576 112 1580
rect 116 1576 118 1580
rect 110 1574 118 1576
rect 134 1580 142 1582
rect 134 1576 136 1580
rect 140 1576 142 1580
rect 134 1574 142 1576
rect 158 1580 166 1582
rect 158 1576 160 1580
rect 164 1576 166 1580
rect 158 1574 166 1576
rect 182 1580 190 1582
rect 182 1576 184 1580
rect 188 1576 190 1580
rect 182 1574 190 1576
rect 206 1580 214 1582
rect 206 1576 208 1580
rect 212 1576 214 1580
rect 206 1574 214 1576
rect 230 1580 238 1582
rect 230 1576 232 1580
rect 236 1576 238 1580
rect 230 1574 238 1576
rect 254 1580 262 1582
rect 254 1576 256 1580
rect 260 1576 262 1580
rect 254 1574 262 1576
rect 278 1580 286 1582
rect 278 1576 280 1580
rect 284 1576 286 1580
rect 278 1574 286 1576
rect 302 1580 310 1582
rect 302 1576 304 1580
rect 308 1576 310 1580
rect 302 1574 310 1576
rect 326 1580 334 1582
rect 326 1576 328 1580
rect 332 1576 334 1580
rect 326 1574 334 1576
rect 350 1580 358 1582
rect 350 1576 352 1580
rect 356 1576 358 1580
rect 350 1574 358 1576
rect 374 1580 382 1582
rect 374 1576 376 1580
rect 380 1576 382 1580
rect 374 1574 382 1576
rect 398 1580 406 1582
rect 398 1576 400 1580
rect 404 1576 406 1580
rect 398 1574 406 1576
rect 422 1580 430 1582
rect 422 1576 424 1580
rect 428 1576 430 1580
rect 422 1574 430 1576
rect 446 1580 454 1582
rect 446 1576 448 1580
rect 452 1576 454 1580
rect 446 1574 454 1576
rect 470 1580 478 1582
rect 470 1576 472 1580
rect 476 1576 478 1580
rect 470 1574 478 1576
rect 494 1580 502 1582
rect 494 1576 496 1580
rect 500 1576 502 1580
rect 494 1574 502 1576
rect 98 1568 106 1570
rect 98 1564 100 1568
rect 104 1564 106 1568
rect 98 1562 106 1564
rect 122 1568 130 1570
rect 122 1564 124 1568
rect 128 1564 130 1568
rect 122 1562 130 1564
rect 146 1568 154 1570
rect 146 1564 148 1568
rect 152 1564 154 1568
rect 146 1562 154 1564
rect 170 1568 178 1570
rect 170 1564 172 1568
rect 176 1564 178 1568
rect 170 1562 178 1564
rect 194 1568 202 1570
rect 194 1564 196 1568
rect 200 1564 202 1568
rect 194 1562 202 1564
rect 218 1568 226 1570
rect 218 1564 220 1568
rect 224 1564 226 1568
rect 218 1562 226 1564
rect 242 1568 250 1570
rect 242 1564 244 1568
rect 248 1564 250 1568
rect 242 1562 250 1564
rect 266 1568 274 1570
rect 266 1564 268 1568
rect 272 1564 274 1568
rect 266 1562 274 1564
rect 290 1568 298 1570
rect 290 1564 292 1568
rect 296 1564 298 1568
rect 290 1562 298 1564
rect 314 1568 322 1570
rect 314 1564 316 1568
rect 320 1564 322 1568
rect 314 1562 322 1564
rect 338 1568 346 1570
rect 338 1564 340 1568
rect 344 1564 346 1568
rect 338 1562 346 1564
rect 362 1568 370 1570
rect 362 1564 364 1568
rect 368 1564 370 1568
rect 362 1562 370 1564
rect 386 1568 394 1570
rect 386 1564 388 1568
rect 392 1564 394 1568
rect 386 1562 394 1564
rect 410 1568 418 1570
rect 410 1564 412 1568
rect 416 1564 418 1568
rect 410 1562 418 1564
rect 434 1568 442 1570
rect 434 1564 436 1568
rect 440 1564 442 1568
rect 434 1562 442 1564
rect 458 1568 466 1570
rect 458 1564 460 1568
rect 464 1564 466 1568
rect 458 1562 466 1564
rect 482 1568 490 1570
rect 482 1564 484 1568
rect 488 1564 490 1568
rect 482 1562 490 1564
rect 110 1556 118 1558
rect 110 1552 112 1556
rect 116 1552 118 1556
rect 110 1550 118 1552
rect 134 1556 142 1558
rect 134 1552 136 1556
rect 140 1552 142 1556
rect 134 1550 142 1552
rect 158 1556 166 1558
rect 158 1552 160 1556
rect 164 1552 166 1556
rect 158 1550 166 1552
rect 182 1556 190 1558
rect 182 1552 184 1556
rect 188 1552 190 1556
rect 182 1550 190 1552
rect 206 1556 214 1558
rect 206 1552 208 1556
rect 212 1552 214 1556
rect 206 1550 214 1552
rect 230 1556 238 1558
rect 230 1552 232 1556
rect 236 1552 238 1556
rect 230 1550 238 1552
rect 254 1556 262 1558
rect 254 1552 256 1556
rect 260 1552 262 1556
rect 254 1550 262 1552
rect 278 1556 286 1558
rect 278 1552 280 1556
rect 284 1552 286 1556
rect 278 1550 286 1552
rect 302 1556 310 1558
rect 302 1552 304 1556
rect 308 1552 310 1556
rect 302 1550 310 1552
rect 326 1556 334 1558
rect 326 1552 328 1556
rect 332 1552 334 1556
rect 326 1550 334 1552
rect 350 1556 358 1558
rect 350 1552 352 1556
rect 356 1552 358 1556
rect 350 1550 358 1552
rect 374 1556 382 1558
rect 374 1552 376 1556
rect 380 1552 382 1556
rect 374 1550 382 1552
rect 398 1556 406 1558
rect 398 1552 400 1556
rect 404 1552 406 1556
rect 398 1550 406 1552
rect 422 1556 430 1558
rect 422 1552 424 1556
rect 428 1552 430 1556
rect 422 1550 430 1552
rect 446 1556 454 1558
rect 446 1552 448 1556
rect 452 1552 454 1556
rect 446 1550 454 1552
rect 470 1556 478 1558
rect 470 1552 472 1556
rect 476 1552 478 1556
rect 470 1550 478 1552
rect 494 1556 502 1558
rect 494 1552 496 1556
rect 500 1552 502 1556
rect 494 1550 502 1552
rect 98 1544 106 1546
rect 98 1540 100 1544
rect 104 1540 106 1544
rect 98 1538 106 1540
rect 122 1544 130 1546
rect 122 1540 124 1544
rect 128 1540 130 1544
rect 122 1538 130 1540
rect 146 1544 154 1546
rect 146 1540 148 1544
rect 152 1540 154 1544
rect 146 1538 154 1540
rect 170 1544 178 1546
rect 170 1540 172 1544
rect 176 1540 178 1544
rect 170 1538 178 1540
rect 194 1544 202 1546
rect 194 1540 196 1544
rect 200 1540 202 1544
rect 194 1538 202 1540
rect 218 1544 226 1546
rect 218 1540 220 1544
rect 224 1540 226 1544
rect 218 1538 226 1540
rect 242 1544 250 1546
rect 242 1540 244 1544
rect 248 1540 250 1544
rect 242 1538 250 1540
rect 266 1544 274 1546
rect 266 1540 268 1544
rect 272 1540 274 1544
rect 266 1538 274 1540
rect 290 1544 298 1546
rect 290 1540 292 1544
rect 296 1540 298 1544
rect 290 1538 298 1540
rect 314 1544 322 1546
rect 314 1540 316 1544
rect 320 1540 322 1544
rect 314 1538 322 1540
rect 338 1544 346 1546
rect 338 1540 340 1544
rect 344 1540 346 1544
rect 338 1538 346 1540
rect 362 1544 370 1546
rect 362 1540 364 1544
rect 368 1540 370 1544
rect 362 1538 370 1540
rect 386 1544 394 1546
rect 386 1540 388 1544
rect 392 1540 394 1544
rect 386 1538 394 1540
rect 410 1544 418 1546
rect 410 1540 412 1544
rect 416 1540 418 1544
rect 410 1538 418 1540
rect 434 1544 442 1546
rect 434 1540 436 1544
rect 440 1540 442 1544
rect 434 1538 442 1540
rect 458 1544 466 1546
rect 458 1540 460 1544
rect 464 1540 466 1544
rect 458 1538 466 1540
rect 482 1544 490 1546
rect 482 1540 484 1544
rect 488 1540 490 1544
rect 482 1538 490 1540
<< nwell >>
rect 34 858 566 1306
rect -6 496 606 660
rect -6 20 22 496
rect 578 20 606 496
rect -6 -8 606 20
<< ntransistor >>
rect 76 430 276 436
rect 324 430 524 436
rect 76 340 276 346
rect 76 298 276 304
rect 324 340 524 346
rect 324 298 524 304
rect 76 210 276 216
rect 76 168 276 174
rect 324 210 524 216
rect 324 168 524 174
rect 76 80 276 86
rect 324 80 524 86
<< ndiffusion >>
rect 76 452 276 454
rect 76 444 82 452
rect 190 444 276 452
rect 76 436 276 444
rect 324 452 524 454
rect 324 444 410 452
rect 518 444 524 452
rect 324 436 524 444
rect 76 398 276 430
rect 76 390 112 398
rect 240 390 276 398
rect 76 386 276 390
rect 76 378 112 386
rect 240 378 276 386
rect 76 346 276 378
rect 76 332 276 340
rect 76 324 82 332
rect 240 324 276 332
rect 76 320 276 324
rect 76 312 82 320
rect 240 312 276 320
rect 76 304 276 312
rect 76 266 276 298
rect 76 248 112 266
rect 240 248 276 266
rect 76 216 276 248
rect 324 398 524 430
rect 324 390 360 398
rect 488 390 524 398
rect 324 386 524 390
rect 324 378 360 386
rect 488 378 524 386
rect 324 346 524 378
rect 324 332 524 340
rect 324 324 360 332
rect 518 324 524 332
rect 324 320 524 324
rect 324 312 360 320
rect 518 312 524 320
rect 324 304 524 312
rect 76 202 276 210
rect 76 194 82 202
rect 240 194 276 202
rect 76 190 276 194
rect 76 182 82 190
rect 240 182 276 190
rect 76 174 276 182
rect 76 136 276 168
rect 76 118 112 136
rect 240 118 276 136
rect 76 86 276 118
rect 324 266 524 298
rect 324 248 360 266
rect 488 248 524 266
rect 324 216 524 248
rect 324 202 524 210
rect 324 194 360 202
rect 518 194 524 202
rect 324 190 524 194
rect 324 182 360 190
rect 518 182 524 190
rect 324 174 524 182
rect 324 136 524 168
rect 324 118 360 136
rect 488 118 524 136
rect 324 86 524 118
rect 76 72 276 80
rect 76 64 82 72
rect 190 64 276 72
rect 76 62 276 64
rect 324 72 524 80
rect 324 64 410 72
rect 518 64 524 72
rect 324 62 524 64
<< ndcontact >>
rect 82 444 190 452
rect 410 444 518 452
rect 112 390 240 398
rect 112 378 240 386
rect 82 324 240 332
rect 82 312 240 320
rect 112 248 240 266
rect 360 390 488 398
rect 360 378 488 386
rect 360 324 518 332
rect 360 312 518 320
rect 82 194 240 202
rect 82 182 240 190
rect 112 118 240 136
rect 360 248 488 266
rect 360 194 518 202
rect 360 182 518 190
rect 360 118 488 136
rect 82 64 190 72
rect 410 64 518 72
<< psubstratepdiff >>
rect 0 1338 600 1340
rect 0 840 2 1338
rect 190 1320 408 1338
rect 576 1320 580 1338
rect 20 1318 580 1320
rect 20 846 22 1318
rect 578 846 580 1318
rect 20 840 580 846
rect 598 840 600 1338
rect 0 836 600 840
rect 0 828 4 836
rect 12 828 24 836
rect 42 828 54 836
rect 72 828 84 836
rect 102 828 114 836
rect 132 828 144 836
rect 162 828 174 836
rect 182 828 296 836
rect 304 828 418 836
rect 426 828 438 836
rect 456 828 468 836
rect 486 828 498 836
rect 516 828 528 836
rect 546 828 558 836
rect 576 828 588 836
rect 596 828 600 836
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 0 818 14 826
rect 22 818 34 826
rect 52 818 64 826
rect 82 818 94 826
rect 112 818 124 826
rect 142 818 154 826
rect 172 818 184 826
rect 192 818 286 826
rect 294 818 306 826
rect 314 818 408 826
rect 416 818 428 826
rect 446 818 458 826
rect 476 818 488 826
rect 506 818 518 826
rect 536 818 548 826
rect 566 818 578 826
rect 586 818 600 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 0 808 4 816
rect 12 808 24 816
rect 42 808 54 816
rect 72 808 84 816
rect 102 808 114 816
rect 132 808 144 816
rect 162 808 174 816
rect 182 808 296 816
rect 304 808 418 816
rect 426 808 438 816
rect 456 808 468 816
rect 486 808 498 816
rect 516 808 528 816
rect 546 808 558 816
rect 576 808 588 816
rect 596 808 600 816
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 0 798 14 806
rect 22 798 34 806
rect 52 798 64 806
rect 82 798 94 806
rect 112 798 124 806
rect 142 798 154 806
rect 172 798 184 806
rect 192 798 286 806
rect 294 798 306 806
rect 314 798 408 806
rect 416 798 428 806
rect 446 798 458 806
rect 476 798 488 806
rect 506 798 518 806
rect 536 798 548 806
rect 566 798 578 806
rect 586 798 600 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 0 788 4 796
rect 12 788 24 796
rect 42 788 54 796
rect 72 788 84 796
rect 102 788 114 796
rect 132 788 144 796
rect 162 788 174 796
rect 182 788 296 796
rect 304 788 418 796
rect 426 788 438 796
rect 456 788 468 796
rect 486 788 498 796
rect 516 788 528 796
rect 546 788 558 796
rect 576 788 588 796
rect 596 788 600 796
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 0 778 14 786
rect 22 778 34 786
rect 52 778 64 786
rect 82 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 776 124 786
rect 142 776 154 786
rect 172 776 184 786
rect 0 768 4 776
rect 12 768 24 776
rect 42 768 54 776
rect 72 768 84 776
rect 192 768 286 786
rect 294 776 306 786
rect 314 768 408 786
rect 416 776 428 786
rect 446 776 458 786
rect 476 776 488 786
rect 506 778 518 786
rect 536 778 548 786
rect 566 778 578 786
rect 586 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 516 768 528 776
rect 546 768 558 776
rect 576 768 588 776
rect 596 768 600 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 14 766
rect 22 758 34 766
rect 52 758 64 766
rect 82 758 94 766
rect 112 758 124 768
rect 142 758 154 768
rect 172 758 184 768
rect 192 758 296 768
rect 304 758 408 768
rect 416 758 428 768
rect 446 758 458 768
rect 476 758 488 768
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 518 766
rect 536 758 548 766
rect 566 758 578 766
rect 586 758 600 766
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 0 748 4 756
rect 12 748 24 756
rect 42 748 54 756
rect 72 748 84 756
rect 102 748 114 756
rect 132 748 144 756
rect 162 748 174 756
rect 182 748 286 756
rect 294 748 306 756
rect 314 748 418 756
rect 426 748 438 756
rect 456 748 468 756
rect 486 748 498 756
rect 516 748 528 756
rect 546 748 558 756
rect 576 748 588 756
rect 596 748 600 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 0 738 14 746
rect 22 738 34 746
rect 52 738 64 746
rect 82 738 94 746
rect 112 738 124 746
rect 142 738 154 746
rect 172 738 184 746
rect 192 738 296 746
rect 304 738 408 746
rect 416 738 428 746
rect 446 738 458 746
rect 476 738 488 746
rect 506 738 518 746
rect 536 738 548 746
rect 566 738 578 746
rect 586 738 600 746
rect 0 736 600 738
rect 0 728 4 736
rect 12 728 24 736
rect 32 728 286 736
rect 294 728 306 736
rect 314 728 568 736
rect 576 728 588 736
rect 596 728 600 736
rect 0 726 600 728
rect 0 718 14 726
rect 22 718 34 726
rect 52 718 64 726
rect 82 718 94 726
rect 112 718 124 726
rect 142 718 154 726
rect 172 718 184 726
rect 192 718 296 726
rect 304 718 408 726
rect 416 718 428 726
rect 446 718 458 726
rect 476 718 488 726
rect 506 718 518 726
rect 536 718 548 726
rect 566 718 578 726
rect 586 718 600 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 0 708 4 716
rect 12 708 24 716
rect 42 708 54 716
rect 72 708 84 716
rect 102 708 114 716
rect 132 708 144 716
rect 162 708 174 716
rect 182 708 286 716
rect 294 708 306 716
rect 314 708 418 716
rect 426 708 438 716
rect 456 708 468 716
rect 486 708 498 716
rect 516 708 528 716
rect 546 708 558 716
rect 576 708 588 716
rect 596 708 600 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 0 698 14 706
rect 22 698 34 706
rect 52 698 64 706
rect 82 698 94 706
rect 112 698 124 706
rect 142 698 154 706
rect 172 698 184 706
rect 192 698 408 706
rect 416 698 428 706
rect 446 698 458 706
rect 476 698 488 706
rect 506 698 518 706
rect 536 698 548 706
rect 566 698 578 706
rect 586 698 600 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 0 688 4 696
rect 12 688 24 696
rect 42 688 54 696
rect 72 688 84 696
rect 102 688 114 696
rect 132 688 144 696
rect 162 688 174 696
rect 182 688 286 696
rect 314 688 418 696
rect 426 688 438 696
rect 456 688 468 696
rect 486 688 498 696
rect 516 688 528 696
rect 546 688 558 696
rect 576 688 588 696
rect 596 688 600 696
rect 0 686 600 688
rect 28 484 572 490
rect 28 456 38 484
rect 56 458 78 466
rect 56 456 60 458
rect 28 444 60 456
rect 28 436 38 444
rect 56 436 60 444
rect 76 456 78 458
rect 196 458 404 484
rect 196 456 276 458
rect 76 454 276 456
rect 284 444 316 458
rect 284 436 291 444
rect 309 436 316 444
rect 324 456 404 458
rect 522 458 544 466
rect 522 456 524 458
rect 324 454 524 456
rect 540 456 544 458
rect 562 456 572 484
rect 540 444 572 456
rect 540 436 544 444
rect 562 436 572 444
rect 28 424 60 436
rect 28 416 38 424
rect 56 416 60 424
rect 28 404 60 416
rect 28 396 38 404
rect 56 396 60 404
rect 28 384 60 396
rect 28 376 38 384
rect 56 376 60 384
rect 28 364 60 376
rect 28 356 38 364
rect 56 356 60 364
rect 28 344 60 356
rect 28 336 38 344
rect 56 336 60 344
rect 28 324 60 336
rect 28 316 38 324
rect 56 316 60 324
rect 28 304 60 316
rect 28 296 38 304
rect 56 296 60 304
rect 28 284 60 296
rect 28 276 38 284
rect 56 276 60 284
rect 28 264 60 276
rect 28 256 38 264
rect 56 256 60 264
rect 28 244 60 256
rect 28 236 38 244
rect 56 236 60 244
rect 28 224 60 236
rect 28 216 38 224
rect 56 216 60 224
rect 28 204 60 216
rect 28 196 38 204
rect 56 196 60 204
rect 28 184 60 196
rect 28 176 38 184
rect 56 176 60 184
rect 28 164 60 176
rect 28 156 38 164
rect 56 156 60 164
rect 28 144 60 156
rect 28 136 38 144
rect 56 136 60 144
rect 28 124 60 136
rect 28 116 38 124
rect 56 116 60 124
rect 28 104 60 116
rect 28 96 38 104
rect 56 96 60 104
rect 28 84 60 96
rect 28 76 38 84
rect 56 76 60 84
rect 284 428 316 436
rect 284 420 291 428
rect 309 420 316 428
rect 284 412 316 420
rect 284 404 291 412
rect 309 404 316 412
rect 284 268 316 404
rect 284 260 291 268
rect 309 260 316 268
rect 284 252 316 260
rect 284 244 291 252
rect 309 244 316 252
rect 284 124 316 244
rect 284 116 291 124
rect 309 116 316 124
rect 284 108 316 116
rect 284 100 291 108
rect 309 100 316 108
rect 284 92 316 100
rect 284 84 291 92
rect 309 84 316 92
rect 28 64 60 76
rect 28 56 38 64
rect 56 58 60 64
rect 76 58 276 62
rect 284 76 316 84
rect 540 424 572 436
rect 540 416 544 424
rect 562 416 572 424
rect 540 404 572 416
rect 540 396 544 404
rect 562 396 572 404
rect 540 384 572 396
rect 540 376 544 384
rect 562 376 572 384
rect 540 364 572 376
rect 540 356 544 364
rect 562 356 572 364
rect 540 344 572 356
rect 540 336 544 344
rect 562 336 572 344
rect 540 324 572 336
rect 540 316 544 324
rect 562 316 572 324
rect 540 304 572 316
rect 540 296 544 304
rect 562 296 572 304
rect 540 284 572 296
rect 540 276 544 284
rect 562 276 572 284
rect 540 264 572 276
rect 540 256 544 264
rect 562 256 572 264
rect 540 244 572 256
rect 540 236 544 244
rect 562 236 572 244
rect 540 224 572 236
rect 540 216 544 224
rect 562 216 572 224
rect 540 204 572 216
rect 540 196 544 204
rect 562 196 572 204
rect 540 184 572 196
rect 540 176 544 184
rect 562 176 572 184
rect 540 164 572 176
rect 540 156 544 164
rect 562 156 572 164
rect 540 144 572 156
rect 540 136 544 144
rect 562 136 572 144
rect 540 124 572 136
rect 540 116 544 124
rect 562 116 572 124
rect 540 104 572 116
rect 540 96 544 104
rect 562 96 572 104
rect 540 84 572 96
rect 284 68 291 76
rect 309 68 316 76
rect 284 58 316 68
rect 324 58 524 62
rect 540 76 544 84
rect 562 76 572 84
rect 540 64 572 76
rect 540 58 544 64
rect 56 56 544 58
rect 562 56 572 64
rect 28 54 572 56
rect 28 46 68 54
rect 76 46 88 54
rect 96 46 108 54
rect 116 46 128 54
rect 136 46 148 54
rect 156 46 168 54
rect 176 46 188 54
rect 196 46 404 54
rect 412 46 424 54
rect 432 46 444 54
rect 452 46 464 54
rect 472 46 484 54
rect 492 46 504 54
rect 512 46 524 54
rect 532 46 572 54
rect 28 44 572 46
rect 28 36 38 44
rect 66 36 78 44
rect 86 36 98 44
rect 106 36 118 44
rect 126 36 138 44
rect 146 36 158 44
rect 166 36 178 44
rect 186 36 414 44
rect 422 36 434 44
rect 442 36 454 44
rect 462 36 474 44
rect 482 36 494 44
rect 502 36 514 44
rect 522 36 534 44
rect 562 36 572 44
rect 28 26 572 36
<< nsubstratendiff >>
rect 40 1298 560 1300
rect 40 1290 46 1298
rect 54 1290 66 1298
rect 84 1290 96 1298
rect 114 1290 126 1298
rect 144 1290 156 1298
rect 174 1290 186 1298
rect 204 1290 216 1298
rect 234 1290 246 1298
rect 264 1290 276 1298
rect 294 1290 306 1298
rect 324 1290 336 1298
rect 354 1290 366 1298
rect 384 1290 396 1298
rect 414 1290 426 1298
rect 444 1290 456 1298
rect 474 1290 486 1298
rect 504 1290 516 1298
rect 534 1290 546 1298
rect 554 1290 560 1298
rect 40 1288 76 1290
rect 84 1288 106 1290
rect 114 1288 136 1290
rect 144 1288 166 1290
rect 174 1288 196 1290
rect 204 1288 226 1290
rect 234 1288 256 1290
rect 264 1288 286 1290
rect 294 1288 316 1290
rect 324 1288 346 1290
rect 354 1288 376 1290
rect 384 1288 406 1290
rect 414 1288 436 1290
rect 444 1288 466 1290
rect 474 1288 496 1290
rect 504 1288 526 1290
rect 534 1288 560 1290
rect 40 1280 56 1288
rect 64 1280 76 1288
rect 94 1280 106 1288
rect 124 1280 136 1288
rect 154 1280 166 1288
rect 184 1280 196 1288
rect 214 1280 226 1288
rect 244 1280 256 1288
rect 274 1280 286 1288
rect 304 1280 316 1288
rect 334 1280 346 1288
rect 364 1280 376 1288
rect 394 1280 406 1288
rect 424 1280 436 1288
rect 454 1280 466 1288
rect 484 1280 496 1288
rect 514 1280 526 1288
rect 544 1280 560 1288
rect 40 1278 76 1280
rect 84 1278 106 1280
rect 114 1278 136 1280
rect 144 1278 166 1280
rect 174 1278 196 1280
rect 204 1278 226 1280
rect 234 1278 256 1280
rect 264 1278 286 1280
rect 294 1278 316 1280
rect 324 1278 346 1280
rect 354 1278 376 1280
rect 384 1278 406 1280
rect 414 1278 436 1280
rect 444 1278 466 1280
rect 474 1278 496 1280
rect 504 1278 526 1280
rect 534 1278 560 1280
rect 40 1270 46 1278
rect 54 1270 66 1278
rect 84 1270 96 1278
rect 114 1270 126 1278
rect 144 1270 156 1278
rect 174 1270 186 1278
rect 204 1270 216 1278
rect 234 1270 246 1278
rect 264 1270 276 1278
rect 294 1270 306 1278
rect 324 1270 336 1278
rect 354 1270 366 1278
rect 384 1270 396 1278
rect 414 1270 426 1278
rect 444 1270 456 1278
rect 474 1270 486 1278
rect 504 1270 516 1278
rect 534 1270 546 1278
rect 554 1270 560 1278
rect 40 1268 76 1270
rect 84 1268 106 1270
rect 114 1268 136 1270
rect 144 1268 166 1270
rect 174 1268 196 1270
rect 204 1268 226 1270
rect 234 1268 256 1270
rect 264 1268 286 1270
rect 294 1268 316 1270
rect 324 1268 346 1270
rect 354 1268 376 1270
rect 384 1268 406 1270
rect 414 1268 436 1270
rect 444 1268 466 1270
rect 474 1268 496 1270
rect 504 1268 526 1270
rect 534 1268 560 1270
rect 40 1260 56 1268
rect 64 1260 76 1268
rect 94 1260 106 1268
rect 124 1260 136 1268
rect 154 1260 166 1268
rect 184 1260 196 1268
rect 214 1260 226 1268
rect 244 1260 256 1268
rect 274 1260 286 1268
rect 304 1260 316 1268
rect 334 1260 346 1268
rect 364 1260 376 1268
rect 394 1260 406 1268
rect 424 1260 436 1268
rect 454 1260 466 1268
rect 484 1260 496 1268
rect 514 1260 526 1268
rect 544 1260 560 1268
rect 40 1258 76 1260
rect 84 1258 106 1260
rect 114 1258 136 1260
rect 144 1258 166 1260
rect 174 1258 196 1260
rect 204 1258 226 1260
rect 234 1258 256 1260
rect 264 1258 286 1260
rect 294 1258 316 1260
rect 324 1258 346 1260
rect 354 1258 376 1260
rect 384 1258 406 1260
rect 414 1258 436 1260
rect 444 1258 466 1260
rect 474 1258 496 1260
rect 504 1258 526 1260
rect 534 1258 560 1260
rect 40 1250 46 1258
rect 54 1250 66 1258
rect 84 1250 96 1258
rect 114 1250 126 1258
rect 144 1250 156 1258
rect 174 1250 186 1258
rect 204 1250 216 1258
rect 234 1250 246 1258
rect 264 1250 276 1258
rect 294 1250 306 1258
rect 324 1250 336 1258
rect 354 1250 366 1258
rect 384 1250 396 1258
rect 414 1250 426 1258
rect 444 1250 456 1258
rect 474 1250 486 1258
rect 504 1250 516 1258
rect 534 1250 546 1258
rect 554 1250 560 1258
rect 40 1248 76 1250
rect 84 1248 106 1250
rect 114 1248 136 1250
rect 144 1248 166 1250
rect 174 1248 196 1250
rect 204 1248 226 1250
rect 234 1248 256 1250
rect 264 1248 286 1250
rect 294 1248 316 1250
rect 324 1248 346 1250
rect 354 1248 376 1250
rect 384 1248 406 1250
rect 414 1248 436 1250
rect 444 1248 466 1250
rect 474 1248 496 1250
rect 504 1248 526 1250
rect 534 1248 560 1250
rect 40 1240 56 1248
rect 64 1240 76 1248
rect 94 1240 106 1248
rect 124 1240 136 1248
rect 154 1240 166 1248
rect 184 1240 196 1248
rect 214 1240 226 1248
rect 244 1240 256 1248
rect 274 1240 286 1248
rect 304 1240 316 1248
rect 334 1240 346 1248
rect 364 1240 376 1248
rect 394 1240 406 1248
rect 424 1240 436 1248
rect 454 1240 466 1248
rect 484 1240 496 1248
rect 514 1240 526 1248
rect 544 1240 560 1248
rect 40 1238 76 1240
rect 84 1238 106 1240
rect 114 1238 136 1240
rect 144 1238 166 1240
rect 174 1238 196 1240
rect 204 1238 226 1240
rect 234 1238 256 1240
rect 264 1238 286 1240
rect 294 1238 316 1240
rect 324 1238 346 1240
rect 354 1238 376 1240
rect 384 1238 406 1240
rect 414 1238 436 1240
rect 444 1238 466 1240
rect 474 1238 496 1240
rect 504 1238 526 1240
rect 534 1238 560 1240
rect 40 1230 46 1238
rect 54 1230 66 1238
rect 84 1230 96 1238
rect 114 1230 126 1238
rect 144 1230 156 1238
rect 174 1230 186 1238
rect 204 1230 216 1238
rect 234 1230 246 1238
rect 264 1230 276 1238
rect 294 1230 306 1238
rect 324 1230 336 1238
rect 354 1230 366 1238
rect 384 1230 396 1238
rect 414 1230 426 1238
rect 444 1230 456 1238
rect 474 1230 486 1238
rect 504 1230 516 1238
rect 534 1230 546 1238
rect 554 1230 560 1238
rect 40 1228 76 1230
rect 84 1228 106 1230
rect 114 1228 136 1230
rect 144 1228 166 1230
rect 174 1228 196 1230
rect 204 1228 226 1230
rect 234 1228 256 1230
rect 264 1228 286 1230
rect 294 1228 316 1230
rect 324 1228 346 1230
rect 354 1228 376 1230
rect 384 1228 406 1230
rect 414 1228 436 1230
rect 444 1228 466 1230
rect 474 1228 496 1230
rect 504 1228 526 1230
rect 534 1228 560 1230
rect 40 1220 56 1228
rect 64 1220 76 1228
rect 94 1220 106 1228
rect 124 1220 136 1228
rect 154 1220 166 1228
rect 184 1220 196 1228
rect 214 1220 226 1228
rect 244 1220 256 1228
rect 274 1220 286 1228
rect 304 1220 316 1228
rect 334 1220 346 1228
rect 364 1220 376 1228
rect 394 1220 406 1228
rect 424 1220 436 1228
rect 454 1220 466 1228
rect 484 1220 496 1228
rect 514 1220 526 1228
rect 544 1220 560 1228
rect 40 1218 76 1220
rect 84 1218 106 1220
rect 114 1218 136 1220
rect 144 1218 166 1220
rect 174 1218 196 1220
rect 204 1218 226 1220
rect 234 1218 256 1220
rect 264 1218 286 1220
rect 294 1218 316 1220
rect 324 1218 346 1220
rect 354 1218 376 1220
rect 384 1218 406 1220
rect 414 1218 436 1220
rect 444 1218 466 1220
rect 474 1218 496 1220
rect 504 1218 526 1220
rect 534 1218 560 1220
rect 40 1210 46 1218
rect 54 1210 66 1218
rect 84 1210 96 1218
rect 114 1210 126 1218
rect 144 1210 156 1218
rect 174 1210 186 1218
rect 204 1210 216 1218
rect 234 1210 246 1218
rect 264 1210 276 1218
rect 294 1210 306 1218
rect 324 1210 336 1218
rect 354 1210 366 1218
rect 384 1210 396 1218
rect 414 1210 426 1218
rect 444 1210 456 1218
rect 474 1210 486 1218
rect 504 1210 516 1218
rect 534 1210 546 1218
rect 554 1210 560 1218
rect 40 1208 76 1210
rect 84 1208 106 1210
rect 114 1208 136 1210
rect 144 1208 166 1210
rect 174 1208 196 1210
rect 204 1208 226 1210
rect 234 1208 256 1210
rect 264 1208 286 1210
rect 294 1208 316 1210
rect 324 1208 346 1210
rect 354 1208 376 1210
rect 384 1208 406 1210
rect 414 1208 436 1210
rect 444 1208 466 1210
rect 474 1208 496 1210
rect 504 1208 526 1210
rect 534 1208 560 1210
rect 40 1200 56 1208
rect 64 1200 76 1208
rect 94 1200 106 1208
rect 124 1200 136 1208
rect 154 1200 166 1208
rect 184 1200 196 1208
rect 214 1200 226 1208
rect 244 1200 256 1208
rect 274 1200 286 1208
rect 304 1200 316 1208
rect 334 1200 346 1208
rect 364 1200 376 1208
rect 394 1200 406 1208
rect 424 1200 436 1208
rect 454 1200 466 1208
rect 484 1200 496 1208
rect 514 1200 526 1208
rect 544 1200 560 1208
rect 40 1198 76 1200
rect 84 1198 106 1200
rect 114 1198 136 1200
rect 144 1198 166 1200
rect 174 1198 196 1200
rect 204 1198 226 1200
rect 234 1198 256 1200
rect 264 1198 286 1200
rect 294 1198 316 1200
rect 324 1198 346 1200
rect 354 1198 376 1200
rect 384 1198 406 1200
rect 414 1198 436 1200
rect 444 1198 466 1200
rect 474 1198 496 1200
rect 504 1198 526 1200
rect 534 1198 560 1200
rect 40 1190 46 1198
rect 54 1190 66 1198
rect 84 1190 96 1198
rect 114 1190 126 1198
rect 144 1190 156 1198
rect 174 1190 186 1198
rect 204 1190 216 1198
rect 234 1190 246 1198
rect 264 1190 276 1198
rect 294 1190 306 1198
rect 324 1190 336 1198
rect 354 1190 366 1198
rect 384 1190 396 1198
rect 414 1190 426 1198
rect 444 1190 456 1198
rect 474 1190 486 1198
rect 504 1190 516 1198
rect 534 1190 546 1198
rect 554 1190 560 1198
rect 40 1188 76 1190
rect 84 1188 526 1190
rect 534 1188 560 1190
rect 40 1180 56 1188
rect 64 1180 76 1188
rect 94 1180 506 1188
rect 514 1180 526 1188
rect 544 1180 560 1188
rect 40 1178 76 1180
rect 84 1178 526 1180
rect 534 1178 560 1180
rect 40 1170 46 1178
rect 54 1170 66 1178
rect 84 1170 96 1178
rect 114 1170 126 1178
rect 144 1170 156 1178
rect 174 1170 186 1178
rect 204 1170 216 1178
rect 234 1170 246 1178
rect 264 1170 276 1178
rect 294 1170 306 1178
rect 324 1170 336 1178
rect 354 1170 366 1178
rect 384 1170 396 1178
rect 414 1170 426 1178
rect 444 1170 456 1178
rect 474 1170 486 1178
rect 504 1170 516 1178
rect 534 1170 546 1178
rect 554 1170 560 1178
rect 40 1168 76 1170
rect 84 1168 106 1170
rect 114 1168 136 1170
rect 144 1168 166 1170
rect 174 1168 196 1170
rect 204 1168 226 1170
rect 234 1168 256 1170
rect 264 1168 286 1170
rect 294 1168 316 1170
rect 324 1168 346 1170
rect 354 1168 376 1170
rect 384 1168 406 1170
rect 414 1168 436 1170
rect 444 1168 466 1170
rect 474 1168 496 1170
rect 504 1168 526 1170
rect 534 1168 560 1170
rect 40 1160 56 1168
rect 64 1160 76 1168
rect 94 1160 106 1168
rect 124 1160 136 1168
rect 154 1160 166 1168
rect 184 1160 196 1168
rect 214 1160 226 1168
rect 244 1160 256 1168
rect 274 1160 286 1168
rect 304 1160 316 1168
rect 334 1160 346 1168
rect 364 1160 376 1168
rect 394 1160 406 1168
rect 424 1160 436 1168
rect 454 1160 466 1168
rect 484 1160 496 1168
rect 514 1160 526 1168
rect 544 1160 560 1168
rect 40 1158 76 1160
rect 84 1158 106 1160
rect 114 1158 136 1160
rect 144 1158 166 1160
rect 174 1158 196 1160
rect 204 1158 226 1160
rect 234 1158 256 1160
rect 264 1158 286 1160
rect 294 1158 316 1160
rect 324 1158 346 1160
rect 354 1158 376 1160
rect 384 1158 406 1160
rect 414 1158 436 1160
rect 444 1158 466 1160
rect 474 1158 496 1160
rect 504 1158 526 1160
rect 534 1158 560 1160
rect 40 1150 46 1158
rect 54 1150 66 1158
rect 84 1150 96 1158
rect 114 1150 126 1158
rect 144 1150 156 1158
rect 174 1150 186 1158
rect 204 1150 216 1158
rect 234 1150 246 1158
rect 264 1150 276 1158
rect 294 1150 306 1158
rect 324 1150 336 1158
rect 354 1150 366 1158
rect 384 1150 396 1158
rect 414 1150 426 1158
rect 444 1150 456 1158
rect 474 1150 486 1158
rect 504 1150 516 1158
rect 534 1150 546 1158
rect 554 1150 560 1158
rect 40 1148 76 1150
rect 84 1148 106 1150
rect 114 1148 136 1150
rect 144 1148 166 1150
rect 174 1148 196 1150
rect 204 1148 226 1150
rect 234 1148 256 1150
rect 264 1148 286 1150
rect 294 1148 316 1150
rect 324 1148 346 1150
rect 354 1148 376 1150
rect 384 1148 406 1150
rect 414 1148 436 1150
rect 444 1148 466 1150
rect 474 1148 496 1150
rect 504 1148 526 1150
rect 534 1148 560 1150
rect 40 1140 56 1148
rect 64 1140 76 1148
rect 94 1140 106 1148
rect 124 1140 136 1148
rect 154 1140 166 1148
rect 184 1140 196 1148
rect 214 1140 226 1148
rect 244 1140 256 1148
rect 274 1140 286 1148
rect 304 1140 316 1148
rect 334 1140 346 1148
rect 364 1140 376 1148
rect 394 1140 406 1148
rect 424 1140 436 1148
rect 454 1140 466 1148
rect 484 1140 496 1148
rect 514 1140 526 1148
rect 544 1140 560 1148
rect 40 1138 76 1140
rect 84 1138 106 1140
rect 114 1138 136 1140
rect 144 1138 166 1140
rect 174 1138 196 1140
rect 204 1138 226 1140
rect 234 1138 256 1140
rect 264 1138 286 1140
rect 294 1138 316 1140
rect 324 1138 346 1140
rect 354 1138 376 1140
rect 384 1138 406 1140
rect 414 1138 436 1140
rect 444 1138 466 1140
rect 474 1138 496 1140
rect 504 1138 526 1140
rect 534 1138 560 1140
rect 40 1130 46 1138
rect 54 1130 66 1138
rect 84 1130 96 1138
rect 114 1130 126 1138
rect 144 1130 156 1138
rect 174 1130 186 1138
rect 204 1130 216 1138
rect 234 1130 246 1138
rect 264 1130 276 1138
rect 294 1130 306 1138
rect 324 1130 336 1138
rect 354 1130 366 1138
rect 384 1130 396 1138
rect 414 1130 426 1138
rect 444 1130 456 1138
rect 474 1130 486 1138
rect 504 1130 516 1138
rect 534 1130 546 1138
rect 554 1130 560 1138
rect 40 1128 76 1130
rect 84 1128 106 1130
rect 114 1128 136 1130
rect 144 1128 166 1130
rect 174 1128 196 1130
rect 204 1128 226 1130
rect 234 1128 256 1130
rect 264 1128 286 1130
rect 294 1128 316 1130
rect 324 1128 346 1130
rect 354 1128 376 1130
rect 384 1128 406 1130
rect 414 1128 436 1130
rect 444 1128 466 1130
rect 474 1128 496 1130
rect 504 1128 526 1130
rect 534 1128 560 1130
rect 40 1120 56 1128
rect 64 1120 76 1128
rect 94 1120 106 1128
rect 124 1120 136 1128
rect 154 1120 166 1128
rect 184 1120 196 1128
rect 214 1120 226 1128
rect 244 1120 256 1128
rect 274 1120 286 1128
rect 304 1120 316 1128
rect 334 1120 346 1128
rect 364 1120 376 1128
rect 394 1120 406 1128
rect 424 1120 436 1128
rect 454 1120 466 1128
rect 484 1120 496 1128
rect 40 1118 86 1120
rect 40 1110 46 1118
rect 54 1110 66 1118
rect 74 1110 86 1118
rect 40 1108 86 1110
rect 94 1108 506 1120
rect 40 1100 56 1108
rect 64 1100 76 1108
rect 94 1100 106 1108
rect 124 1100 136 1108
rect 154 1100 166 1108
rect 184 1100 196 1108
rect 214 1100 226 1108
rect 244 1100 256 1108
rect 274 1100 286 1108
rect 304 1100 316 1108
rect 334 1100 346 1108
rect 364 1100 376 1108
rect 394 1100 406 1108
rect 424 1100 436 1108
rect 454 1100 466 1108
rect 484 1100 496 1108
rect 514 1100 526 1128
rect 544 1120 560 1128
rect 534 1118 560 1120
rect 534 1110 546 1118
rect 554 1110 560 1118
rect 534 1108 560 1110
rect 544 1100 560 1108
rect 40 1098 76 1100
rect 84 1098 106 1100
rect 114 1098 136 1100
rect 144 1098 166 1100
rect 174 1098 196 1100
rect 204 1098 226 1100
rect 234 1098 256 1100
rect 264 1098 286 1100
rect 294 1098 316 1100
rect 324 1098 346 1100
rect 354 1098 376 1100
rect 384 1098 406 1100
rect 414 1098 436 1100
rect 444 1098 466 1100
rect 474 1098 496 1100
rect 504 1098 526 1100
rect 534 1098 560 1100
rect 40 1090 46 1098
rect 54 1090 66 1098
rect 84 1090 96 1098
rect 114 1090 126 1098
rect 144 1090 156 1098
rect 174 1090 186 1098
rect 204 1090 216 1098
rect 234 1090 246 1098
rect 264 1090 276 1098
rect 294 1090 306 1098
rect 324 1090 336 1098
rect 354 1090 366 1098
rect 384 1090 396 1098
rect 414 1090 426 1098
rect 444 1090 456 1098
rect 474 1090 486 1098
rect 504 1090 516 1098
rect 534 1090 546 1098
rect 554 1090 560 1098
rect 40 1088 76 1090
rect 84 1088 106 1090
rect 114 1088 136 1090
rect 144 1088 166 1090
rect 174 1088 196 1090
rect 204 1088 226 1090
rect 234 1088 256 1090
rect 264 1088 286 1090
rect 294 1088 316 1090
rect 324 1088 346 1090
rect 354 1088 376 1090
rect 384 1088 406 1090
rect 414 1088 436 1090
rect 444 1088 466 1090
rect 474 1088 496 1090
rect 504 1088 526 1090
rect 534 1088 560 1090
rect 40 1080 56 1088
rect 64 1080 76 1088
rect 94 1080 106 1088
rect 124 1080 136 1088
rect 154 1080 166 1088
rect 184 1080 196 1088
rect 214 1080 226 1088
rect 244 1080 256 1088
rect 274 1080 286 1088
rect 304 1080 316 1088
rect 334 1080 346 1088
rect 364 1080 376 1088
rect 394 1080 406 1088
rect 424 1080 436 1088
rect 454 1080 466 1088
rect 484 1080 496 1088
rect 514 1080 526 1088
rect 544 1080 560 1088
rect 40 1078 76 1080
rect 84 1078 106 1080
rect 114 1078 136 1080
rect 144 1078 166 1080
rect 174 1078 196 1080
rect 204 1078 226 1080
rect 234 1078 256 1080
rect 264 1078 286 1080
rect 294 1078 316 1080
rect 324 1078 346 1080
rect 354 1078 376 1080
rect 384 1078 406 1080
rect 414 1078 436 1080
rect 444 1078 466 1080
rect 474 1078 496 1080
rect 504 1078 526 1080
rect 534 1078 560 1080
rect 40 1070 46 1078
rect 54 1070 66 1078
rect 84 1070 96 1078
rect 114 1070 126 1078
rect 144 1070 156 1078
rect 174 1070 186 1078
rect 204 1070 216 1078
rect 234 1070 246 1078
rect 264 1070 276 1078
rect 294 1070 306 1078
rect 324 1070 336 1078
rect 354 1070 366 1078
rect 384 1070 396 1078
rect 414 1070 426 1078
rect 444 1070 456 1078
rect 474 1070 486 1078
rect 504 1070 516 1078
rect 534 1070 546 1078
rect 554 1070 560 1078
rect 40 1068 76 1070
rect 84 1068 106 1070
rect 114 1068 136 1070
rect 144 1068 166 1070
rect 174 1068 196 1070
rect 204 1068 226 1070
rect 234 1068 256 1070
rect 264 1068 286 1070
rect 294 1068 316 1070
rect 324 1068 346 1070
rect 354 1068 376 1070
rect 384 1068 406 1070
rect 414 1068 436 1070
rect 444 1068 466 1070
rect 474 1068 496 1070
rect 504 1068 526 1070
rect 534 1068 560 1070
rect 40 1060 56 1068
rect 64 1060 76 1068
rect 94 1060 106 1068
rect 124 1060 136 1068
rect 154 1060 166 1068
rect 184 1060 196 1068
rect 214 1060 226 1068
rect 244 1060 256 1068
rect 274 1060 286 1068
rect 304 1060 316 1068
rect 334 1060 346 1068
rect 364 1060 376 1068
rect 394 1060 406 1068
rect 424 1060 436 1068
rect 454 1060 466 1068
rect 484 1060 496 1068
rect 514 1060 526 1068
rect 544 1060 560 1068
rect 40 1058 76 1060
rect 84 1058 106 1060
rect 114 1058 136 1060
rect 144 1058 166 1060
rect 174 1058 196 1060
rect 204 1058 226 1060
rect 234 1058 256 1060
rect 264 1058 286 1060
rect 294 1058 316 1060
rect 324 1058 346 1060
rect 354 1058 376 1060
rect 384 1058 406 1060
rect 414 1058 436 1060
rect 444 1058 466 1060
rect 474 1058 496 1060
rect 504 1058 526 1060
rect 534 1058 560 1060
rect 40 1050 46 1058
rect 54 1050 66 1058
rect 84 1050 96 1058
rect 114 1050 126 1058
rect 144 1050 156 1058
rect 174 1050 186 1058
rect 204 1050 216 1058
rect 234 1050 246 1058
rect 264 1050 276 1058
rect 294 1050 306 1058
rect 324 1050 336 1058
rect 354 1050 366 1058
rect 384 1050 396 1058
rect 414 1050 426 1058
rect 444 1050 456 1058
rect 474 1050 486 1058
rect 504 1050 516 1058
rect 534 1050 546 1058
rect 554 1050 560 1058
rect 40 1048 76 1050
rect 84 1048 106 1050
rect 114 1048 136 1050
rect 144 1048 166 1050
rect 174 1048 196 1050
rect 204 1048 226 1050
rect 234 1048 256 1050
rect 264 1048 286 1050
rect 294 1048 316 1050
rect 324 1048 346 1050
rect 354 1048 376 1050
rect 384 1048 406 1050
rect 414 1048 436 1050
rect 444 1048 466 1050
rect 474 1048 496 1050
rect 504 1048 526 1050
rect 534 1048 560 1050
rect 40 1040 56 1048
rect 64 1040 76 1048
rect 94 1040 106 1048
rect 124 1040 136 1048
rect 154 1040 166 1048
rect 184 1040 196 1048
rect 214 1040 226 1048
rect 244 1040 256 1048
rect 274 1040 286 1048
rect 304 1040 316 1048
rect 334 1040 346 1048
rect 364 1040 376 1048
rect 394 1040 406 1048
rect 424 1040 436 1048
rect 454 1040 466 1048
rect 484 1040 496 1048
rect 40 1038 76 1040
rect 40 1030 46 1038
rect 54 1030 66 1038
rect 40 1028 76 1030
rect 84 1028 506 1040
rect 40 1020 56 1028
rect 64 1020 76 1028
rect 94 1020 106 1028
rect 124 1020 136 1028
rect 154 1020 166 1028
rect 184 1020 196 1028
rect 214 1020 226 1028
rect 244 1020 256 1028
rect 274 1020 286 1028
rect 304 1020 316 1028
rect 334 1020 346 1028
rect 364 1020 376 1028
rect 394 1020 406 1028
rect 424 1020 436 1028
rect 454 1020 466 1028
rect 484 1020 496 1028
rect 514 1020 526 1048
rect 544 1040 560 1048
rect 534 1038 560 1040
rect 534 1030 546 1038
rect 554 1030 560 1038
rect 534 1028 560 1030
rect 544 1020 560 1028
rect 40 1018 76 1020
rect 84 1018 106 1020
rect 114 1018 136 1020
rect 144 1018 166 1020
rect 174 1018 196 1020
rect 204 1018 226 1020
rect 234 1018 256 1020
rect 264 1018 286 1020
rect 294 1018 316 1020
rect 324 1018 346 1020
rect 354 1018 376 1020
rect 384 1018 406 1020
rect 414 1018 436 1020
rect 444 1018 466 1020
rect 474 1018 496 1020
rect 504 1018 526 1020
rect 534 1018 560 1020
rect 40 1010 46 1018
rect 54 1010 66 1018
rect 84 1010 96 1018
rect 114 1010 126 1018
rect 144 1010 156 1018
rect 174 1010 186 1018
rect 204 1010 216 1018
rect 234 1010 246 1018
rect 264 1010 276 1018
rect 294 1010 306 1018
rect 324 1010 336 1018
rect 354 1010 366 1018
rect 384 1010 396 1018
rect 414 1010 426 1018
rect 444 1010 456 1018
rect 474 1010 486 1018
rect 504 1010 516 1018
rect 534 1010 546 1018
rect 554 1010 560 1018
rect 40 1008 76 1010
rect 84 1008 106 1010
rect 114 1008 136 1010
rect 144 1008 166 1010
rect 174 1008 196 1010
rect 204 1008 226 1010
rect 234 1008 256 1010
rect 264 1008 286 1010
rect 294 1008 316 1010
rect 324 1008 346 1010
rect 354 1008 376 1010
rect 384 1008 406 1010
rect 414 1008 436 1010
rect 444 1008 466 1010
rect 474 1008 496 1010
rect 504 1008 526 1010
rect 534 1008 560 1010
rect 40 1000 56 1008
rect 64 1000 76 1008
rect 94 1000 106 1008
rect 124 1000 136 1008
rect 154 1000 166 1008
rect 184 1000 196 1008
rect 214 1000 226 1008
rect 244 1000 256 1008
rect 274 1000 286 1008
rect 304 1000 316 1008
rect 334 1000 346 1008
rect 364 1000 376 1008
rect 394 1000 406 1008
rect 424 1000 436 1008
rect 454 1000 466 1008
rect 484 1000 496 1008
rect 514 1000 526 1008
rect 544 1000 560 1008
rect 40 998 76 1000
rect 84 998 106 1000
rect 114 998 136 1000
rect 144 998 166 1000
rect 174 998 196 1000
rect 204 998 226 1000
rect 234 998 256 1000
rect 264 998 286 1000
rect 294 998 316 1000
rect 324 998 346 1000
rect 354 998 376 1000
rect 384 998 406 1000
rect 414 998 436 1000
rect 444 998 466 1000
rect 474 998 496 1000
rect 504 998 526 1000
rect 534 998 560 1000
rect 40 990 46 998
rect 54 990 66 998
rect 84 990 96 998
rect 114 990 126 998
rect 144 990 156 998
rect 174 990 186 998
rect 204 990 216 998
rect 234 990 246 998
rect 264 990 276 998
rect 294 990 306 998
rect 324 990 336 998
rect 354 990 366 998
rect 384 990 396 998
rect 414 990 426 998
rect 444 990 456 998
rect 474 990 486 998
rect 504 990 516 998
rect 534 990 546 998
rect 554 990 560 998
rect 40 988 76 990
rect 84 988 106 990
rect 114 988 136 990
rect 144 988 166 990
rect 174 988 196 990
rect 204 988 226 990
rect 234 988 256 990
rect 264 988 286 990
rect 294 988 316 990
rect 324 988 346 990
rect 354 988 376 990
rect 384 988 406 990
rect 414 988 436 990
rect 444 988 466 990
rect 474 988 496 990
rect 504 988 526 990
rect 534 988 560 990
rect 40 980 56 988
rect 64 980 76 988
rect 94 980 106 988
rect 124 980 136 988
rect 154 980 166 988
rect 184 980 196 988
rect 214 980 226 988
rect 244 980 256 988
rect 274 980 286 988
rect 304 980 316 988
rect 334 980 346 988
rect 364 980 376 988
rect 394 980 406 988
rect 424 980 436 988
rect 454 980 466 988
rect 484 980 496 988
rect 514 980 526 988
rect 544 980 560 988
rect 40 978 76 980
rect 84 978 106 980
rect 114 978 136 980
rect 144 978 166 980
rect 174 978 196 980
rect 204 978 226 980
rect 234 978 256 980
rect 264 978 286 980
rect 294 978 316 980
rect 324 978 346 980
rect 354 978 376 980
rect 384 978 406 980
rect 414 978 436 980
rect 444 978 466 980
rect 474 978 496 980
rect 504 978 526 980
rect 534 978 560 980
rect 40 970 46 978
rect 54 970 66 978
rect 84 970 96 978
rect 114 970 126 978
rect 144 970 156 978
rect 174 970 186 978
rect 204 970 216 978
rect 234 970 246 978
rect 264 970 276 978
rect 294 970 306 978
rect 324 970 336 978
rect 354 970 366 978
rect 384 970 396 978
rect 414 970 426 978
rect 444 970 456 978
rect 474 970 486 978
rect 504 970 516 978
rect 534 970 546 978
rect 554 970 560 978
rect 40 968 560 970
rect 40 960 536 968
rect 544 960 560 968
rect 40 958 560 960
rect 40 950 46 958
rect 54 950 66 958
rect 84 950 96 958
rect 114 950 126 958
rect 144 950 156 958
rect 174 950 186 958
rect 204 950 216 958
rect 234 950 246 958
rect 264 950 276 958
rect 294 950 306 958
rect 324 950 336 958
rect 354 950 366 958
rect 384 950 396 958
rect 414 950 426 958
rect 444 950 456 958
rect 474 950 486 958
rect 504 950 516 958
rect 534 950 546 958
rect 554 950 560 958
rect 40 948 76 950
rect 84 948 106 950
rect 114 948 136 950
rect 144 948 166 950
rect 174 948 196 950
rect 204 948 226 950
rect 234 948 256 950
rect 264 948 286 950
rect 294 948 316 950
rect 324 948 346 950
rect 354 948 376 950
rect 384 948 406 950
rect 414 948 436 950
rect 444 948 466 950
rect 474 948 496 950
rect 504 948 526 950
rect 534 948 560 950
rect 40 940 56 948
rect 64 940 76 948
rect 94 940 106 948
rect 124 940 136 948
rect 154 940 166 948
rect 184 940 196 948
rect 214 940 226 948
rect 244 940 256 948
rect 274 940 286 948
rect 304 940 316 948
rect 334 940 346 948
rect 364 940 376 948
rect 394 940 406 948
rect 424 940 436 948
rect 454 940 466 948
rect 484 940 496 948
rect 514 940 526 948
rect 544 940 560 948
rect 40 938 76 940
rect 84 938 106 940
rect 114 938 136 940
rect 144 938 166 940
rect 174 938 196 940
rect 204 938 226 940
rect 234 938 256 940
rect 264 938 286 940
rect 294 938 316 940
rect 324 938 346 940
rect 354 938 376 940
rect 384 938 406 940
rect 414 938 436 940
rect 444 938 466 940
rect 474 938 496 940
rect 504 938 526 940
rect 534 938 560 940
rect 40 930 46 938
rect 54 930 66 938
rect 84 930 96 938
rect 114 930 126 938
rect 144 930 156 938
rect 174 930 186 938
rect 204 930 216 938
rect 234 930 246 938
rect 264 930 276 938
rect 294 930 306 938
rect 324 930 336 938
rect 354 930 366 938
rect 384 930 396 938
rect 414 930 426 938
rect 444 930 456 938
rect 474 930 486 938
rect 504 930 516 938
rect 534 930 546 938
rect 554 930 560 938
rect 40 928 76 930
rect 84 928 106 930
rect 114 928 136 930
rect 144 928 166 930
rect 174 928 196 930
rect 204 928 226 930
rect 234 928 256 930
rect 264 928 286 930
rect 294 928 316 930
rect 324 928 346 930
rect 354 928 376 930
rect 384 928 406 930
rect 414 928 436 930
rect 444 928 466 930
rect 474 928 496 930
rect 504 928 526 930
rect 534 928 560 930
rect 40 920 56 928
rect 64 920 76 928
rect 94 920 106 928
rect 124 920 136 928
rect 154 920 166 928
rect 184 920 196 928
rect 214 920 226 928
rect 244 920 256 928
rect 274 920 286 928
rect 304 920 316 928
rect 334 920 346 928
rect 364 920 376 928
rect 394 920 406 928
rect 424 920 436 928
rect 454 920 466 928
rect 484 920 496 928
rect 514 920 526 928
rect 544 920 560 928
rect 40 918 76 920
rect 84 918 106 920
rect 114 918 136 920
rect 144 918 166 920
rect 174 918 196 920
rect 204 918 226 920
rect 234 918 256 920
rect 264 918 286 920
rect 294 918 316 920
rect 324 918 346 920
rect 354 918 376 920
rect 384 918 406 920
rect 414 918 436 920
rect 444 918 466 920
rect 474 918 496 920
rect 504 918 526 920
rect 534 918 560 920
rect 40 910 46 918
rect 54 910 66 918
rect 84 910 96 918
rect 114 910 126 918
rect 144 910 156 918
rect 174 910 186 918
rect 204 910 216 918
rect 234 910 246 918
rect 264 910 276 918
rect 294 910 306 918
rect 324 910 336 918
rect 354 910 366 918
rect 384 910 396 918
rect 414 910 426 918
rect 444 910 456 918
rect 474 910 486 918
rect 504 910 516 918
rect 534 910 546 918
rect 554 910 560 918
rect 40 908 76 910
rect 84 908 106 910
rect 114 908 136 910
rect 144 908 166 910
rect 174 908 196 910
rect 204 908 226 910
rect 234 908 256 910
rect 264 908 286 910
rect 294 908 316 910
rect 324 908 346 910
rect 354 908 376 910
rect 384 908 406 910
rect 414 908 436 910
rect 444 908 466 910
rect 474 908 496 910
rect 504 908 526 910
rect 534 908 560 910
rect 40 900 56 908
rect 64 900 76 908
rect 94 900 106 908
rect 124 900 136 908
rect 154 900 166 908
rect 184 900 196 908
rect 214 900 226 908
rect 244 900 256 908
rect 274 900 286 908
rect 304 900 316 908
rect 334 900 346 908
rect 364 900 376 908
rect 394 900 406 908
rect 424 900 436 908
rect 454 900 466 908
rect 484 900 496 908
rect 514 900 526 908
rect 544 900 560 908
rect 40 898 76 900
rect 84 898 106 900
rect 114 898 136 900
rect 144 898 166 900
rect 174 898 196 900
rect 204 898 226 900
rect 234 898 256 900
rect 264 898 286 900
rect 294 898 316 900
rect 324 898 346 900
rect 354 898 376 900
rect 384 898 406 900
rect 414 898 436 900
rect 444 898 466 900
rect 474 898 496 900
rect 504 898 526 900
rect 534 898 560 900
rect 40 890 46 898
rect 54 890 66 898
rect 84 890 96 898
rect 114 890 126 898
rect 144 890 156 898
rect 174 890 186 898
rect 204 890 216 898
rect 234 890 246 898
rect 264 890 276 898
rect 294 890 306 898
rect 324 890 336 898
rect 354 890 366 898
rect 384 890 396 898
rect 414 890 426 898
rect 444 890 456 898
rect 474 890 486 898
rect 504 890 516 898
rect 534 890 546 898
rect 554 890 560 898
rect 40 888 76 890
rect 84 888 106 890
rect 114 888 136 890
rect 144 888 166 890
rect 174 888 196 890
rect 204 888 226 890
rect 234 888 256 890
rect 264 888 286 890
rect 294 888 316 890
rect 324 888 346 890
rect 354 888 376 890
rect 384 888 406 890
rect 414 888 436 890
rect 444 888 466 890
rect 474 888 496 890
rect 504 888 526 890
rect 534 888 560 890
rect 40 878 56 888
rect 64 878 76 888
rect 94 878 106 888
rect 124 878 136 888
rect 154 878 166 888
rect 184 878 196 888
rect 214 878 226 888
rect 244 878 256 888
rect 274 878 286 888
rect 304 878 316 888
rect 334 878 346 888
rect 364 878 376 888
rect 394 878 406 888
rect 424 878 436 888
rect 454 878 466 888
rect 484 878 496 888
rect 514 878 526 888
rect 544 878 560 888
rect 40 870 46 878
rect 554 870 560 878
rect 40 864 560 870
rect 0 652 600 654
rect 0 644 4 652
rect 12 644 24 652
rect 42 644 54 652
rect 72 644 84 652
rect 102 644 114 652
rect 132 644 144 652
rect 162 644 174 652
rect 192 644 204 652
rect 222 644 234 652
rect 242 644 256 652
rect 264 644 276 652
rect 294 644 306 652
rect 324 644 336 652
rect 344 644 358 652
rect 366 644 378 652
rect 396 644 408 652
rect 426 644 438 652
rect 456 644 468 652
rect 486 644 498 652
rect 516 644 528 652
rect 546 644 558 652
rect 576 644 588 652
rect 596 644 600 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 192 642 214 644
rect 222 642 286 644
rect 294 642 316 644
rect 324 642 378 644
rect 386 642 408 644
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 0 634 14 642
rect 22 634 34 642
rect 52 634 64 642
rect 82 634 94 642
rect 112 634 124 642
rect 142 634 154 642
rect 172 634 184 642
rect 202 634 214 642
rect 232 634 244 642
rect 252 634 266 642
rect 274 634 286 642
rect 304 634 316 642
rect 334 634 348 642
rect 356 634 368 642
rect 386 634 398 642
rect 416 634 428 642
rect 446 634 458 642
rect 476 634 488 642
rect 506 634 518 642
rect 536 634 548 642
rect 566 634 578 642
rect 586 634 600 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 192 632 214 634
rect 222 632 286 634
rect 294 632 316 634
rect 324 632 378 634
rect 386 632 408 634
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 0 624 4 632
rect 12 624 24 632
rect 42 624 54 632
rect 72 624 84 632
rect 102 624 114 632
rect 132 624 144 632
rect 162 624 174 632
rect 192 624 204 632
rect 222 624 234 632
rect 242 624 256 632
rect 264 624 276 632
rect 294 624 306 632
rect 324 624 336 632
rect 344 624 358 632
rect 366 624 378 632
rect 396 624 408 632
rect 426 624 438 632
rect 456 624 468 632
rect 486 624 498 632
rect 516 624 528 632
rect 546 624 558 632
rect 576 624 588 632
rect 596 624 600 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 192 622 214 624
rect 222 622 286 624
rect 294 622 316 624
rect 324 622 378 624
rect 386 622 408 624
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 0 614 14 622
rect 22 614 34 622
rect 52 614 64 622
rect 82 614 94 622
rect 112 614 124 622
rect 142 614 154 622
rect 172 614 184 622
rect 202 614 214 622
rect 232 614 244 622
rect 252 614 266 622
rect 274 614 286 622
rect 304 614 316 622
rect 334 614 348 622
rect 356 614 368 622
rect 386 614 398 622
rect 416 614 428 622
rect 446 614 458 622
rect 476 614 488 622
rect 506 614 518 622
rect 536 614 548 622
rect 566 614 578 622
rect 586 614 600 622
rect 0 612 214 614
rect 0 604 4 612
rect 12 604 24 612
rect 32 604 214 612
rect 0 602 214 604
rect 222 612 286 614
rect 294 612 316 614
rect 324 612 378 614
rect 222 604 234 612
rect 242 604 256 612
rect 264 604 276 612
rect 294 604 306 612
rect 324 604 336 612
rect 344 604 358 612
rect 366 604 378 612
rect 222 602 286 604
rect 294 602 316 604
rect 324 602 378 604
rect 386 612 600 614
rect 386 604 568 612
rect 576 604 588 612
rect 596 604 600 612
rect 386 602 600 604
rect 0 594 14 602
rect 22 594 34 602
rect 52 594 64 602
rect 82 594 94 602
rect 112 594 124 602
rect 142 594 154 602
rect 172 594 184 602
rect 202 594 214 602
rect 232 594 244 602
rect 252 594 266 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 192 592 214 594
rect 222 592 266 594
rect 274 592 286 602
rect 304 592 316 602
rect 334 594 348 602
rect 356 594 368 602
rect 386 594 398 602
rect 416 594 428 602
rect 446 594 458 602
rect 476 594 488 602
rect 506 594 518 602
rect 536 594 548 602
rect 566 594 578 602
rect 586 594 600 602
rect 334 592 378 594
rect 386 592 408 594
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 0 584 4 592
rect 12 584 24 592
rect 42 584 54 592
rect 72 584 84 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 592
rect 132 582 144 592
rect 162 582 174 592
rect 192 582 204 592
rect 222 582 234 592
rect 242 582 256 592
rect 0 574 14 582
rect 22 574 34 582
rect 52 574 64 582
rect 82 574 94 582
rect 252 574 256 582
rect 344 582 358 592
rect 366 582 378 592
rect 396 582 408 592
rect 426 582 438 592
rect 456 582 468 592
rect 486 582 498 592
rect 516 584 528 592
rect 546 584 558 592
rect 576 584 588 592
rect 596 584 600 592
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 344 574 348 582
rect 506 574 518 582
rect 536 574 548 582
rect 566 574 578 582
rect 586 574 600 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 0 564 4 572
rect 12 564 24 572
rect 42 564 54 572
rect 72 564 84 572
rect 102 564 114 574
rect 132 564 144 574
rect 162 564 174 574
rect 192 564 204 574
rect 222 564 234 574
rect 242 564 256 574
rect 264 564 276 574
rect 294 564 306 574
rect 324 564 336 574
rect 344 564 358 574
rect 366 564 378 574
rect 396 564 408 574
rect 426 564 438 574
rect 456 564 468 574
rect 486 564 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 516 564 528 572
rect 546 564 558 572
rect 576 564 588 572
rect 596 564 600 572
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 192 562 214 564
rect 222 562 286 564
rect 294 562 316 564
rect 324 562 378 564
rect 386 562 408 564
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 0 554 14 562
rect 22 554 34 562
rect 52 554 64 562
rect 82 554 94 562
rect 112 554 124 562
rect 142 554 154 562
rect 172 554 184 562
rect 202 554 214 562
rect 232 554 244 562
rect 252 554 266 562
rect 274 554 286 562
rect 304 554 316 562
rect 334 554 348 562
rect 356 554 368 562
rect 386 554 398 562
rect 416 554 428 562
rect 446 554 458 562
rect 476 554 488 562
rect 506 554 518 562
rect 536 554 548 562
rect 566 554 578 562
rect 586 554 600 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 192 552 214 554
rect 222 552 286 554
rect 294 552 316 554
rect 324 552 378 554
rect 386 552 408 554
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 0 544 4 552
rect 12 544 24 552
rect 42 544 54 552
rect 72 544 84 552
rect 102 544 114 552
rect 132 544 144 552
rect 162 544 174 552
rect 192 544 204 552
rect 222 544 234 552
rect 242 544 256 552
rect 264 544 276 552
rect 294 544 306 552
rect 324 544 336 552
rect 344 544 358 552
rect 366 544 378 552
rect 396 544 408 552
rect 426 544 438 552
rect 456 544 468 552
rect 486 544 498 552
rect 516 544 528 552
rect 546 544 558 552
rect 576 544 588 552
rect 596 544 600 552
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 192 542 214 544
rect 222 542 286 544
rect 294 542 316 544
rect 324 542 378 544
rect 386 542 408 544
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 0 534 14 542
rect 22 534 34 542
rect 52 534 64 542
rect 82 534 94 542
rect 112 534 124 542
rect 142 534 154 542
rect 172 534 184 542
rect 202 534 214 542
rect 232 534 244 542
rect 252 534 266 542
rect 274 534 286 542
rect 304 534 316 542
rect 334 534 348 542
rect 356 534 368 542
rect 386 534 398 542
rect 416 534 428 542
rect 446 534 458 542
rect 476 534 488 542
rect 506 534 518 542
rect 536 534 548 542
rect 566 534 578 542
rect 586 534 600 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 192 532 214 534
rect 222 532 286 534
rect 294 532 316 534
rect 324 532 378 534
rect 386 532 408 534
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 0 524 4 532
rect 12 524 24 532
rect 42 524 54 532
rect 72 524 84 532
rect 102 524 114 532
rect 132 524 144 532
rect 162 524 174 532
rect 192 524 204 532
rect 222 524 234 532
rect 242 524 256 532
rect 264 524 276 532
rect 294 524 306 532
rect 324 524 336 532
rect 344 524 358 532
rect 366 524 378 532
rect 396 524 408 532
rect 426 524 438 532
rect 456 524 468 532
rect 486 524 498 532
rect 516 524 528 532
rect 546 524 558 532
rect 576 524 588 532
rect 596 524 600 532
rect 0 516 600 524
rect 0 8 4 516
rect 12 508 24 516
rect 32 508 44 516
rect 52 508 64 516
rect 72 508 84 516
rect 92 508 104 516
rect 112 508 124 516
rect 132 508 144 516
rect 152 508 164 516
rect 172 508 184 516
rect 192 508 204 516
rect 212 508 224 516
rect 232 508 244 516
rect 252 508 264 516
rect 272 508 284 516
rect 292 508 318 516
rect 326 508 338 516
rect 346 508 358 516
rect 366 508 378 516
rect 386 508 398 516
rect 406 508 418 516
rect 426 508 438 516
rect 446 508 458 516
rect 466 508 478 516
rect 486 508 498 516
rect 506 508 518 516
rect 526 508 538 516
rect 546 508 558 516
rect 566 508 578 516
rect 12 502 588 508
rect 12 14 16 502
rect 584 14 588 502
rect 12 12 588 14
rect 0 4 14 8
rect 182 4 408 12
rect 596 8 600 516
rect 586 4 600 8
rect 0 -2 600 4
<< psubstratepcontact >>
rect 2 1320 190 1338
rect 408 1320 576 1338
rect 2 840 20 1320
rect 580 840 598 1338
rect 4 828 12 836
rect 24 828 42 836
rect 54 828 72 836
rect 84 828 102 836
rect 114 828 132 836
rect 144 828 162 836
rect 174 828 182 836
rect 296 828 304 836
rect 418 828 426 836
rect 438 828 456 836
rect 468 828 486 836
rect 498 828 516 836
rect 528 828 546 836
rect 558 828 576 836
rect 588 828 596 836
rect 34 826 42 828
rect 64 826 72 828
rect 94 826 102 828
rect 124 826 132 828
rect 154 826 162 828
rect 438 826 446 828
rect 468 826 476 828
rect 498 826 506 828
rect 528 826 536 828
rect 558 826 566 828
rect 14 818 22 826
rect 34 818 52 826
rect 64 818 82 826
rect 94 818 112 826
rect 124 818 142 826
rect 154 818 172 826
rect 184 818 192 826
rect 286 818 294 826
rect 306 818 314 826
rect 408 818 416 826
rect 428 818 446 826
rect 458 818 476 826
rect 488 818 506 826
rect 518 818 536 826
rect 548 818 566 826
rect 578 818 586 826
rect 34 816 42 818
rect 64 816 72 818
rect 94 816 102 818
rect 124 816 132 818
rect 154 816 162 818
rect 438 816 446 818
rect 468 816 476 818
rect 498 816 506 818
rect 528 816 536 818
rect 558 816 566 818
rect 4 808 12 816
rect 24 808 42 816
rect 54 808 72 816
rect 84 808 102 816
rect 114 808 132 816
rect 144 808 162 816
rect 174 808 182 816
rect 296 808 304 816
rect 418 808 426 816
rect 438 808 456 816
rect 468 808 486 816
rect 498 808 516 816
rect 528 808 546 816
rect 558 808 576 816
rect 588 808 596 816
rect 34 806 42 808
rect 64 806 72 808
rect 94 806 102 808
rect 124 806 132 808
rect 154 806 162 808
rect 438 806 446 808
rect 468 806 476 808
rect 498 806 506 808
rect 528 806 536 808
rect 558 806 566 808
rect 14 798 22 806
rect 34 798 52 806
rect 64 798 82 806
rect 94 798 112 806
rect 124 798 142 806
rect 154 798 172 806
rect 184 798 192 806
rect 286 798 294 806
rect 306 798 314 806
rect 408 798 416 806
rect 428 798 446 806
rect 458 798 476 806
rect 488 798 506 806
rect 518 798 536 806
rect 548 798 566 806
rect 578 798 586 806
rect 34 796 42 798
rect 64 796 72 798
rect 94 796 102 798
rect 124 796 132 798
rect 154 796 162 798
rect 438 796 446 798
rect 468 796 476 798
rect 498 796 506 798
rect 528 796 536 798
rect 558 796 566 798
rect 4 788 12 796
rect 24 788 42 796
rect 54 788 72 796
rect 84 788 102 796
rect 114 788 132 796
rect 144 788 162 796
rect 174 788 182 796
rect 296 788 304 796
rect 418 788 426 796
rect 438 788 456 796
rect 468 788 486 796
rect 498 788 516 796
rect 528 788 546 796
rect 558 788 576 796
rect 588 788 596 796
rect 34 786 42 788
rect 64 786 72 788
rect 94 786 102 788
rect 124 786 132 788
rect 154 786 162 788
rect 438 786 446 788
rect 468 786 476 788
rect 498 786 506 788
rect 528 786 536 788
rect 558 786 566 788
rect 14 778 22 786
rect 34 778 52 786
rect 64 778 82 786
rect 34 776 42 778
rect 64 776 72 778
rect 94 776 112 786
rect 124 776 142 786
rect 154 776 172 786
rect 184 776 192 786
rect 4 768 12 776
rect 24 768 42 776
rect 54 768 72 776
rect 84 768 192 776
rect 286 776 294 786
rect 306 776 314 786
rect 286 768 314 776
rect 408 776 416 786
rect 428 776 446 786
rect 458 776 476 786
rect 488 776 506 786
rect 518 778 536 786
rect 548 778 566 786
rect 578 778 586 786
rect 528 776 536 778
rect 558 776 566 778
rect 408 768 516 776
rect 528 768 546 776
rect 558 768 576 776
rect 588 768 596 776
rect 34 766 42 768
rect 64 766 72 768
rect 14 758 22 766
rect 34 758 52 766
rect 64 758 82 766
rect 94 758 112 768
rect 124 758 142 768
rect 154 758 172 768
rect 184 758 192 768
rect 296 758 304 768
rect 408 758 416 768
rect 428 758 446 768
rect 458 758 476 768
rect 488 758 506 768
rect 528 766 536 768
rect 558 766 566 768
rect 518 758 536 766
rect 548 758 566 766
rect 578 758 586 766
rect 34 756 42 758
rect 64 756 72 758
rect 94 756 102 758
rect 124 756 132 758
rect 154 756 162 758
rect 438 756 446 758
rect 468 756 476 758
rect 498 756 506 758
rect 528 756 536 758
rect 558 756 566 758
rect 4 748 12 756
rect 24 748 42 756
rect 54 748 72 756
rect 84 748 102 756
rect 114 748 132 756
rect 144 748 162 756
rect 174 748 182 756
rect 286 748 294 756
rect 306 748 314 756
rect 418 748 426 756
rect 438 748 456 756
rect 468 748 486 756
rect 498 748 516 756
rect 528 748 546 756
rect 558 748 576 756
rect 588 748 596 756
rect 34 746 42 748
rect 64 746 72 748
rect 94 746 102 748
rect 124 746 132 748
rect 154 746 162 748
rect 438 746 446 748
rect 468 746 476 748
rect 498 746 506 748
rect 528 746 536 748
rect 558 746 566 748
rect 14 738 22 746
rect 34 738 52 746
rect 64 738 82 746
rect 94 738 112 746
rect 124 738 142 746
rect 154 738 172 746
rect 184 738 192 746
rect 296 738 304 746
rect 408 738 416 746
rect 428 738 446 746
rect 458 738 476 746
rect 488 738 506 746
rect 518 738 536 746
rect 548 738 566 746
rect 578 738 586 746
rect 4 728 12 736
rect 24 728 32 736
rect 286 728 294 736
rect 306 728 314 736
rect 568 728 576 736
rect 588 728 596 736
rect 14 718 22 726
rect 34 718 52 726
rect 64 718 82 726
rect 94 718 112 726
rect 124 718 142 726
rect 154 718 172 726
rect 184 718 192 726
rect 296 718 304 726
rect 408 718 416 726
rect 428 718 446 726
rect 458 718 476 726
rect 488 718 506 726
rect 518 718 536 726
rect 548 718 566 726
rect 578 718 586 726
rect 34 716 42 718
rect 64 716 72 718
rect 94 716 102 718
rect 124 716 132 718
rect 154 716 162 718
rect 438 716 446 718
rect 468 716 476 718
rect 498 716 506 718
rect 528 716 536 718
rect 558 716 566 718
rect 4 708 12 716
rect 24 708 42 716
rect 54 708 72 716
rect 84 708 102 716
rect 114 708 132 716
rect 144 708 162 716
rect 174 708 182 716
rect 286 708 294 716
rect 306 708 314 716
rect 418 708 426 716
rect 438 708 456 716
rect 468 708 486 716
rect 498 708 516 716
rect 528 708 546 716
rect 558 708 576 716
rect 588 708 596 716
rect 34 706 42 708
rect 64 706 72 708
rect 94 706 102 708
rect 124 706 132 708
rect 154 706 162 708
rect 438 706 446 708
rect 468 706 476 708
rect 498 706 506 708
rect 528 706 536 708
rect 558 706 566 708
rect 14 698 22 706
rect 34 698 52 706
rect 64 698 82 706
rect 94 698 112 706
rect 124 698 142 706
rect 154 698 172 706
rect 184 698 192 706
rect 408 698 416 706
rect 428 698 446 706
rect 458 698 476 706
rect 488 698 506 706
rect 518 698 536 706
rect 548 698 566 706
rect 578 698 586 706
rect 34 696 42 698
rect 64 696 72 698
rect 94 696 102 698
rect 124 696 132 698
rect 154 696 162 698
rect 438 696 446 698
rect 468 696 476 698
rect 498 696 506 698
rect 528 696 536 698
rect 558 696 566 698
rect 4 688 12 696
rect 24 688 42 696
rect 54 688 72 696
rect 84 688 102 696
rect 114 688 132 696
rect 144 688 162 696
rect 174 688 182 696
rect 286 688 314 696
rect 418 688 426 696
rect 438 688 456 696
rect 468 688 486 696
rect 498 688 516 696
rect 528 688 546 696
rect 558 688 576 696
rect 588 688 596 696
rect 38 466 196 484
rect 38 456 56 466
rect 38 436 56 444
rect 78 456 196 466
rect 404 466 562 484
rect 291 436 309 444
rect 404 456 522 466
rect 544 456 562 466
rect 544 436 562 444
rect 38 416 56 424
rect 38 396 56 404
rect 38 376 56 384
rect 38 356 56 364
rect 38 336 56 344
rect 38 316 56 324
rect 38 296 56 304
rect 38 276 56 284
rect 38 256 56 264
rect 38 236 56 244
rect 38 216 56 224
rect 38 196 56 204
rect 38 176 56 184
rect 38 156 56 164
rect 38 136 56 144
rect 38 116 56 124
rect 38 96 56 104
rect 38 76 56 84
rect 291 420 309 428
rect 291 404 309 412
rect 291 260 309 268
rect 291 244 309 252
rect 291 116 309 124
rect 291 100 309 108
rect 291 84 309 92
rect 38 56 56 64
rect 544 416 562 424
rect 544 396 562 404
rect 544 376 562 384
rect 544 356 562 364
rect 544 336 562 344
rect 544 316 562 324
rect 544 296 562 304
rect 544 276 562 284
rect 544 256 562 264
rect 544 236 562 244
rect 544 216 562 224
rect 544 196 562 204
rect 544 176 562 184
rect 544 156 562 164
rect 544 136 562 144
rect 544 116 562 124
rect 544 96 562 104
rect 291 68 309 76
rect 544 76 562 84
rect 544 56 562 64
rect 68 46 76 54
rect 88 46 96 54
rect 108 46 116 54
rect 128 46 136 54
rect 148 46 156 54
rect 168 46 176 54
rect 188 46 196 54
rect 404 46 412 54
rect 424 46 432 54
rect 444 46 452 54
rect 464 46 472 54
rect 484 46 492 54
rect 504 46 512 54
rect 524 46 532 54
rect 38 36 66 44
rect 78 36 86 44
rect 98 36 106 44
rect 118 36 126 44
rect 138 36 146 44
rect 158 36 166 44
rect 178 36 186 44
rect 414 36 422 44
rect 434 36 442 44
rect 454 36 462 44
rect 474 36 482 44
rect 494 36 502 44
rect 514 36 522 44
rect 534 36 562 44
<< nsubstratencontact >>
rect 46 1290 54 1298
rect 66 1290 84 1298
rect 96 1290 114 1298
rect 126 1290 144 1298
rect 156 1290 174 1298
rect 186 1290 204 1298
rect 216 1290 234 1298
rect 246 1290 264 1298
rect 276 1290 294 1298
rect 306 1290 324 1298
rect 336 1290 354 1298
rect 366 1290 384 1298
rect 396 1290 414 1298
rect 426 1290 444 1298
rect 456 1290 474 1298
rect 486 1290 504 1298
rect 516 1290 534 1298
rect 546 1290 554 1298
rect 76 1288 84 1290
rect 106 1288 114 1290
rect 136 1288 144 1290
rect 166 1288 174 1290
rect 196 1288 204 1290
rect 226 1288 234 1290
rect 256 1288 264 1290
rect 286 1288 294 1290
rect 316 1288 324 1290
rect 346 1288 354 1290
rect 376 1288 384 1290
rect 406 1288 414 1290
rect 436 1288 444 1290
rect 466 1288 474 1290
rect 496 1288 504 1290
rect 526 1288 534 1290
rect 56 1280 64 1288
rect 76 1280 94 1288
rect 106 1280 124 1288
rect 136 1280 154 1288
rect 166 1280 184 1288
rect 196 1280 214 1288
rect 226 1280 244 1288
rect 256 1280 274 1288
rect 286 1280 304 1288
rect 316 1280 334 1288
rect 346 1280 364 1288
rect 376 1280 394 1288
rect 406 1280 424 1288
rect 436 1280 454 1288
rect 466 1280 484 1288
rect 496 1280 514 1288
rect 526 1280 544 1288
rect 76 1278 84 1280
rect 106 1278 114 1280
rect 136 1278 144 1280
rect 166 1278 174 1280
rect 196 1278 204 1280
rect 226 1278 234 1280
rect 256 1278 264 1280
rect 286 1278 294 1280
rect 316 1278 324 1280
rect 346 1278 354 1280
rect 376 1278 384 1280
rect 406 1278 414 1280
rect 436 1278 444 1280
rect 466 1278 474 1280
rect 496 1278 504 1280
rect 526 1278 534 1280
rect 46 1270 54 1278
rect 66 1270 84 1278
rect 96 1270 114 1278
rect 126 1270 144 1278
rect 156 1270 174 1278
rect 186 1270 204 1278
rect 216 1270 234 1278
rect 246 1270 264 1278
rect 276 1270 294 1278
rect 306 1270 324 1278
rect 336 1270 354 1278
rect 366 1270 384 1278
rect 396 1270 414 1278
rect 426 1270 444 1278
rect 456 1270 474 1278
rect 486 1270 504 1278
rect 516 1270 534 1278
rect 546 1270 554 1278
rect 76 1268 84 1270
rect 106 1268 114 1270
rect 136 1268 144 1270
rect 166 1268 174 1270
rect 196 1268 204 1270
rect 226 1268 234 1270
rect 256 1268 264 1270
rect 286 1268 294 1270
rect 316 1268 324 1270
rect 346 1268 354 1270
rect 376 1268 384 1270
rect 406 1268 414 1270
rect 436 1268 444 1270
rect 466 1268 474 1270
rect 496 1268 504 1270
rect 526 1268 534 1270
rect 56 1260 64 1268
rect 76 1260 94 1268
rect 106 1260 124 1268
rect 136 1260 154 1268
rect 166 1260 184 1268
rect 196 1260 214 1268
rect 226 1260 244 1268
rect 256 1260 274 1268
rect 286 1260 304 1268
rect 316 1260 334 1268
rect 346 1260 364 1268
rect 376 1260 394 1268
rect 406 1260 424 1268
rect 436 1260 454 1268
rect 466 1260 484 1268
rect 496 1260 514 1268
rect 526 1260 544 1268
rect 76 1258 84 1260
rect 106 1258 114 1260
rect 136 1258 144 1260
rect 166 1258 174 1260
rect 196 1258 204 1260
rect 226 1258 234 1260
rect 256 1258 264 1260
rect 286 1258 294 1260
rect 316 1258 324 1260
rect 346 1258 354 1260
rect 376 1258 384 1260
rect 406 1258 414 1260
rect 436 1258 444 1260
rect 466 1258 474 1260
rect 496 1258 504 1260
rect 526 1258 534 1260
rect 46 1250 54 1258
rect 66 1250 84 1258
rect 96 1250 114 1258
rect 126 1250 144 1258
rect 156 1250 174 1258
rect 186 1250 204 1258
rect 216 1250 234 1258
rect 246 1250 264 1258
rect 276 1250 294 1258
rect 306 1250 324 1258
rect 336 1250 354 1258
rect 366 1250 384 1258
rect 396 1250 414 1258
rect 426 1250 444 1258
rect 456 1250 474 1258
rect 486 1250 504 1258
rect 516 1250 534 1258
rect 546 1250 554 1258
rect 76 1248 84 1250
rect 106 1248 114 1250
rect 136 1248 144 1250
rect 166 1248 174 1250
rect 196 1248 204 1250
rect 226 1248 234 1250
rect 256 1248 264 1250
rect 286 1248 294 1250
rect 316 1248 324 1250
rect 346 1248 354 1250
rect 376 1248 384 1250
rect 406 1248 414 1250
rect 436 1248 444 1250
rect 466 1248 474 1250
rect 496 1248 504 1250
rect 526 1248 534 1250
rect 56 1240 64 1248
rect 76 1240 94 1248
rect 106 1240 124 1248
rect 136 1240 154 1248
rect 166 1240 184 1248
rect 196 1240 214 1248
rect 226 1240 244 1248
rect 256 1240 274 1248
rect 286 1240 304 1248
rect 316 1240 334 1248
rect 346 1240 364 1248
rect 376 1240 394 1248
rect 406 1240 424 1248
rect 436 1240 454 1248
rect 466 1240 484 1248
rect 496 1240 514 1248
rect 526 1240 544 1248
rect 76 1238 84 1240
rect 106 1238 114 1240
rect 136 1238 144 1240
rect 166 1238 174 1240
rect 196 1238 204 1240
rect 226 1238 234 1240
rect 256 1238 264 1240
rect 286 1238 294 1240
rect 316 1238 324 1240
rect 346 1238 354 1240
rect 376 1238 384 1240
rect 406 1238 414 1240
rect 436 1238 444 1240
rect 466 1238 474 1240
rect 496 1238 504 1240
rect 526 1238 534 1240
rect 46 1230 54 1238
rect 66 1230 84 1238
rect 96 1230 114 1238
rect 126 1230 144 1238
rect 156 1230 174 1238
rect 186 1230 204 1238
rect 216 1230 234 1238
rect 246 1230 264 1238
rect 276 1230 294 1238
rect 306 1230 324 1238
rect 336 1230 354 1238
rect 366 1230 384 1238
rect 396 1230 414 1238
rect 426 1230 444 1238
rect 456 1230 474 1238
rect 486 1230 504 1238
rect 516 1230 534 1238
rect 546 1230 554 1238
rect 76 1228 84 1230
rect 106 1228 114 1230
rect 136 1228 144 1230
rect 166 1228 174 1230
rect 196 1228 204 1230
rect 226 1228 234 1230
rect 256 1228 264 1230
rect 286 1228 294 1230
rect 316 1228 324 1230
rect 346 1228 354 1230
rect 376 1228 384 1230
rect 406 1228 414 1230
rect 436 1228 444 1230
rect 466 1228 474 1230
rect 496 1228 504 1230
rect 526 1228 534 1230
rect 56 1220 64 1228
rect 76 1220 94 1228
rect 106 1220 124 1228
rect 136 1220 154 1228
rect 166 1220 184 1228
rect 196 1220 214 1228
rect 226 1220 244 1228
rect 256 1220 274 1228
rect 286 1220 304 1228
rect 316 1220 334 1228
rect 346 1220 364 1228
rect 376 1220 394 1228
rect 406 1220 424 1228
rect 436 1220 454 1228
rect 466 1220 484 1228
rect 496 1220 514 1228
rect 526 1220 544 1228
rect 76 1218 84 1220
rect 106 1218 114 1220
rect 136 1218 144 1220
rect 166 1218 174 1220
rect 196 1218 204 1220
rect 226 1218 234 1220
rect 256 1218 264 1220
rect 286 1218 294 1220
rect 316 1218 324 1220
rect 346 1218 354 1220
rect 376 1218 384 1220
rect 406 1218 414 1220
rect 436 1218 444 1220
rect 466 1218 474 1220
rect 496 1218 504 1220
rect 526 1218 534 1220
rect 46 1210 54 1218
rect 66 1210 84 1218
rect 96 1210 114 1218
rect 126 1210 144 1218
rect 156 1210 174 1218
rect 186 1210 204 1218
rect 216 1210 234 1218
rect 246 1210 264 1218
rect 276 1210 294 1218
rect 306 1210 324 1218
rect 336 1210 354 1218
rect 366 1210 384 1218
rect 396 1210 414 1218
rect 426 1210 444 1218
rect 456 1210 474 1218
rect 486 1210 504 1218
rect 516 1210 534 1218
rect 546 1210 554 1218
rect 76 1208 84 1210
rect 106 1208 114 1210
rect 136 1208 144 1210
rect 166 1208 174 1210
rect 196 1208 204 1210
rect 226 1208 234 1210
rect 256 1208 264 1210
rect 286 1208 294 1210
rect 316 1208 324 1210
rect 346 1208 354 1210
rect 376 1208 384 1210
rect 406 1208 414 1210
rect 436 1208 444 1210
rect 466 1208 474 1210
rect 496 1208 504 1210
rect 526 1208 534 1210
rect 56 1200 64 1208
rect 76 1200 94 1208
rect 106 1200 124 1208
rect 136 1200 154 1208
rect 166 1200 184 1208
rect 196 1200 214 1208
rect 226 1200 244 1208
rect 256 1200 274 1208
rect 286 1200 304 1208
rect 316 1200 334 1208
rect 346 1200 364 1208
rect 376 1200 394 1208
rect 406 1200 424 1208
rect 436 1200 454 1208
rect 466 1200 484 1208
rect 496 1200 514 1208
rect 526 1200 544 1208
rect 76 1198 84 1200
rect 106 1198 114 1200
rect 136 1198 144 1200
rect 166 1198 174 1200
rect 196 1198 204 1200
rect 226 1198 234 1200
rect 256 1198 264 1200
rect 286 1198 294 1200
rect 316 1198 324 1200
rect 346 1198 354 1200
rect 376 1198 384 1200
rect 406 1198 414 1200
rect 436 1198 444 1200
rect 466 1198 474 1200
rect 496 1198 504 1200
rect 526 1198 534 1200
rect 46 1190 54 1198
rect 66 1190 84 1198
rect 96 1190 114 1198
rect 126 1190 144 1198
rect 156 1190 174 1198
rect 186 1190 204 1198
rect 216 1190 234 1198
rect 246 1190 264 1198
rect 276 1190 294 1198
rect 306 1190 324 1198
rect 336 1190 354 1198
rect 366 1190 384 1198
rect 396 1190 414 1198
rect 426 1190 444 1198
rect 456 1190 474 1198
rect 486 1190 504 1198
rect 516 1190 534 1198
rect 546 1190 554 1198
rect 76 1188 84 1190
rect 526 1188 534 1190
rect 56 1180 64 1188
rect 76 1180 94 1188
rect 506 1180 514 1188
rect 526 1180 544 1188
rect 76 1178 84 1180
rect 526 1178 534 1180
rect 46 1170 54 1178
rect 66 1170 84 1178
rect 96 1170 114 1178
rect 126 1170 144 1178
rect 156 1170 174 1178
rect 186 1170 204 1178
rect 216 1170 234 1178
rect 246 1170 264 1178
rect 276 1170 294 1178
rect 306 1170 324 1178
rect 336 1170 354 1178
rect 366 1170 384 1178
rect 396 1170 414 1178
rect 426 1170 444 1178
rect 456 1170 474 1178
rect 486 1170 504 1178
rect 516 1170 534 1178
rect 546 1170 554 1178
rect 76 1168 84 1170
rect 106 1168 114 1170
rect 136 1168 144 1170
rect 166 1168 174 1170
rect 196 1168 204 1170
rect 226 1168 234 1170
rect 256 1168 264 1170
rect 286 1168 294 1170
rect 316 1168 324 1170
rect 346 1168 354 1170
rect 376 1168 384 1170
rect 406 1168 414 1170
rect 436 1168 444 1170
rect 466 1168 474 1170
rect 496 1168 504 1170
rect 526 1168 534 1170
rect 56 1160 64 1168
rect 76 1160 94 1168
rect 106 1160 124 1168
rect 136 1160 154 1168
rect 166 1160 184 1168
rect 196 1160 214 1168
rect 226 1160 244 1168
rect 256 1160 274 1168
rect 286 1160 304 1168
rect 316 1160 334 1168
rect 346 1160 364 1168
rect 376 1160 394 1168
rect 406 1160 424 1168
rect 436 1160 454 1168
rect 466 1160 484 1168
rect 496 1160 514 1168
rect 526 1160 544 1168
rect 76 1158 84 1160
rect 106 1158 114 1160
rect 136 1158 144 1160
rect 166 1158 174 1160
rect 196 1158 204 1160
rect 226 1158 234 1160
rect 256 1158 264 1160
rect 286 1158 294 1160
rect 316 1158 324 1160
rect 346 1158 354 1160
rect 376 1158 384 1160
rect 406 1158 414 1160
rect 436 1158 444 1160
rect 466 1158 474 1160
rect 496 1158 504 1160
rect 526 1158 534 1160
rect 46 1150 54 1158
rect 66 1150 84 1158
rect 96 1150 114 1158
rect 126 1150 144 1158
rect 156 1150 174 1158
rect 186 1150 204 1158
rect 216 1150 234 1158
rect 246 1150 264 1158
rect 276 1150 294 1158
rect 306 1150 324 1158
rect 336 1150 354 1158
rect 366 1150 384 1158
rect 396 1150 414 1158
rect 426 1150 444 1158
rect 456 1150 474 1158
rect 486 1150 504 1158
rect 516 1150 534 1158
rect 546 1150 554 1158
rect 76 1148 84 1150
rect 106 1148 114 1150
rect 136 1148 144 1150
rect 166 1148 174 1150
rect 196 1148 204 1150
rect 226 1148 234 1150
rect 256 1148 264 1150
rect 286 1148 294 1150
rect 316 1148 324 1150
rect 346 1148 354 1150
rect 376 1148 384 1150
rect 406 1148 414 1150
rect 436 1148 444 1150
rect 466 1148 474 1150
rect 496 1148 504 1150
rect 526 1148 534 1150
rect 56 1140 64 1148
rect 76 1140 94 1148
rect 106 1140 124 1148
rect 136 1140 154 1148
rect 166 1140 184 1148
rect 196 1140 214 1148
rect 226 1140 244 1148
rect 256 1140 274 1148
rect 286 1140 304 1148
rect 316 1140 334 1148
rect 346 1140 364 1148
rect 376 1140 394 1148
rect 406 1140 424 1148
rect 436 1140 454 1148
rect 466 1140 484 1148
rect 496 1140 514 1148
rect 526 1140 544 1148
rect 76 1138 84 1140
rect 106 1138 114 1140
rect 136 1138 144 1140
rect 166 1138 174 1140
rect 196 1138 204 1140
rect 226 1138 234 1140
rect 256 1138 264 1140
rect 286 1138 294 1140
rect 316 1138 324 1140
rect 346 1138 354 1140
rect 376 1138 384 1140
rect 406 1138 414 1140
rect 436 1138 444 1140
rect 466 1138 474 1140
rect 496 1138 504 1140
rect 526 1138 534 1140
rect 46 1130 54 1138
rect 66 1130 84 1138
rect 96 1130 114 1138
rect 126 1130 144 1138
rect 156 1130 174 1138
rect 186 1130 204 1138
rect 216 1130 234 1138
rect 246 1130 264 1138
rect 276 1130 294 1138
rect 306 1130 324 1138
rect 336 1130 354 1138
rect 366 1130 384 1138
rect 396 1130 414 1138
rect 426 1130 444 1138
rect 456 1130 474 1138
rect 486 1130 504 1138
rect 516 1130 534 1138
rect 546 1130 554 1138
rect 76 1128 84 1130
rect 106 1128 114 1130
rect 136 1128 144 1130
rect 166 1128 174 1130
rect 196 1128 204 1130
rect 226 1128 234 1130
rect 256 1128 264 1130
rect 286 1128 294 1130
rect 316 1128 324 1130
rect 346 1128 354 1130
rect 376 1128 384 1130
rect 406 1128 414 1130
rect 436 1128 444 1130
rect 466 1128 474 1130
rect 496 1128 504 1130
rect 526 1128 534 1130
rect 56 1120 64 1128
rect 76 1120 94 1128
rect 106 1120 124 1128
rect 136 1120 154 1128
rect 166 1120 184 1128
rect 196 1120 214 1128
rect 226 1120 244 1128
rect 256 1120 274 1128
rect 286 1120 304 1128
rect 316 1120 334 1128
rect 346 1120 364 1128
rect 376 1120 394 1128
rect 406 1120 424 1128
rect 436 1120 454 1128
rect 466 1120 484 1128
rect 496 1120 514 1128
rect 46 1110 54 1118
rect 66 1110 74 1118
rect 86 1108 94 1120
rect 506 1108 514 1120
rect 56 1100 64 1108
rect 76 1100 94 1108
rect 106 1100 124 1108
rect 136 1100 154 1108
rect 166 1100 184 1108
rect 196 1100 214 1108
rect 226 1100 244 1108
rect 256 1100 274 1108
rect 286 1100 304 1108
rect 316 1100 334 1108
rect 346 1100 364 1108
rect 376 1100 394 1108
rect 406 1100 424 1108
rect 436 1100 454 1108
rect 466 1100 484 1108
rect 496 1100 514 1108
rect 526 1120 544 1128
rect 526 1108 534 1120
rect 546 1110 554 1118
rect 526 1100 544 1108
rect 76 1098 84 1100
rect 106 1098 114 1100
rect 136 1098 144 1100
rect 166 1098 174 1100
rect 196 1098 204 1100
rect 226 1098 234 1100
rect 256 1098 264 1100
rect 286 1098 294 1100
rect 316 1098 324 1100
rect 346 1098 354 1100
rect 376 1098 384 1100
rect 406 1098 414 1100
rect 436 1098 444 1100
rect 466 1098 474 1100
rect 496 1098 504 1100
rect 526 1098 534 1100
rect 46 1090 54 1098
rect 66 1090 84 1098
rect 96 1090 114 1098
rect 126 1090 144 1098
rect 156 1090 174 1098
rect 186 1090 204 1098
rect 216 1090 234 1098
rect 246 1090 264 1098
rect 276 1090 294 1098
rect 306 1090 324 1098
rect 336 1090 354 1098
rect 366 1090 384 1098
rect 396 1090 414 1098
rect 426 1090 444 1098
rect 456 1090 474 1098
rect 486 1090 504 1098
rect 516 1090 534 1098
rect 546 1090 554 1098
rect 76 1088 84 1090
rect 106 1088 114 1090
rect 136 1088 144 1090
rect 166 1088 174 1090
rect 196 1088 204 1090
rect 226 1088 234 1090
rect 256 1088 264 1090
rect 286 1088 294 1090
rect 316 1088 324 1090
rect 346 1088 354 1090
rect 376 1088 384 1090
rect 406 1088 414 1090
rect 436 1088 444 1090
rect 466 1088 474 1090
rect 496 1088 504 1090
rect 526 1088 534 1090
rect 56 1080 64 1088
rect 76 1080 94 1088
rect 106 1080 124 1088
rect 136 1080 154 1088
rect 166 1080 184 1088
rect 196 1080 214 1088
rect 226 1080 244 1088
rect 256 1080 274 1088
rect 286 1080 304 1088
rect 316 1080 334 1088
rect 346 1080 364 1088
rect 376 1080 394 1088
rect 406 1080 424 1088
rect 436 1080 454 1088
rect 466 1080 484 1088
rect 496 1080 514 1088
rect 526 1080 544 1088
rect 76 1078 84 1080
rect 106 1078 114 1080
rect 136 1078 144 1080
rect 166 1078 174 1080
rect 196 1078 204 1080
rect 226 1078 234 1080
rect 256 1078 264 1080
rect 286 1078 294 1080
rect 316 1078 324 1080
rect 346 1078 354 1080
rect 376 1078 384 1080
rect 406 1078 414 1080
rect 436 1078 444 1080
rect 466 1078 474 1080
rect 496 1078 504 1080
rect 526 1078 534 1080
rect 46 1070 54 1078
rect 66 1070 84 1078
rect 96 1070 114 1078
rect 126 1070 144 1078
rect 156 1070 174 1078
rect 186 1070 204 1078
rect 216 1070 234 1078
rect 246 1070 264 1078
rect 276 1070 294 1078
rect 306 1070 324 1078
rect 336 1070 354 1078
rect 366 1070 384 1078
rect 396 1070 414 1078
rect 426 1070 444 1078
rect 456 1070 474 1078
rect 486 1070 504 1078
rect 516 1070 534 1078
rect 546 1070 554 1078
rect 76 1068 84 1070
rect 106 1068 114 1070
rect 136 1068 144 1070
rect 166 1068 174 1070
rect 196 1068 204 1070
rect 226 1068 234 1070
rect 256 1068 264 1070
rect 286 1068 294 1070
rect 316 1068 324 1070
rect 346 1068 354 1070
rect 376 1068 384 1070
rect 406 1068 414 1070
rect 436 1068 444 1070
rect 466 1068 474 1070
rect 496 1068 504 1070
rect 526 1068 534 1070
rect 56 1060 64 1068
rect 76 1060 94 1068
rect 106 1060 124 1068
rect 136 1060 154 1068
rect 166 1060 184 1068
rect 196 1060 214 1068
rect 226 1060 244 1068
rect 256 1060 274 1068
rect 286 1060 304 1068
rect 316 1060 334 1068
rect 346 1060 364 1068
rect 376 1060 394 1068
rect 406 1060 424 1068
rect 436 1060 454 1068
rect 466 1060 484 1068
rect 496 1060 514 1068
rect 526 1060 544 1068
rect 76 1058 84 1060
rect 106 1058 114 1060
rect 136 1058 144 1060
rect 166 1058 174 1060
rect 196 1058 204 1060
rect 226 1058 234 1060
rect 256 1058 264 1060
rect 286 1058 294 1060
rect 316 1058 324 1060
rect 346 1058 354 1060
rect 376 1058 384 1060
rect 406 1058 414 1060
rect 436 1058 444 1060
rect 466 1058 474 1060
rect 496 1058 504 1060
rect 526 1058 534 1060
rect 46 1050 54 1058
rect 66 1050 84 1058
rect 96 1050 114 1058
rect 126 1050 144 1058
rect 156 1050 174 1058
rect 186 1050 204 1058
rect 216 1050 234 1058
rect 246 1050 264 1058
rect 276 1050 294 1058
rect 306 1050 324 1058
rect 336 1050 354 1058
rect 366 1050 384 1058
rect 396 1050 414 1058
rect 426 1050 444 1058
rect 456 1050 474 1058
rect 486 1050 504 1058
rect 516 1050 534 1058
rect 546 1050 554 1058
rect 76 1048 84 1050
rect 106 1048 114 1050
rect 136 1048 144 1050
rect 166 1048 174 1050
rect 196 1048 204 1050
rect 226 1048 234 1050
rect 256 1048 264 1050
rect 286 1048 294 1050
rect 316 1048 324 1050
rect 346 1048 354 1050
rect 376 1048 384 1050
rect 406 1048 414 1050
rect 436 1048 444 1050
rect 466 1048 474 1050
rect 496 1048 504 1050
rect 526 1048 534 1050
rect 56 1040 64 1048
rect 76 1040 94 1048
rect 106 1040 124 1048
rect 136 1040 154 1048
rect 166 1040 184 1048
rect 196 1040 214 1048
rect 226 1040 244 1048
rect 256 1040 274 1048
rect 286 1040 304 1048
rect 316 1040 334 1048
rect 346 1040 364 1048
rect 376 1040 394 1048
rect 406 1040 424 1048
rect 436 1040 454 1048
rect 466 1040 484 1048
rect 496 1040 514 1048
rect 76 1038 84 1040
rect 46 1030 54 1038
rect 66 1030 84 1038
rect 76 1028 84 1030
rect 506 1028 514 1040
rect 56 1020 64 1028
rect 76 1020 94 1028
rect 106 1020 124 1028
rect 136 1020 154 1028
rect 166 1020 184 1028
rect 196 1020 214 1028
rect 226 1020 244 1028
rect 256 1020 274 1028
rect 286 1020 304 1028
rect 316 1020 334 1028
rect 346 1020 364 1028
rect 376 1020 394 1028
rect 406 1020 424 1028
rect 436 1020 454 1028
rect 466 1020 484 1028
rect 496 1020 514 1028
rect 526 1040 544 1048
rect 526 1028 534 1040
rect 546 1030 554 1038
rect 526 1020 544 1028
rect 76 1018 84 1020
rect 106 1018 114 1020
rect 136 1018 144 1020
rect 166 1018 174 1020
rect 196 1018 204 1020
rect 226 1018 234 1020
rect 256 1018 264 1020
rect 286 1018 294 1020
rect 316 1018 324 1020
rect 346 1018 354 1020
rect 376 1018 384 1020
rect 406 1018 414 1020
rect 436 1018 444 1020
rect 466 1018 474 1020
rect 496 1018 504 1020
rect 526 1018 534 1020
rect 46 1010 54 1018
rect 66 1010 84 1018
rect 96 1010 114 1018
rect 126 1010 144 1018
rect 156 1010 174 1018
rect 186 1010 204 1018
rect 216 1010 234 1018
rect 246 1010 264 1018
rect 276 1010 294 1018
rect 306 1010 324 1018
rect 336 1010 354 1018
rect 366 1010 384 1018
rect 396 1010 414 1018
rect 426 1010 444 1018
rect 456 1010 474 1018
rect 486 1010 504 1018
rect 516 1010 534 1018
rect 546 1010 554 1018
rect 76 1008 84 1010
rect 106 1008 114 1010
rect 136 1008 144 1010
rect 166 1008 174 1010
rect 196 1008 204 1010
rect 226 1008 234 1010
rect 256 1008 264 1010
rect 286 1008 294 1010
rect 316 1008 324 1010
rect 346 1008 354 1010
rect 376 1008 384 1010
rect 406 1008 414 1010
rect 436 1008 444 1010
rect 466 1008 474 1010
rect 496 1008 504 1010
rect 526 1008 534 1010
rect 56 1000 64 1008
rect 76 1000 94 1008
rect 106 1000 124 1008
rect 136 1000 154 1008
rect 166 1000 184 1008
rect 196 1000 214 1008
rect 226 1000 244 1008
rect 256 1000 274 1008
rect 286 1000 304 1008
rect 316 1000 334 1008
rect 346 1000 364 1008
rect 376 1000 394 1008
rect 406 1000 424 1008
rect 436 1000 454 1008
rect 466 1000 484 1008
rect 496 1000 514 1008
rect 526 1000 544 1008
rect 76 998 84 1000
rect 106 998 114 1000
rect 136 998 144 1000
rect 166 998 174 1000
rect 196 998 204 1000
rect 226 998 234 1000
rect 256 998 264 1000
rect 286 998 294 1000
rect 316 998 324 1000
rect 346 998 354 1000
rect 376 998 384 1000
rect 406 998 414 1000
rect 436 998 444 1000
rect 466 998 474 1000
rect 496 998 504 1000
rect 526 998 534 1000
rect 46 990 54 998
rect 66 990 84 998
rect 96 990 114 998
rect 126 990 144 998
rect 156 990 174 998
rect 186 990 204 998
rect 216 990 234 998
rect 246 990 264 998
rect 276 990 294 998
rect 306 990 324 998
rect 336 990 354 998
rect 366 990 384 998
rect 396 990 414 998
rect 426 990 444 998
rect 456 990 474 998
rect 486 990 504 998
rect 516 990 534 998
rect 546 990 554 998
rect 76 988 84 990
rect 106 988 114 990
rect 136 988 144 990
rect 166 988 174 990
rect 196 988 204 990
rect 226 988 234 990
rect 256 988 264 990
rect 286 988 294 990
rect 316 988 324 990
rect 346 988 354 990
rect 376 988 384 990
rect 406 988 414 990
rect 436 988 444 990
rect 466 988 474 990
rect 496 988 504 990
rect 526 988 534 990
rect 56 980 64 988
rect 76 980 94 988
rect 106 980 124 988
rect 136 980 154 988
rect 166 980 184 988
rect 196 980 214 988
rect 226 980 244 988
rect 256 980 274 988
rect 286 980 304 988
rect 316 980 334 988
rect 346 980 364 988
rect 376 980 394 988
rect 406 980 424 988
rect 436 980 454 988
rect 466 980 484 988
rect 496 980 514 988
rect 526 980 544 988
rect 76 978 84 980
rect 106 978 114 980
rect 136 978 144 980
rect 166 978 174 980
rect 196 978 204 980
rect 226 978 234 980
rect 256 978 264 980
rect 286 978 294 980
rect 316 978 324 980
rect 346 978 354 980
rect 376 978 384 980
rect 406 978 414 980
rect 436 978 444 980
rect 466 978 474 980
rect 496 978 504 980
rect 526 978 534 980
rect 46 970 54 978
rect 66 970 84 978
rect 96 970 114 978
rect 126 970 144 978
rect 156 970 174 978
rect 186 970 204 978
rect 216 970 234 978
rect 246 970 264 978
rect 276 970 294 978
rect 306 970 324 978
rect 336 970 354 978
rect 366 970 384 978
rect 396 970 414 978
rect 426 970 444 978
rect 456 970 474 978
rect 486 970 504 978
rect 516 970 534 978
rect 546 970 554 978
rect 536 960 544 968
rect 46 950 54 958
rect 66 950 84 958
rect 96 950 114 958
rect 126 950 144 958
rect 156 950 174 958
rect 186 950 204 958
rect 216 950 234 958
rect 246 950 264 958
rect 276 950 294 958
rect 306 950 324 958
rect 336 950 354 958
rect 366 950 384 958
rect 396 950 414 958
rect 426 950 444 958
rect 456 950 474 958
rect 486 950 504 958
rect 516 950 534 958
rect 546 950 554 958
rect 76 948 84 950
rect 106 948 114 950
rect 136 948 144 950
rect 166 948 174 950
rect 196 948 204 950
rect 226 948 234 950
rect 256 948 264 950
rect 286 948 294 950
rect 316 948 324 950
rect 346 948 354 950
rect 376 948 384 950
rect 406 948 414 950
rect 436 948 444 950
rect 466 948 474 950
rect 496 948 504 950
rect 526 948 534 950
rect 56 940 64 948
rect 76 940 94 948
rect 106 940 124 948
rect 136 940 154 948
rect 166 940 184 948
rect 196 940 214 948
rect 226 940 244 948
rect 256 940 274 948
rect 286 940 304 948
rect 316 940 334 948
rect 346 940 364 948
rect 376 940 394 948
rect 406 940 424 948
rect 436 940 454 948
rect 466 940 484 948
rect 496 940 514 948
rect 526 940 544 948
rect 76 938 84 940
rect 106 938 114 940
rect 136 938 144 940
rect 166 938 174 940
rect 196 938 204 940
rect 226 938 234 940
rect 256 938 264 940
rect 286 938 294 940
rect 316 938 324 940
rect 346 938 354 940
rect 376 938 384 940
rect 406 938 414 940
rect 436 938 444 940
rect 466 938 474 940
rect 496 938 504 940
rect 526 938 534 940
rect 46 930 54 938
rect 66 930 84 938
rect 96 930 114 938
rect 126 930 144 938
rect 156 930 174 938
rect 186 930 204 938
rect 216 930 234 938
rect 246 930 264 938
rect 276 930 294 938
rect 306 930 324 938
rect 336 930 354 938
rect 366 930 384 938
rect 396 930 414 938
rect 426 930 444 938
rect 456 930 474 938
rect 486 930 504 938
rect 516 930 534 938
rect 546 930 554 938
rect 76 928 84 930
rect 106 928 114 930
rect 136 928 144 930
rect 166 928 174 930
rect 196 928 204 930
rect 226 928 234 930
rect 256 928 264 930
rect 286 928 294 930
rect 316 928 324 930
rect 346 928 354 930
rect 376 928 384 930
rect 406 928 414 930
rect 436 928 444 930
rect 466 928 474 930
rect 496 928 504 930
rect 526 928 534 930
rect 56 920 64 928
rect 76 920 94 928
rect 106 920 124 928
rect 136 920 154 928
rect 166 920 184 928
rect 196 920 214 928
rect 226 920 244 928
rect 256 920 274 928
rect 286 920 304 928
rect 316 920 334 928
rect 346 920 364 928
rect 376 920 394 928
rect 406 920 424 928
rect 436 920 454 928
rect 466 920 484 928
rect 496 920 514 928
rect 526 920 544 928
rect 76 918 84 920
rect 106 918 114 920
rect 136 918 144 920
rect 166 918 174 920
rect 196 918 204 920
rect 226 918 234 920
rect 256 918 264 920
rect 286 918 294 920
rect 316 918 324 920
rect 346 918 354 920
rect 376 918 384 920
rect 406 918 414 920
rect 436 918 444 920
rect 466 918 474 920
rect 496 918 504 920
rect 526 918 534 920
rect 46 910 54 918
rect 66 910 84 918
rect 96 910 114 918
rect 126 910 144 918
rect 156 910 174 918
rect 186 910 204 918
rect 216 910 234 918
rect 246 910 264 918
rect 276 910 294 918
rect 306 910 324 918
rect 336 910 354 918
rect 366 910 384 918
rect 396 910 414 918
rect 426 910 444 918
rect 456 910 474 918
rect 486 910 504 918
rect 516 910 534 918
rect 546 910 554 918
rect 76 908 84 910
rect 106 908 114 910
rect 136 908 144 910
rect 166 908 174 910
rect 196 908 204 910
rect 226 908 234 910
rect 256 908 264 910
rect 286 908 294 910
rect 316 908 324 910
rect 346 908 354 910
rect 376 908 384 910
rect 406 908 414 910
rect 436 908 444 910
rect 466 908 474 910
rect 496 908 504 910
rect 526 908 534 910
rect 56 900 64 908
rect 76 900 94 908
rect 106 900 124 908
rect 136 900 154 908
rect 166 900 184 908
rect 196 900 214 908
rect 226 900 244 908
rect 256 900 274 908
rect 286 900 304 908
rect 316 900 334 908
rect 346 900 364 908
rect 376 900 394 908
rect 406 900 424 908
rect 436 900 454 908
rect 466 900 484 908
rect 496 900 514 908
rect 526 900 544 908
rect 76 898 84 900
rect 106 898 114 900
rect 136 898 144 900
rect 166 898 174 900
rect 196 898 204 900
rect 226 898 234 900
rect 256 898 264 900
rect 286 898 294 900
rect 316 898 324 900
rect 346 898 354 900
rect 376 898 384 900
rect 406 898 414 900
rect 436 898 444 900
rect 466 898 474 900
rect 496 898 504 900
rect 526 898 534 900
rect 46 890 54 898
rect 66 890 84 898
rect 96 890 114 898
rect 126 890 144 898
rect 156 890 174 898
rect 186 890 204 898
rect 216 890 234 898
rect 246 890 264 898
rect 276 890 294 898
rect 306 890 324 898
rect 336 890 354 898
rect 366 890 384 898
rect 396 890 414 898
rect 426 890 444 898
rect 456 890 474 898
rect 486 890 504 898
rect 516 890 534 898
rect 546 890 554 898
rect 76 888 84 890
rect 106 888 114 890
rect 136 888 144 890
rect 166 888 174 890
rect 196 888 204 890
rect 226 888 234 890
rect 256 888 264 890
rect 286 888 294 890
rect 316 888 324 890
rect 346 888 354 890
rect 376 888 384 890
rect 406 888 414 890
rect 436 888 444 890
rect 466 888 474 890
rect 496 888 504 890
rect 526 888 534 890
rect 56 878 64 888
rect 76 878 94 888
rect 106 878 124 888
rect 136 878 154 888
rect 166 878 184 888
rect 196 878 214 888
rect 226 878 244 888
rect 256 878 274 888
rect 286 878 304 888
rect 316 878 334 888
rect 346 878 364 888
rect 376 878 394 888
rect 406 878 424 888
rect 436 878 454 888
rect 466 878 484 888
rect 496 878 514 888
rect 526 878 544 888
rect 46 870 554 878
rect 4 644 12 652
rect 24 644 42 652
rect 54 644 72 652
rect 84 644 102 652
rect 114 644 132 652
rect 144 644 162 652
rect 174 644 192 652
rect 204 644 222 652
rect 234 644 242 652
rect 256 644 264 652
rect 276 644 294 652
rect 306 644 324 652
rect 336 644 344 652
rect 358 644 366 652
rect 378 644 396 652
rect 408 644 426 652
rect 438 644 456 652
rect 468 644 486 652
rect 498 644 516 652
rect 528 644 546 652
rect 558 644 576 652
rect 588 644 596 652
rect 34 642 42 644
rect 64 642 72 644
rect 94 642 102 644
rect 124 642 132 644
rect 154 642 162 644
rect 184 642 192 644
rect 214 642 222 644
rect 286 642 294 644
rect 316 642 324 644
rect 378 642 386 644
rect 408 642 416 644
rect 438 642 446 644
rect 468 642 476 644
rect 498 642 506 644
rect 528 642 536 644
rect 558 642 566 644
rect 14 634 22 642
rect 34 634 52 642
rect 64 634 82 642
rect 94 634 112 642
rect 124 634 142 642
rect 154 634 172 642
rect 184 634 202 642
rect 214 634 232 642
rect 244 634 252 642
rect 266 634 274 642
rect 286 634 304 642
rect 316 634 334 642
rect 348 634 356 642
rect 368 634 386 642
rect 398 634 416 642
rect 428 634 446 642
rect 458 634 476 642
rect 488 634 506 642
rect 518 634 536 642
rect 548 634 566 642
rect 578 634 586 642
rect 34 632 42 634
rect 64 632 72 634
rect 94 632 102 634
rect 124 632 132 634
rect 154 632 162 634
rect 184 632 192 634
rect 214 632 222 634
rect 286 632 294 634
rect 316 632 324 634
rect 378 632 386 634
rect 408 632 416 634
rect 438 632 446 634
rect 468 632 476 634
rect 498 632 506 634
rect 528 632 536 634
rect 558 632 566 634
rect 4 624 12 632
rect 24 624 42 632
rect 54 624 72 632
rect 84 624 102 632
rect 114 624 132 632
rect 144 624 162 632
rect 174 624 192 632
rect 204 624 222 632
rect 234 624 242 632
rect 256 624 264 632
rect 276 624 294 632
rect 306 624 324 632
rect 336 624 344 632
rect 358 624 366 632
rect 378 624 396 632
rect 408 624 426 632
rect 438 624 456 632
rect 468 624 486 632
rect 498 624 516 632
rect 528 624 546 632
rect 558 624 576 632
rect 588 624 596 632
rect 34 622 42 624
rect 64 622 72 624
rect 94 622 102 624
rect 124 622 132 624
rect 154 622 162 624
rect 184 622 192 624
rect 214 622 222 624
rect 286 622 294 624
rect 316 622 324 624
rect 378 622 386 624
rect 408 622 416 624
rect 438 622 446 624
rect 468 622 476 624
rect 498 622 506 624
rect 528 622 536 624
rect 558 622 566 624
rect 14 614 22 622
rect 34 614 52 622
rect 64 614 82 622
rect 94 614 112 622
rect 124 614 142 622
rect 154 614 172 622
rect 184 614 202 622
rect 214 614 232 622
rect 244 614 252 622
rect 266 614 274 622
rect 286 614 304 622
rect 316 614 334 622
rect 348 614 356 622
rect 368 614 386 622
rect 398 614 416 622
rect 428 614 446 622
rect 458 614 476 622
rect 488 614 506 622
rect 518 614 536 622
rect 548 614 566 622
rect 578 614 586 622
rect 4 604 12 612
rect 24 604 32 612
rect 214 602 222 614
rect 286 612 294 614
rect 316 612 324 614
rect 234 604 242 612
rect 256 604 264 612
rect 276 604 294 612
rect 306 604 324 612
rect 336 604 344 612
rect 358 604 366 612
rect 286 602 294 604
rect 316 602 324 604
rect 378 602 386 614
rect 568 604 576 612
rect 588 604 596 612
rect 14 594 22 602
rect 34 594 52 602
rect 64 594 82 602
rect 94 594 112 602
rect 124 594 142 602
rect 154 594 172 602
rect 184 594 202 602
rect 214 594 232 602
rect 244 594 252 602
rect 34 592 42 594
rect 64 592 72 594
rect 94 592 102 594
rect 124 592 132 594
rect 154 592 162 594
rect 184 592 192 594
rect 214 592 222 594
rect 266 592 274 602
rect 286 592 304 602
rect 316 592 334 602
rect 348 594 356 602
rect 368 594 386 602
rect 398 594 416 602
rect 428 594 446 602
rect 458 594 476 602
rect 488 594 506 602
rect 518 594 536 602
rect 548 594 566 602
rect 578 594 586 602
rect 378 592 386 594
rect 408 592 416 594
rect 438 592 446 594
rect 468 592 476 594
rect 498 592 506 594
rect 528 592 536 594
rect 558 592 566 594
rect 4 584 12 592
rect 24 584 42 592
rect 54 584 72 592
rect 84 584 102 592
rect 34 582 42 584
rect 64 582 72 584
rect 94 582 102 584
rect 114 582 132 592
rect 144 582 162 592
rect 174 582 192 592
rect 204 582 222 592
rect 234 582 242 592
rect 14 574 22 582
rect 34 574 52 582
rect 64 574 82 582
rect 94 574 252 582
rect 256 574 344 592
rect 358 582 366 592
rect 378 582 396 592
rect 408 582 426 592
rect 438 582 456 592
rect 468 582 486 592
rect 498 584 516 592
rect 528 584 546 592
rect 558 584 576 592
rect 588 584 596 592
rect 498 582 506 584
rect 528 582 536 584
rect 558 582 566 584
rect 348 574 506 582
rect 518 574 536 582
rect 548 574 566 582
rect 578 574 586 582
rect 34 572 42 574
rect 64 572 72 574
rect 94 572 102 574
rect 4 564 12 572
rect 24 564 42 572
rect 54 564 72 572
rect 84 564 102 572
rect 114 564 132 574
rect 144 564 162 574
rect 174 564 192 574
rect 204 564 222 574
rect 234 564 242 574
rect 256 564 264 574
rect 276 564 294 574
rect 306 564 324 574
rect 336 564 344 574
rect 358 564 366 574
rect 378 564 396 574
rect 408 564 426 574
rect 438 564 456 574
rect 468 564 486 574
rect 498 572 506 574
rect 528 572 536 574
rect 558 572 566 574
rect 498 564 516 572
rect 528 564 546 572
rect 558 564 576 572
rect 588 564 596 572
rect 34 562 42 564
rect 64 562 72 564
rect 94 562 102 564
rect 124 562 132 564
rect 154 562 162 564
rect 184 562 192 564
rect 214 562 222 564
rect 286 562 294 564
rect 316 562 324 564
rect 378 562 386 564
rect 408 562 416 564
rect 438 562 446 564
rect 468 562 476 564
rect 498 562 506 564
rect 528 562 536 564
rect 558 562 566 564
rect 14 554 22 562
rect 34 554 52 562
rect 64 554 82 562
rect 94 554 112 562
rect 124 554 142 562
rect 154 554 172 562
rect 184 554 202 562
rect 214 554 232 562
rect 244 554 252 562
rect 266 554 274 562
rect 286 554 304 562
rect 316 554 334 562
rect 348 554 356 562
rect 368 554 386 562
rect 398 554 416 562
rect 428 554 446 562
rect 458 554 476 562
rect 488 554 506 562
rect 518 554 536 562
rect 548 554 566 562
rect 578 554 586 562
rect 34 552 42 554
rect 64 552 72 554
rect 94 552 102 554
rect 124 552 132 554
rect 154 552 162 554
rect 184 552 192 554
rect 214 552 222 554
rect 286 552 294 554
rect 316 552 324 554
rect 378 552 386 554
rect 408 552 416 554
rect 438 552 446 554
rect 468 552 476 554
rect 498 552 506 554
rect 528 552 536 554
rect 558 552 566 554
rect 4 544 12 552
rect 24 544 42 552
rect 54 544 72 552
rect 84 544 102 552
rect 114 544 132 552
rect 144 544 162 552
rect 174 544 192 552
rect 204 544 222 552
rect 234 544 242 552
rect 256 544 264 552
rect 276 544 294 552
rect 306 544 324 552
rect 336 544 344 552
rect 358 544 366 552
rect 378 544 396 552
rect 408 544 426 552
rect 438 544 456 552
rect 468 544 486 552
rect 498 544 516 552
rect 528 544 546 552
rect 558 544 576 552
rect 588 544 596 552
rect 34 542 42 544
rect 64 542 72 544
rect 94 542 102 544
rect 124 542 132 544
rect 154 542 162 544
rect 184 542 192 544
rect 214 542 222 544
rect 286 542 294 544
rect 316 542 324 544
rect 378 542 386 544
rect 408 542 416 544
rect 438 542 446 544
rect 468 542 476 544
rect 498 542 506 544
rect 528 542 536 544
rect 558 542 566 544
rect 14 534 22 542
rect 34 534 52 542
rect 64 534 82 542
rect 94 534 112 542
rect 124 534 142 542
rect 154 534 172 542
rect 184 534 202 542
rect 214 534 232 542
rect 244 534 252 542
rect 266 534 274 542
rect 286 534 304 542
rect 316 534 334 542
rect 348 534 356 542
rect 368 534 386 542
rect 398 534 416 542
rect 428 534 446 542
rect 458 534 476 542
rect 488 534 506 542
rect 518 534 536 542
rect 548 534 566 542
rect 578 534 586 542
rect 34 532 42 534
rect 64 532 72 534
rect 94 532 102 534
rect 124 532 132 534
rect 154 532 162 534
rect 184 532 192 534
rect 214 532 222 534
rect 286 532 294 534
rect 316 532 324 534
rect 378 532 386 534
rect 408 532 416 534
rect 438 532 446 534
rect 468 532 476 534
rect 498 532 506 534
rect 528 532 536 534
rect 558 532 566 534
rect 4 524 12 532
rect 24 524 42 532
rect 54 524 72 532
rect 84 524 102 532
rect 114 524 132 532
rect 144 524 162 532
rect 174 524 192 532
rect 204 524 222 532
rect 234 524 242 532
rect 256 524 264 532
rect 276 524 294 532
rect 306 524 324 532
rect 336 524 344 532
rect 358 524 366 532
rect 378 524 396 532
rect 408 524 426 532
rect 438 524 456 532
rect 468 524 486 532
rect 498 524 516 532
rect 528 524 546 532
rect 558 524 576 532
rect 588 524 596 532
rect 4 12 12 516
rect 24 508 32 516
rect 44 508 52 516
rect 64 508 72 516
rect 84 508 92 516
rect 104 508 112 516
rect 124 508 132 516
rect 144 508 152 516
rect 164 508 172 516
rect 184 508 192 516
rect 204 508 212 516
rect 224 508 232 516
rect 244 508 252 516
rect 264 508 272 516
rect 284 508 292 516
rect 318 508 326 516
rect 338 508 346 516
rect 358 508 366 516
rect 378 508 386 516
rect 398 508 406 516
rect 418 508 426 516
rect 438 508 446 516
rect 458 508 466 516
rect 478 508 486 516
rect 498 508 506 516
rect 518 508 526 516
rect 538 508 546 516
rect 558 508 566 516
rect 578 508 596 516
rect 588 12 596 508
rect 4 8 182 12
rect 14 4 182 8
rect 408 8 596 12
rect 408 4 586 8
<< polysilicon >>
rect 62 432 76 436
rect 62 84 64 432
rect 72 430 76 432
rect 276 430 280 436
rect 72 346 74 430
rect 320 430 324 436
rect 524 432 538 436
rect 524 430 528 432
rect 72 340 76 346
rect 276 340 280 346
rect 72 304 74 340
rect 72 298 76 304
rect 276 298 280 304
rect 72 216 74 298
rect 526 346 528 430
rect 320 340 324 346
rect 524 340 528 346
rect 526 304 528 340
rect 320 298 324 304
rect 524 298 528 304
rect 72 210 76 216
rect 276 210 280 216
rect 72 174 74 210
rect 72 168 76 174
rect 276 168 280 174
rect 72 86 74 168
rect 526 216 528 298
rect 320 210 324 216
rect 524 210 528 216
rect 526 174 528 210
rect 320 168 324 174
rect 524 168 528 174
rect 72 84 76 86
rect 62 80 76 84
rect 276 80 280 86
rect 526 86 528 168
rect 320 80 324 86
rect 524 84 528 86
rect 536 84 538 432
rect 524 80 538 84
<< polycontact >>
rect 64 84 72 432
rect 528 84 536 432
<< metal1 >>
rect 124 1460 476 1480
rect 144 1440 456 1460
rect 164 1420 436 1440
rect 184 1400 416 1420
rect 0 1338 198 1340
rect 0 840 2 1338
rect 190 1320 198 1338
rect 20 1319 198 1320
rect 20 840 21 1319
rect 204 1300 396 1400
rect 402 1338 600 1340
rect 402 1320 408 1338
rect 576 1320 580 1338
rect 402 1319 580 1320
rect 100 1298 560 1300
rect 42 1290 46 1298
rect 54 1290 56 1298
rect 64 1290 66 1298
rect 84 1290 86 1298
rect 94 1290 96 1298
rect 114 1290 116 1298
rect 124 1290 126 1298
rect 144 1290 146 1298
rect 154 1290 156 1298
rect 174 1290 176 1298
rect 184 1290 186 1298
rect 204 1290 206 1298
rect 214 1290 216 1298
rect 234 1290 236 1298
rect 244 1290 246 1298
rect 264 1290 266 1298
rect 274 1290 276 1298
rect 294 1290 296 1298
rect 304 1290 306 1298
rect 324 1290 326 1298
rect 334 1290 336 1298
rect 354 1290 356 1298
rect 364 1290 366 1298
rect 384 1290 386 1298
rect 394 1290 396 1298
rect 414 1290 416 1298
rect 424 1290 426 1298
rect 444 1290 446 1298
rect 454 1290 456 1298
rect 474 1290 476 1298
rect 484 1290 486 1298
rect 504 1290 506 1298
rect 514 1290 516 1298
rect 534 1290 536 1298
rect 544 1290 546 1298
rect 554 1290 560 1298
rect 42 1288 76 1290
rect 84 1288 106 1290
rect 114 1288 136 1290
rect 144 1288 166 1290
rect 174 1288 196 1290
rect 204 1288 226 1290
rect 234 1288 256 1290
rect 264 1288 286 1290
rect 294 1288 316 1290
rect 324 1288 346 1290
rect 354 1288 376 1290
rect 384 1288 406 1290
rect 414 1288 436 1290
rect 444 1288 466 1290
rect 474 1288 496 1290
rect 504 1288 526 1290
rect 534 1288 560 1290
rect 42 1280 46 1288
rect 54 1280 56 1288
rect 64 1280 66 1288
rect 74 1280 76 1288
rect 94 1280 96 1288
rect 104 1280 106 1288
rect 124 1280 126 1288
rect 134 1280 136 1288
rect 154 1280 156 1288
rect 164 1280 166 1288
rect 184 1280 186 1288
rect 194 1280 196 1288
rect 214 1280 216 1288
rect 224 1280 226 1288
rect 244 1280 246 1288
rect 254 1280 256 1288
rect 274 1280 276 1288
rect 284 1280 286 1288
rect 304 1280 306 1288
rect 314 1280 316 1288
rect 334 1280 336 1288
rect 344 1280 346 1288
rect 364 1280 366 1288
rect 374 1280 376 1288
rect 394 1280 396 1288
rect 404 1280 406 1288
rect 424 1280 426 1288
rect 434 1280 436 1288
rect 454 1280 456 1288
rect 464 1280 466 1288
rect 484 1280 486 1288
rect 494 1280 496 1288
rect 514 1280 516 1288
rect 524 1280 526 1288
rect 544 1280 546 1288
rect 554 1280 560 1288
rect 42 1278 76 1280
rect 84 1278 106 1280
rect 114 1278 136 1280
rect 144 1278 166 1280
rect 174 1278 196 1280
rect 204 1278 226 1280
rect 234 1278 256 1280
rect 264 1278 286 1280
rect 294 1278 316 1280
rect 324 1278 346 1280
rect 354 1278 376 1280
rect 384 1278 406 1280
rect 414 1278 436 1280
rect 444 1278 466 1280
rect 474 1278 496 1280
rect 504 1278 526 1280
rect 534 1278 560 1280
rect 42 1270 46 1278
rect 54 1270 56 1278
rect 64 1270 66 1278
rect 84 1270 86 1278
rect 94 1270 96 1278
rect 114 1270 116 1278
rect 124 1270 126 1278
rect 144 1270 146 1278
rect 154 1270 156 1278
rect 174 1270 176 1278
rect 184 1270 186 1278
rect 204 1270 206 1278
rect 214 1270 216 1278
rect 234 1270 236 1278
rect 244 1270 246 1278
rect 264 1270 266 1278
rect 274 1270 276 1278
rect 294 1270 296 1278
rect 304 1270 306 1278
rect 324 1270 326 1278
rect 334 1270 336 1278
rect 354 1270 356 1278
rect 364 1270 366 1278
rect 384 1270 386 1278
rect 394 1270 396 1278
rect 414 1270 416 1278
rect 424 1270 426 1278
rect 444 1270 446 1278
rect 454 1270 456 1278
rect 474 1270 476 1278
rect 484 1270 486 1278
rect 504 1270 506 1278
rect 514 1270 516 1278
rect 534 1270 536 1278
rect 544 1270 546 1278
rect 554 1270 560 1278
rect 42 1268 76 1270
rect 84 1268 106 1270
rect 114 1268 136 1270
rect 144 1268 166 1270
rect 174 1268 196 1270
rect 204 1268 226 1270
rect 234 1268 256 1270
rect 264 1268 286 1270
rect 294 1268 316 1270
rect 324 1268 346 1270
rect 354 1268 376 1270
rect 384 1268 406 1270
rect 414 1268 436 1270
rect 444 1268 466 1270
rect 474 1268 496 1270
rect 504 1268 526 1270
rect 534 1268 560 1270
rect 42 1260 46 1268
rect 54 1260 56 1268
rect 64 1260 66 1268
rect 74 1260 76 1268
rect 94 1260 96 1268
rect 104 1260 106 1268
rect 124 1260 126 1268
rect 134 1260 136 1268
rect 154 1260 156 1268
rect 164 1260 166 1268
rect 184 1260 186 1268
rect 194 1260 196 1268
rect 214 1260 216 1268
rect 224 1260 226 1268
rect 244 1260 246 1268
rect 254 1260 256 1268
rect 274 1260 276 1268
rect 284 1260 286 1268
rect 304 1260 306 1268
rect 314 1260 316 1268
rect 334 1260 336 1268
rect 344 1260 346 1268
rect 364 1260 366 1268
rect 374 1260 376 1268
rect 394 1260 396 1268
rect 404 1260 406 1268
rect 424 1260 426 1268
rect 434 1260 436 1268
rect 454 1260 456 1268
rect 464 1260 466 1268
rect 484 1260 486 1268
rect 494 1260 496 1268
rect 514 1260 516 1268
rect 524 1260 526 1268
rect 544 1260 546 1268
rect 554 1260 560 1268
rect 42 1258 76 1260
rect 84 1258 106 1260
rect 114 1258 136 1260
rect 144 1258 166 1260
rect 174 1258 196 1260
rect 204 1258 226 1260
rect 234 1258 256 1260
rect 264 1258 286 1260
rect 294 1258 316 1260
rect 324 1258 346 1260
rect 354 1258 376 1260
rect 384 1258 406 1260
rect 414 1258 436 1260
rect 444 1258 466 1260
rect 474 1258 496 1260
rect 504 1258 526 1260
rect 534 1258 560 1260
rect 42 1250 46 1258
rect 54 1250 56 1258
rect 64 1250 66 1258
rect 84 1250 86 1258
rect 94 1250 96 1258
rect 114 1250 116 1258
rect 124 1250 126 1258
rect 144 1250 146 1258
rect 154 1250 156 1258
rect 174 1250 176 1258
rect 184 1250 186 1258
rect 204 1250 206 1258
rect 214 1250 216 1258
rect 234 1250 236 1258
rect 244 1250 246 1258
rect 264 1250 266 1258
rect 274 1250 276 1258
rect 294 1250 296 1258
rect 304 1250 306 1258
rect 324 1250 326 1258
rect 334 1250 336 1258
rect 354 1250 356 1258
rect 364 1250 366 1258
rect 384 1250 386 1258
rect 394 1250 396 1258
rect 414 1250 416 1258
rect 424 1250 426 1258
rect 444 1250 446 1258
rect 454 1250 456 1258
rect 474 1250 476 1258
rect 484 1250 486 1258
rect 504 1250 506 1258
rect 514 1250 516 1258
rect 534 1250 536 1258
rect 544 1250 546 1258
rect 554 1250 560 1258
rect 42 1248 76 1250
rect 84 1248 106 1250
rect 114 1248 136 1250
rect 144 1248 166 1250
rect 174 1248 196 1250
rect 204 1248 226 1250
rect 234 1248 256 1250
rect 264 1248 286 1250
rect 294 1248 316 1250
rect 324 1248 346 1250
rect 354 1248 376 1250
rect 384 1248 406 1250
rect 414 1248 436 1250
rect 444 1248 466 1250
rect 474 1248 496 1250
rect 504 1248 526 1250
rect 534 1248 560 1250
rect 42 1240 46 1248
rect 54 1240 56 1248
rect 64 1240 66 1248
rect 74 1240 76 1248
rect 94 1240 96 1248
rect 104 1240 106 1248
rect 124 1240 126 1248
rect 134 1240 136 1248
rect 154 1240 156 1248
rect 164 1240 166 1248
rect 184 1240 186 1248
rect 194 1240 196 1248
rect 214 1240 216 1248
rect 224 1240 226 1248
rect 244 1240 246 1248
rect 254 1240 256 1248
rect 274 1240 276 1248
rect 284 1240 286 1248
rect 304 1240 306 1248
rect 314 1240 316 1248
rect 334 1240 336 1248
rect 344 1240 346 1248
rect 364 1240 366 1248
rect 374 1240 376 1248
rect 394 1240 396 1248
rect 404 1240 406 1248
rect 424 1240 426 1248
rect 434 1240 436 1248
rect 454 1240 456 1248
rect 464 1240 466 1248
rect 484 1240 486 1248
rect 494 1240 496 1248
rect 514 1240 516 1248
rect 524 1240 526 1248
rect 544 1240 546 1248
rect 554 1240 560 1248
rect 42 1238 76 1240
rect 84 1238 106 1240
rect 114 1238 136 1240
rect 144 1238 166 1240
rect 174 1238 196 1240
rect 204 1238 226 1240
rect 234 1238 256 1240
rect 264 1238 286 1240
rect 294 1238 316 1240
rect 324 1238 346 1240
rect 354 1238 376 1240
rect 384 1238 406 1240
rect 414 1238 436 1240
rect 444 1238 466 1240
rect 474 1238 496 1240
rect 504 1238 526 1240
rect 534 1238 560 1240
rect 42 1230 46 1238
rect 54 1230 56 1238
rect 64 1230 66 1238
rect 84 1230 86 1238
rect 94 1230 96 1238
rect 114 1230 116 1238
rect 124 1230 126 1238
rect 144 1230 146 1238
rect 154 1230 156 1238
rect 174 1230 176 1238
rect 184 1230 186 1238
rect 204 1230 206 1238
rect 214 1230 216 1238
rect 234 1230 236 1238
rect 244 1230 246 1238
rect 264 1230 266 1238
rect 274 1230 276 1238
rect 294 1230 296 1238
rect 304 1230 306 1238
rect 324 1230 326 1238
rect 334 1230 336 1238
rect 354 1230 356 1238
rect 364 1230 366 1238
rect 384 1230 386 1238
rect 394 1230 396 1238
rect 414 1230 416 1238
rect 424 1230 426 1238
rect 444 1230 446 1238
rect 454 1230 456 1238
rect 474 1230 476 1238
rect 484 1230 486 1238
rect 504 1230 506 1238
rect 514 1230 516 1238
rect 534 1230 536 1238
rect 544 1230 546 1238
rect 554 1230 560 1238
rect 42 1228 76 1230
rect 84 1228 106 1230
rect 114 1228 136 1230
rect 144 1228 166 1230
rect 174 1228 196 1230
rect 204 1228 226 1230
rect 234 1228 256 1230
rect 264 1228 286 1230
rect 294 1228 316 1230
rect 324 1228 346 1230
rect 354 1228 376 1230
rect 384 1228 406 1230
rect 414 1228 436 1230
rect 444 1228 466 1230
rect 474 1228 496 1230
rect 504 1228 526 1230
rect 534 1228 560 1230
rect 42 1220 46 1228
rect 54 1220 56 1228
rect 64 1220 66 1228
rect 74 1220 76 1228
rect 94 1220 96 1228
rect 104 1220 106 1228
rect 124 1220 126 1228
rect 134 1220 136 1228
rect 154 1220 156 1228
rect 164 1220 166 1228
rect 184 1220 186 1228
rect 194 1220 196 1228
rect 214 1220 216 1228
rect 224 1220 226 1228
rect 244 1220 246 1228
rect 254 1220 256 1228
rect 274 1220 276 1228
rect 284 1220 286 1228
rect 304 1220 306 1228
rect 314 1220 316 1228
rect 334 1220 336 1228
rect 344 1220 346 1228
rect 364 1220 366 1228
rect 374 1220 376 1228
rect 394 1220 396 1228
rect 404 1220 406 1228
rect 424 1220 426 1228
rect 434 1220 436 1228
rect 454 1220 456 1228
rect 464 1220 466 1228
rect 484 1220 486 1228
rect 494 1220 496 1228
rect 514 1220 516 1228
rect 524 1220 526 1228
rect 544 1220 546 1228
rect 554 1220 560 1228
rect 42 1218 76 1220
rect 84 1218 106 1220
rect 114 1218 136 1220
rect 144 1218 166 1220
rect 174 1218 196 1220
rect 204 1218 226 1220
rect 234 1218 256 1220
rect 264 1218 286 1220
rect 294 1218 316 1220
rect 324 1218 346 1220
rect 354 1218 376 1220
rect 384 1218 406 1220
rect 414 1218 436 1220
rect 444 1218 466 1220
rect 474 1218 496 1220
rect 504 1218 526 1220
rect 534 1218 560 1220
rect 42 1210 46 1218
rect 54 1210 56 1218
rect 64 1210 66 1218
rect 84 1210 86 1218
rect 94 1210 96 1218
rect 114 1210 116 1218
rect 124 1210 126 1218
rect 144 1210 146 1218
rect 154 1210 156 1218
rect 174 1210 176 1218
rect 184 1210 186 1218
rect 204 1210 206 1218
rect 214 1210 216 1218
rect 234 1210 236 1218
rect 244 1210 246 1218
rect 264 1210 266 1218
rect 274 1210 276 1218
rect 294 1210 296 1218
rect 304 1210 306 1218
rect 324 1210 326 1218
rect 334 1210 336 1218
rect 354 1210 356 1218
rect 364 1210 366 1218
rect 384 1210 386 1218
rect 394 1210 396 1218
rect 414 1210 416 1218
rect 424 1210 426 1218
rect 444 1210 446 1218
rect 454 1210 456 1218
rect 474 1210 476 1218
rect 484 1210 486 1218
rect 504 1210 506 1218
rect 514 1210 516 1218
rect 534 1210 536 1218
rect 544 1210 546 1218
rect 554 1210 560 1218
rect 42 1208 76 1210
rect 84 1208 106 1210
rect 114 1208 136 1210
rect 144 1208 166 1210
rect 174 1208 196 1210
rect 204 1208 226 1210
rect 234 1208 256 1210
rect 264 1208 286 1210
rect 294 1208 316 1210
rect 324 1208 346 1210
rect 354 1208 376 1210
rect 384 1208 406 1210
rect 414 1208 436 1210
rect 444 1208 466 1210
rect 474 1208 496 1210
rect 504 1208 526 1210
rect 534 1208 560 1210
rect 42 1200 46 1208
rect 54 1200 56 1208
rect 64 1200 66 1208
rect 74 1200 76 1208
rect 94 1200 96 1208
rect 104 1200 106 1208
rect 124 1200 126 1208
rect 134 1200 136 1208
rect 154 1200 156 1208
rect 164 1200 166 1208
rect 184 1200 186 1208
rect 194 1200 196 1208
rect 214 1200 216 1208
rect 224 1200 226 1208
rect 244 1200 246 1208
rect 254 1200 256 1208
rect 274 1200 276 1208
rect 284 1200 286 1208
rect 304 1200 306 1208
rect 314 1200 316 1208
rect 334 1200 336 1208
rect 344 1200 346 1208
rect 364 1200 366 1208
rect 374 1200 376 1208
rect 394 1200 396 1208
rect 404 1200 406 1208
rect 424 1200 426 1208
rect 434 1200 436 1208
rect 454 1200 456 1208
rect 464 1200 466 1208
rect 484 1200 486 1208
rect 494 1200 496 1208
rect 514 1200 516 1208
rect 524 1200 526 1208
rect 544 1200 546 1208
rect 554 1200 560 1208
rect 42 1198 76 1200
rect 84 1198 106 1200
rect 114 1198 136 1200
rect 144 1198 166 1200
rect 174 1198 196 1200
rect 204 1198 226 1200
rect 234 1198 256 1200
rect 264 1198 286 1200
rect 294 1198 316 1200
rect 324 1198 346 1200
rect 354 1198 376 1200
rect 384 1198 406 1200
rect 414 1198 436 1200
rect 444 1198 466 1200
rect 474 1198 496 1200
rect 504 1198 526 1200
rect 534 1198 560 1200
rect 42 1190 46 1198
rect 54 1190 56 1198
rect 64 1190 66 1198
rect 84 1190 86 1198
rect 94 1190 96 1198
rect 114 1190 116 1198
rect 124 1190 126 1198
rect 144 1190 146 1198
rect 154 1190 156 1198
rect 174 1190 176 1198
rect 184 1190 186 1198
rect 204 1190 206 1198
rect 214 1190 216 1198
rect 234 1190 236 1198
rect 244 1190 246 1198
rect 264 1190 266 1198
rect 274 1190 276 1198
rect 294 1190 296 1198
rect 304 1190 306 1198
rect 324 1190 326 1198
rect 334 1190 336 1198
rect 354 1190 356 1198
rect 364 1190 366 1198
rect 384 1190 386 1198
rect 394 1190 396 1198
rect 414 1190 416 1198
rect 424 1190 426 1198
rect 444 1190 446 1198
rect 454 1190 456 1198
rect 474 1190 476 1198
rect 484 1190 486 1198
rect 504 1190 506 1198
rect 514 1190 516 1198
rect 534 1190 536 1198
rect 544 1190 546 1198
rect 554 1190 560 1198
rect 42 1188 76 1190
rect 84 1188 526 1190
rect 534 1188 560 1190
rect 42 1180 46 1188
rect 54 1180 56 1188
rect 64 1180 66 1188
rect 74 1180 76 1188
rect 94 1180 506 1188
rect 514 1180 516 1188
rect 524 1180 526 1188
rect 544 1180 546 1188
rect 554 1180 560 1188
rect 42 1178 76 1180
rect 84 1178 526 1180
rect 534 1178 560 1180
rect 42 1170 46 1178
rect 54 1170 56 1178
rect 64 1170 66 1178
rect 84 1170 86 1178
rect 94 1170 96 1178
rect 114 1170 116 1178
rect 124 1170 126 1178
rect 144 1170 146 1178
rect 154 1170 156 1178
rect 174 1170 176 1178
rect 184 1170 186 1178
rect 204 1170 206 1178
rect 214 1170 216 1178
rect 234 1170 236 1178
rect 244 1170 246 1178
rect 264 1170 266 1178
rect 274 1170 276 1178
rect 294 1170 296 1178
rect 304 1170 306 1178
rect 324 1170 326 1178
rect 334 1170 336 1178
rect 354 1170 356 1178
rect 364 1170 366 1178
rect 384 1170 386 1178
rect 394 1170 396 1178
rect 414 1170 416 1178
rect 424 1170 426 1178
rect 444 1170 446 1178
rect 454 1170 456 1178
rect 474 1170 476 1178
rect 484 1170 486 1178
rect 504 1170 506 1178
rect 514 1170 516 1178
rect 534 1170 536 1178
rect 544 1170 546 1178
rect 554 1170 560 1178
rect 42 1168 76 1170
rect 84 1168 106 1170
rect 114 1168 136 1170
rect 144 1168 166 1170
rect 174 1168 196 1170
rect 204 1168 226 1170
rect 234 1168 256 1170
rect 264 1168 286 1170
rect 294 1168 316 1170
rect 324 1168 346 1170
rect 354 1168 376 1170
rect 384 1168 406 1170
rect 414 1168 436 1170
rect 444 1168 466 1170
rect 474 1168 496 1170
rect 504 1168 526 1170
rect 534 1168 560 1170
rect 42 1160 46 1168
rect 54 1160 56 1168
rect 64 1160 66 1168
rect 74 1160 76 1168
rect 94 1160 96 1168
rect 104 1160 106 1168
rect 124 1160 126 1168
rect 134 1160 136 1168
rect 154 1160 156 1168
rect 164 1160 166 1168
rect 184 1160 186 1168
rect 194 1160 196 1168
rect 214 1160 216 1168
rect 224 1160 226 1168
rect 244 1160 246 1168
rect 254 1160 256 1168
rect 274 1160 276 1168
rect 284 1160 286 1168
rect 304 1160 306 1168
rect 314 1160 316 1168
rect 334 1160 336 1168
rect 344 1160 346 1168
rect 364 1160 366 1168
rect 374 1160 376 1168
rect 394 1160 396 1168
rect 404 1160 406 1168
rect 424 1160 426 1168
rect 434 1160 436 1168
rect 454 1160 456 1168
rect 464 1160 466 1168
rect 484 1160 486 1168
rect 494 1160 496 1168
rect 514 1160 516 1168
rect 524 1160 526 1168
rect 544 1160 546 1168
rect 554 1160 560 1168
rect 42 1158 76 1160
rect 84 1158 106 1160
rect 114 1158 136 1160
rect 144 1158 166 1160
rect 174 1158 196 1160
rect 204 1158 226 1160
rect 234 1158 256 1160
rect 264 1158 286 1160
rect 294 1158 316 1160
rect 324 1158 346 1160
rect 354 1158 376 1160
rect 384 1158 406 1160
rect 414 1158 436 1160
rect 444 1158 466 1160
rect 474 1158 496 1160
rect 504 1158 526 1160
rect 534 1158 560 1160
rect 42 1150 46 1158
rect 54 1150 56 1158
rect 64 1150 66 1158
rect 84 1150 86 1158
rect 94 1150 96 1158
rect 114 1150 116 1158
rect 124 1150 126 1158
rect 144 1150 146 1158
rect 154 1150 156 1158
rect 174 1150 176 1158
rect 184 1150 186 1158
rect 204 1150 206 1158
rect 214 1150 216 1158
rect 234 1150 236 1158
rect 244 1150 246 1158
rect 264 1150 266 1158
rect 274 1150 276 1158
rect 294 1150 296 1158
rect 304 1150 306 1158
rect 324 1150 326 1158
rect 334 1150 336 1158
rect 354 1150 356 1158
rect 364 1150 366 1158
rect 384 1150 386 1158
rect 394 1150 396 1158
rect 414 1150 416 1158
rect 424 1150 426 1158
rect 444 1150 446 1158
rect 454 1150 456 1158
rect 474 1150 476 1158
rect 484 1150 486 1158
rect 504 1150 506 1158
rect 514 1150 516 1158
rect 534 1150 536 1158
rect 544 1150 546 1158
rect 554 1150 560 1158
rect 42 1148 76 1150
rect 84 1148 106 1150
rect 114 1148 136 1150
rect 144 1148 166 1150
rect 174 1148 196 1150
rect 204 1148 226 1150
rect 234 1148 256 1150
rect 264 1148 286 1150
rect 294 1148 316 1150
rect 324 1148 346 1150
rect 354 1148 376 1150
rect 384 1148 406 1150
rect 414 1148 436 1150
rect 444 1148 466 1150
rect 474 1148 496 1150
rect 504 1148 526 1150
rect 534 1148 560 1150
rect 42 1140 46 1148
rect 54 1140 56 1148
rect 64 1140 66 1148
rect 74 1140 76 1148
rect 94 1140 96 1148
rect 104 1140 106 1148
rect 124 1140 126 1148
rect 134 1140 136 1148
rect 154 1140 156 1148
rect 164 1140 166 1148
rect 184 1140 186 1148
rect 194 1140 196 1148
rect 214 1140 216 1148
rect 224 1140 226 1148
rect 244 1140 246 1148
rect 254 1140 256 1148
rect 274 1140 276 1148
rect 284 1140 286 1148
rect 304 1140 306 1148
rect 314 1140 316 1148
rect 334 1140 336 1148
rect 344 1140 346 1148
rect 364 1140 366 1148
rect 374 1140 376 1148
rect 394 1140 396 1148
rect 404 1140 406 1148
rect 424 1140 426 1148
rect 434 1140 436 1148
rect 454 1140 456 1148
rect 464 1140 466 1148
rect 484 1140 486 1148
rect 494 1140 496 1148
rect 514 1140 516 1148
rect 524 1140 526 1148
rect 544 1140 546 1148
rect 554 1140 560 1148
rect 42 1138 76 1140
rect 84 1138 106 1140
rect 114 1138 136 1140
rect 144 1138 166 1140
rect 174 1138 196 1140
rect 204 1138 226 1140
rect 234 1138 256 1140
rect 264 1138 286 1140
rect 294 1138 316 1140
rect 324 1138 346 1140
rect 354 1138 376 1140
rect 384 1138 406 1140
rect 414 1138 436 1140
rect 444 1138 466 1140
rect 474 1138 496 1140
rect 504 1138 526 1140
rect 534 1138 560 1140
rect 42 1130 46 1138
rect 54 1130 56 1138
rect 64 1130 66 1138
rect 84 1130 86 1138
rect 94 1130 96 1138
rect 114 1130 116 1138
rect 124 1130 126 1138
rect 144 1130 146 1138
rect 154 1130 156 1138
rect 174 1130 176 1138
rect 184 1130 186 1138
rect 204 1130 206 1138
rect 214 1130 216 1138
rect 234 1130 236 1138
rect 244 1130 246 1138
rect 264 1130 266 1138
rect 274 1130 276 1138
rect 294 1130 296 1138
rect 304 1130 306 1138
rect 324 1130 326 1138
rect 334 1130 336 1138
rect 354 1130 356 1138
rect 364 1130 366 1138
rect 384 1130 386 1138
rect 394 1130 396 1138
rect 414 1130 416 1138
rect 424 1130 426 1138
rect 444 1130 446 1138
rect 454 1130 456 1138
rect 474 1130 476 1138
rect 484 1130 486 1138
rect 504 1130 506 1138
rect 514 1130 516 1138
rect 534 1130 536 1138
rect 544 1130 546 1138
rect 554 1130 560 1138
rect 42 1128 76 1130
rect 84 1128 106 1130
rect 114 1128 136 1130
rect 144 1128 166 1130
rect 174 1128 196 1130
rect 204 1128 226 1130
rect 234 1128 256 1130
rect 264 1128 286 1130
rect 294 1128 316 1130
rect 324 1128 346 1130
rect 354 1128 376 1130
rect 384 1128 406 1130
rect 414 1128 436 1130
rect 444 1128 466 1130
rect 474 1128 496 1130
rect 504 1128 526 1130
rect 534 1128 560 1130
rect 42 1120 46 1128
rect 54 1120 56 1128
rect 64 1120 66 1128
rect 74 1120 76 1128
rect 94 1120 96 1128
rect 104 1120 106 1128
rect 124 1120 126 1128
rect 134 1120 136 1128
rect 154 1120 156 1128
rect 164 1120 166 1128
rect 184 1120 186 1128
rect 194 1120 196 1128
rect 214 1120 216 1128
rect 224 1120 226 1128
rect 244 1120 246 1128
rect 254 1120 256 1128
rect 274 1120 276 1128
rect 284 1120 286 1128
rect 304 1120 306 1128
rect 314 1120 316 1128
rect 334 1120 336 1128
rect 344 1120 346 1128
rect 364 1120 366 1128
rect 374 1120 376 1128
rect 394 1120 396 1128
rect 404 1120 406 1128
rect 424 1120 426 1128
rect 434 1120 436 1128
rect 454 1120 456 1128
rect 464 1120 466 1128
rect 484 1120 486 1128
rect 494 1120 496 1128
rect 42 1118 86 1120
rect 42 1110 46 1118
rect 54 1110 56 1118
rect 64 1110 66 1118
rect 74 1110 76 1118
rect 84 1110 86 1118
rect 42 1108 86 1110
rect 94 1110 100 1120
rect 204 1110 396 1120
rect 500 1110 506 1120
rect 94 1108 506 1110
rect 42 1100 46 1108
rect 54 1100 56 1108
rect 64 1100 66 1108
rect 74 1100 76 1108
rect 94 1100 96 1108
rect 104 1100 106 1108
rect 124 1100 126 1108
rect 134 1100 136 1108
rect 154 1100 156 1108
rect 164 1100 166 1108
rect 184 1100 186 1108
rect 194 1100 196 1108
rect 214 1100 216 1108
rect 224 1100 226 1108
rect 244 1100 246 1108
rect 254 1100 256 1108
rect 274 1100 276 1108
rect 284 1100 286 1108
rect 304 1100 306 1108
rect 314 1100 316 1108
rect 334 1100 336 1108
rect 344 1100 346 1108
rect 364 1100 366 1108
rect 374 1100 376 1108
rect 394 1100 396 1108
rect 404 1100 406 1108
rect 424 1100 426 1108
rect 434 1100 436 1108
rect 454 1100 456 1108
rect 464 1100 466 1108
rect 484 1100 486 1108
rect 494 1100 496 1108
rect 514 1100 516 1128
rect 524 1100 526 1128
rect 544 1120 546 1128
rect 554 1120 560 1128
rect 534 1118 560 1120
rect 534 1110 536 1118
rect 544 1110 546 1118
rect 554 1110 560 1118
rect 534 1108 560 1110
rect 544 1100 546 1108
rect 554 1100 560 1108
rect 42 1098 76 1100
rect 84 1098 106 1100
rect 114 1098 136 1100
rect 144 1098 166 1100
rect 174 1098 196 1100
rect 204 1098 226 1100
rect 234 1098 256 1100
rect 264 1098 286 1100
rect 294 1098 316 1100
rect 324 1098 346 1100
rect 354 1098 376 1100
rect 384 1098 406 1100
rect 414 1098 436 1100
rect 444 1098 466 1100
rect 474 1098 496 1100
rect 504 1098 526 1100
rect 534 1098 560 1100
rect 42 1090 46 1098
rect 54 1090 56 1098
rect 64 1090 66 1098
rect 84 1090 86 1098
rect 94 1090 96 1098
rect 114 1090 116 1098
rect 124 1090 126 1098
rect 144 1090 146 1098
rect 154 1090 156 1098
rect 174 1090 176 1098
rect 184 1090 186 1098
rect 204 1090 206 1098
rect 214 1090 216 1098
rect 234 1090 236 1098
rect 244 1090 246 1098
rect 264 1090 266 1098
rect 274 1090 276 1098
rect 294 1090 296 1098
rect 304 1090 306 1098
rect 324 1090 326 1098
rect 334 1090 336 1098
rect 354 1090 356 1098
rect 364 1090 366 1098
rect 384 1090 386 1098
rect 394 1090 396 1098
rect 414 1090 416 1098
rect 424 1090 426 1098
rect 444 1090 446 1098
rect 454 1090 456 1098
rect 474 1090 476 1098
rect 484 1090 486 1098
rect 504 1090 506 1098
rect 514 1090 516 1098
rect 534 1090 536 1098
rect 544 1090 546 1098
rect 554 1090 560 1098
rect 42 1088 76 1090
rect 84 1088 106 1090
rect 114 1088 136 1090
rect 144 1088 166 1090
rect 174 1088 196 1090
rect 204 1088 226 1090
rect 234 1088 256 1090
rect 264 1088 286 1090
rect 294 1088 316 1090
rect 324 1088 346 1090
rect 354 1088 376 1090
rect 384 1088 406 1090
rect 414 1088 436 1090
rect 444 1088 466 1090
rect 474 1088 496 1090
rect 504 1088 526 1090
rect 534 1088 560 1090
rect 42 1080 46 1088
rect 54 1080 56 1088
rect 64 1080 66 1088
rect 74 1080 76 1088
rect 94 1080 96 1088
rect 104 1080 106 1088
rect 124 1080 126 1088
rect 134 1080 136 1088
rect 154 1080 156 1088
rect 164 1080 166 1088
rect 184 1080 186 1088
rect 194 1080 196 1088
rect 214 1080 216 1088
rect 224 1080 226 1088
rect 244 1080 246 1088
rect 254 1080 256 1088
rect 274 1080 276 1088
rect 284 1080 286 1088
rect 304 1080 306 1088
rect 314 1080 316 1088
rect 334 1080 336 1088
rect 344 1080 346 1088
rect 364 1080 366 1088
rect 374 1080 376 1088
rect 394 1080 396 1088
rect 404 1080 406 1088
rect 424 1080 426 1088
rect 434 1080 436 1088
rect 454 1080 456 1088
rect 464 1080 466 1088
rect 484 1080 486 1088
rect 494 1080 496 1088
rect 514 1080 516 1088
rect 524 1080 526 1088
rect 544 1080 546 1088
rect 554 1080 560 1088
rect 42 1078 76 1080
rect 84 1078 106 1080
rect 114 1078 136 1080
rect 144 1078 166 1080
rect 174 1078 196 1080
rect 204 1078 226 1080
rect 234 1078 256 1080
rect 264 1078 286 1080
rect 294 1078 316 1080
rect 324 1078 346 1080
rect 354 1078 376 1080
rect 384 1078 406 1080
rect 414 1078 436 1080
rect 444 1078 466 1080
rect 474 1078 496 1080
rect 504 1078 526 1080
rect 534 1078 560 1080
rect 42 1070 46 1078
rect 54 1070 56 1078
rect 64 1070 66 1078
rect 84 1070 86 1078
rect 94 1070 96 1078
rect 114 1070 116 1078
rect 124 1070 126 1078
rect 144 1070 146 1078
rect 154 1070 156 1078
rect 174 1070 176 1078
rect 184 1070 186 1078
rect 204 1070 206 1078
rect 214 1070 216 1078
rect 234 1070 236 1078
rect 244 1070 246 1078
rect 264 1070 266 1078
rect 274 1070 276 1078
rect 294 1070 296 1078
rect 304 1070 306 1078
rect 324 1070 326 1078
rect 334 1070 336 1078
rect 354 1070 356 1078
rect 364 1070 366 1078
rect 384 1070 386 1078
rect 394 1070 396 1078
rect 414 1070 416 1078
rect 424 1070 426 1078
rect 444 1070 446 1078
rect 454 1070 456 1078
rect 474 1070 476 1078
rect 484 1070 486 1078
rect 504 1070 506 1078
rect 514 1070 516 1078
rect 534 1070 536 1078
rect 544 1070 546 1078
rect 554 1070 560 1078
rect 42 1068 76 1070
rect 84 1068 106 1070
rect 114 1068 136 1070
rect 144 1068 166 1070
rect 174 1068 196 1070
rect 204 1068 226 1070
rect 234 1068 256 1070
rect 264 1068 286 1070
rect 294 1068 316 1070
rect 324 1068 346 1070
rect 354 1068 376 1070
rect 384 1068 406 1070
rect 414 1068 436 1070
rect 444 1068 466 1070
rect 474 1068 496 1070
rect 504 1068 526 1070
rect 534 1068 560 1070
rect 42 1060 46 1068
rect 54 1060 56 1068
rect 64 1060 66 1068
rect 74 1060 76 1068
rect 94 1060 96 1068
rect 104 1060 106 1068
rect 124 1060 126 1068
rect 134 1060 136 1068
rect 154 1060 156 1068
rect 164 1060 166 1068
rect 184 1060 186 1068
rect 194 1060 196 1068
rect 214 1060 216 1068
rect 224 1060 226 1068
rect 244 1060 246 1068
rect 254 1060 256 1068
rect 274 1060 276 1068
rect 284 1060 286 1068
rect 304 1060 306 1068
rect 314 1060 316 1068
rect 334 1060 336 1068
rect 344 1060 346 1068
rect 364 1060 366 1068
rect 374 1060 376 1068
rect 394 1060 396 1068
rect 404 1060 406 1068
rect 424 1060 426 1068
rect 434 1060 436 1068
rect 454 1060 456 1068
rect 464 1060 466 1068
rect 484 1060 486 1068
rect 494 1060 496 1068
rect 514 1060 516 1068
rect 524 1060 526 1068
rect 544 1060 546 1068
rect 554 1060 560 1068
rect 42 1058 76 1060
rect 84 1058 106 1060
rect 114 1058 136 1060
rect 144 1058 166 1060
rect 174 1058 196 1060
rect 204 1058 226 1060
rect 234 1058 256 1060
rect 264 1058 286 1060
rect 294 1058 316 1060
rect 324 1058 346 1060
rect 354 1058 376 1060
rect 384 1058 406 1060
rect 414 1058 436 1060
rect 444 1058 466 1060
rect 474 1058 496 1060
rect 504 1058 526 1060
rect 534 1058 560 1060
rect 42 1050 46 1058
rect 54 1050 56 1058
rect 64 1050 66 1058
rect 84 1050 86 1058
rect 94 1050 96 1058
rect 114 1050 116 1058
rect 124 1050 126 1058
rect 144 1050 146 1058
rect 154 1050 156 1058
rect 174 1050 176 1058
rect 184 1050 186 1058
rect 204 1050 206 1058
rect 214 1050 216 1058
rect 234 1050 236 1058
rect 244 1050 246 1058
rect 264 1050 266 1058
rect 274 1050 276 1058
rect 294 1050 296 1058
rect 304 1050 306 1058
rect 324 1050 326 1058
rect 334 1050 336 1058
rect 354 1050 356 1058
rect 364 1050 366 1058
rect 384 1050 386 1058
rect 394 1050 396 1058
rect 414 1050 416 1058
rect 424 1050 426 1058
rect 444 1050 446 1058
rect 454 1050 456 1058
rect 474 1050 476 1058
rect 484 1050 486 1058
rect 504 1050 506 1058
rect 514 1050 516 1058
rect 534 1050 536 1058
rect 544 1050 546 1058
rect 554 1050 560 1058
rect 42 1048 76 1050
rect 84 1048 106 1050
rect 114 1048 136 1050
rect 144 1048 166 1050
rect 174 1048 196 1050
rect 204 1048 226 1050
rect 234 1048 256 1050
rect 264 1048 286 1050
rect 294 1048 316 1050
rect 324 1048 346 1050
rect 354 1048 376 1050
rect 384 1048 406 1050
rect 414 1048 436 1050
rect 444 1048 466 1050
rect 474 1048 496 1050
rect 504 1048 526 1050
rect 534 1048 560 1050
rect 42 1040 46 1048
rect 54 1040 56 1048
rect 64 1040 66 1048
rect 74 1040 76 1048
rect 94 1040 96 1048
rect 104 1040 106 1048
rect 124 1040 126 1048
rect 134 1040 136 1048
rect 154 1040 156 1048
rect 164 1040 166 1048
rect 184 1040 186 1048
rect 194 1040 196 1048
rect 214 1040 216 1048
rect 224 1040 226 1048
rect 244 1040 246 1048
rect 254 1040 256 1048
rect 274 1040 276 1048
rect 284 1040 286 1048
rect 304 1040 306 1048
rect 314 1040 316 1048
rect 334 1040 336 1048
rect 344 1040 346 1048
rect 364 1040 366 1048
rect 374 1040 376 1048
rect 394 1040 396 1048
rect 404 1040 406 1048
rect 424 1040 426 1048
rect 434 1040 436 1048
rect 454 1040 456 1048
rect 464 1040 466 1048
rect 484 1040 486 1048
rect 494 1040 496 1048
rect 42 1038 76 1040
rect 84 1038 506 1040
rect 42 1030 46 1038
rect 54 1030 56 1038
rect 64 1030 66 1038
rect 84 1030 86 1038
rect 94 1030 506 1038
rect 42 1028 76 1030
rect 84 1028 506 1030
rect 42 1020 46 1028
rect 54 1020 56 1028
rect 64 1020 66 1028
rect 74 1020 76 1028
rect 94 1020 96 1028
rect 104 1020 106 1028
rect 124 1020 126 1028
rect 134 1020 136 1028
rect 154 1020 156 1028
rect 164 1020 166 1028
rect 184 1020 186 1028
rect 194 1020 196 1028
rect 214 1020 216 1028
rect 224 1020 226 1028
rect 244 1020 246 1028
rect 254 1020 256 1028
rect 274 1020 276 1028
rect 284 1020 286 1028
rect 304 1020 306 1028
rect 314 1020 316 1028
rect 334 1020 336 1028
rect 344 1020 346 1028
rect 364 1020 366 1028
rect 374 1020 376 1028
rect 394 1020 396 1028
rect 404 1020 406 1028
rect 424 1020 426 1028
rect 434 1020 436 1028
rect 454 1020 456 1028
rect 464 1020 466 1028
rect 484 1020 486 1028
rect 494 1020 496 1028
rect 514 1020 516 1048
rect 524 1020 526 1048
rect 544 1040 546 1048
rect 554 1040 560 1048
rect 534 1038 560 1040
rect 534 1030 536 1038
rect 544 1030 546 1038
rect 554 1030 560 1038
rect 534 1028 560 1030
rect 544 1020 546 1028
rect 554 1020 560 1028
rect 42 1018 76 1020
rect 84 1018 106 1020
rect 114 1018 136 1020
rect 144 1018 166 1020
rect 174 1018 196 1020
rect 204 1018 226 1020
rect 234 1018 256 1020
rect 264 1018 286 1020
rect 294 1018 316 1020
rect 324 1018 346 1020
rect 354 1018 376 1020
rect 384 1018 406 1020
rect 414 1018 436 1020
rect 444 1018 466 1020
rect 474 1018 496 1020
rect 504 1018 526 1020
rect 534 1018 560 1020
rect 42 1010 46 1018
rect 54 1010 56 1018
rect 64 1010 66 1018
rect 84 1010 86 1018
rect 94 1010 96 1018
rect 114 1010 116 1018
rect 124 1010 126 1018
rect 144 1010 146 1018
rect 154 1010 156 1018
rect 174 1010 176 1018
rect 184 1010 186 1018
rect 204 1010 206 1018
rect 214 1010 216 1018
rect 234 1010 236 1018
rect 244 1010 246 1018
rect 264 1010 266 1018
rect 274 1010 276 1018
rect 294 1010 296 1018
rect 304 1010 306 1018
rect 324 1010 326 1018
rect 334 1010 336 1018
rect 354 1010 356 1018
rect 364 1010 366 1018
rect 384 1010 386 1018
rect 394 1010 396 1018
rect 414 1010 416 1018
rect 424 1010 426 1018
rect 444 1010 446 1018
rect 454 1010 456 1018
rect 474 1010 476 1018
rect 484 1010 486 1018
rect 504 1010 506 1018
rect 514 1010 516 1018
rect 534 1010 536 1018
rect 544 1010 546 1018
rect 554 1010 560 1018
rect 42 1008 76 1010
rect 84 1008 106 1010
rect 114 1008 136 1010
rect 144 1008 166 1010
rect 174 1008 196 1010
rect 204 1008 226 1010
rect 234 1008 256 1010
rect 264 1008 286 1010
rect 294 1008 316 1010
rect 324 1008 346 1010
rect 354 1008 376 1010
rect 384 1008 406 1010
rect 414 1008 436 1010
rect 444 1008 466 1010
rect 474 1008 496 1010
rect 504 1008 526 1010
rect 534 1008 560 1010
rect 42 1000 46 1008
rect 54 1000 56 1008
rect 64 1000 66 1008
rect 74 1000 76 1008
rect 94 1000 96 1008
rect 104 1000 106 1008
rect 124 1000 126 1008
rect 134 1000 136 1008
rect 154 1000 156 1008
rect 164 1000 166 1008
rect 184 1000 186 1008
rect 194 1000 196 1008
rect 214 1000 216 1008
rect 224 1000 226 1008
rect 244 1000 246 1008
rect 254 1000 256 1008
rect 274 1000 276 1008
rect 284 1000 286 1008
rect 304 1000 306 1008
rect 314 1000 316 1008
rect 334 1000 336 1008
rect 344 1000 346 1008
rect 364 1000 366 1008
rect 374 1000 376 1008
rect 394 1000 396 1008
rect 404 1000 406 1008
rect 424 1000 426 1008
rect 434 1000 436 1008
rect 454 1000 456 1008
rect 464 1000 466 1008
rect 484 1000 486 1008
rect 494 1000 496 1008
rect 514 1000 516 1008
rect 524 1000 526 1008
rect 544 1000 546 1008
rect 554 1000 560 1008
rect 42 998 76 1000
rect 84 998 106 1000
rect 114 998 136 1000
rect 144 998 166 1000
rect 174 998 196 1000
rect 204 998 226 1000
rect 234 998 256 1000
rect 264 998 286 1000
rect 294 998 316 1000
rect 324 998 346 1000
rect 354 998 376 1000
rect 384 998 406 1000
rect 414 998 436 1000
rect 444 998 466 1000
rect 474 998 496 1000
rect 504 998 526 1000
rect 534 998 560 1000
rect 42 990 46 998
rect 54 990 56 998
rect 64 990 66 998
rect 84 990 86 998
rect 94 990 96 998
rect 114 990 116 998
rect 124 990 126 998
rect 144 990 146 998
rect 154 990 156 998
rect 174 990 176 998
rect 184 990 186 998
rect 204 990 206 998
rect 214 990 216 998
rect 234 990 236 998
rect 244 990 246 998
rect 264 990 266 998
rect 274 990 276 998
rect 294 990 296 998
rect 304 990 306 998
rect 324 990 326 998
rect 334 990 336 998
rect 354 990 356 998
rect 364 990 366 998
rect 384 990 386 998
rect 394 990 396 998
rect 414 990 416 998
rect 424 990 426 998
rect 444 990 446 998
rect 454 990 456 998
rect 474 990 476 998
rect 484 990 486 998
rect 504 990 506 998
rect 514 990 516 998
rect 534 990 536 998
rect 544 990 546 998
rect 554 990 560 998
rect 42 988 76 990
rect 84 988 106 990
rect 114 988 136 990
rect 144 988 166 990
rect 174 988 196 990
rect 204 988 226 990
rect 234 988 256 990
rect 264 988 286 990
rect 294 988 316 990
rect 324 988 346 990
rect 354 988 376 990
rect 384 988 406 990
rect 414 988 436 990
rect 444 988 466 990
rect 474 988 496 990
rect 504 988 526 990
rect 534 988 560 990
rect 42 980 46 988
rect 54 980 56 988
rect 64 980 66 988
rect 74 980 76 988
rect 94 980 96 988
rect 104 980 106 988
rect 124 980 126 988
rect 134 980 136 988
rect 154 980 156 988
rect 164 980 166 988
rect 184 980 186 988
rect 194 980 196 988
rect 214 980 216 988
rect 224 980 226 988
rect 244 980 246 988
rect 254 980 256 988
rect 274 980 276 988
rect 284 980 286 988
rect 304 980 306 988
rect 314 980 316 988
rect 334 980 336 988
rect 344 980 346 988
rect 364 980 366 988
rect 374 980 376 988
rect 394 980 396 988
rect 404 980 406 988
rect 424 980 426 988
rect 434 980 436 988
rect 454 980 456 988
rect 464 980 466 988
rect 484 980 486 988
rect 494 980 496 988
rect 514 980 516 988
rect 524 980 526 988
rect 544 980 546 988
rect 554 980 560 988
rect 42 978 76 980
rect 84 978 106 980
rect 114 978 136 980
rect 144 978 166 980
rect 174 978 196 980
rect 204 978 226 980
rect 234 978 256 980
rect 264 978 286 980
rect 294 978 316 980
rect 324 978 346 980
rect 354 978 376 980
rect 384 978 406 980
rect 414 978 436 980
rect 444 978 466 980
rect 474 978 496 980
rect 504 978 526 980
rect 534 978 560 980
rect 42 970 46 978
rect 54 970 56 978
rect 64 970 66 978
rect 84 970 86 978
rect 94 970 96 978
rect 114 970 116 978
rect 124 970 126 978
rect 144 970 146 978
rect 154 970 156 978
rect 174 970 176 978
rect 184 970 186 978
rect 204 970 206 978
rect 214 970 216 978
rect 234 970 236 978
rect 244 970 246 978
rect 264 970 266 978
rect 274 970 276 978
rect 294 970 296 978
rect 304 970 306 978
rect 324 970 326 978
rect 334 970 336 978
rect 354 970 356 978
rect 364 970 366 978
rect 384 970 386 978
rect 394 970 396 978
rect 414 970 416 978
rect 424 970 426 978
rect 444 970 446 978
rect 454 970 456 978
rect 474 970 476 978
rect 484 970 486 978
rect 504 970 506 978
rect 514 970 516 978
rect 534 970 536 978
rect 544 970 546 978
rect 554 970 560 978
rect 42 968 100 970
rect 42 960 46 968
rect 54 960 100 968
rect 204 960 396 970
rect 500 968 560 970
rect 500 960 536 968
rect 544 960 546 968
rect 554 960 560 968
rect 42 958 560 960
rect 42 950 46 958
rect 54 950 56 958
rect 64 950 66 958
rect 84 950 86 958
rect 94 950 96 958
rect 114 950 116 958
rect 124 950 126 958
rect 144 950 146 958
rect 154 950 156 958
rect 174 950 176 958
rect 184 950 186 958
rect 204 950 206 958
rect 214 950 216 958
rect 234 950 236 958
rect 244 950 246 958
rect 264 950 266 958
rect 274 950 276 958
rect 294 950 296 958
rect 304 950 306 958
rect 324 950 326 958
rect 334 950 336 958
rect 354 950 356 958
rect 364 950 366 958
rect 384 950 386 958
rect 394 950 396 958
rect 414 950 416 958
rect 424 950 426 958
rect 444 950 446 958
rect 454 950 456 958
rect 474 950 476 958
rect 484 950 486 958
rect 504 950 506 958
rect 514 950 516 958
rect 534 950 536 958
rect 544 950 546 958
rect 554 950 560 958
rect 42 948 76 950
rect 84 948 106 950
rect 114 948 136 950
rect 144 948 166 950
rect 174 948 196 950
rect 204 948 226 950
rect 234 948 256 950
rect 264 948 286 950
rect 294 948 316 950
rect 324 948 346 950
rect 354 948 376 950
rect 384 948 406 950
rect 414 948 436 950
rect 444 948 466 950
rect 474 948 496 950
rect 504 948 526 950
rect 534 948 560 950
rect 42 940 46 948
rect 54 940 56 948
rect 64 940 66 948
rect 74 940 76 948
rect 94 940 96 948
rect 104 940 106 948
rect 124 940 126 948
rect 134 940 136 948
rect 154 940 156 948
rect 164 940 166 948
rect 184 940 186 948
rect 194 940 196 948
rect 214 940 216 948
rect 224 940 226 948
rect 244 940 246 948
rect 254 940 256 948
rect 274 940 276 948
rect 284 940 286 948
rect 304 940 306 948
rect 314 940 316 948
rect 334 940 336 948
rect 344 940 346 948
rect 364 940 366 948
rect 374 940 376 948
rect 394 940 396 948
rect 404 940 406 948
rect 424 940 426 948
rect 434 940 436 948
rect 454 940 456 948
rect 464 940 466 948
rect 484 940 486 948
rect 494 940 496 948
rect 514 940 516 948
rect 524 940 526 948
rect 544 940 546 948
rect 554 940 560 948
rect 42 938 76 940
rect 84 938 106 940
rect 114 938 136 940
rect 144 938 166 940
rect 174 938 196 940
rect 204 938 226 940
rect 234 938 256 940
rect 264 938 286 940
rect 294 938 316 940
rect 324 938 346 940
rect 354 938 376 940
rect 384 938 406 940
rect 414 938 436 940
rect 444 938 466 940
rect 474 938 496 940
rect 504 938 526 940
rect 534 938 560 940
rect 42 930 46 938
rect 54 930 56 938
rect 64 930 66 938
rect 84 930 86 938
rect 94 930 96 938
rect 114 930 116 938
rect 124 930 126 938
rect 144 930 146 938
rect 154 930 156 938
rect 174 930 176 938
rect 184 930 186 938
rect 204 930 206 938
rect 214 930 216 938
rect 234 930 236 938
rect 244 930 246 938
rect 264 930 266 938
rect 274 930 276 938
rect 294 930 296 938
rect 304 930 306 938
rect 324 930 326 938
rect 334 930 336 938
rect 354 930 356 938
rect 364 930 366 938
rect 384 930 386 938
rect 394 930 396 938
rect 414 930 416 938
rect 424 930 426 938
rect 444 930 446 938
rect 454 930 456 938
rect 474 930 476 938
rect 484 930 486 938
rect 504 930 506 938
rect 514 930 516 938
rect 534 930 536 938
rect 544 930 546 938
rect 554 930 560 938
rect 42 928 76 930
rect 84 928 106 930
rect 114 928 136 930
rect 144 928 166 930
rect 174 928 196 930
rect 204 928 226 930
rect 234 928 256 930
rect 264 928 286 930
rect 294 928 316 930
rect 324 928 346 930
rect 354 928 376 930
rect 384 928 406 930
rect 414 928 436 930
rect 444 928 466 930
rect 474 928 496 930
rect 504 928 526 930
rect 534 928 560 930
rect 42 920 46 928
rect 54 920 56 928
rect 64 920 66 928
rect 74 920 76 928
rect 94 920 96 928
rect 104 920 106 928
rect 124 920 126 928
rect 134 920 136 928
rect 154 920 156 928
rect 164 920 166 928
rect 184 920 186 928
rect 194 920 196 928
rect 214 920 216 928
rect 224 920 226 928
rect 244 920 246 928
rect 254 920 256 928
rect 274 920 276 928
rect 284 920 286 928
rect 304 920 306 928
rect 314 920 316 928
rect 334 920 336 928
rect 344 920 346 928
rect 364 920 366 928
rect 374 920 376 928
rect 394 920 396 928
rect 404 920 406 928
rect 424 920 426 928
rect 434 920 436 928
rect 454 920 456 928
rect 464 920 466 928
rect 484 920 486 928
rect 494 920 496 928
rect 514 920 516 928
rect 524 920 526 928
rect 544 920 546 928
rect 554 920 560 928
rect 42 918 76 920
rect 84 918 106 920
rect 114 918 136 920
rect 144 918 166 920
rect 174 918 196 920
rect 204 918 226 920
rect 234 918 256 920
rect 264 918 286 920
rect 294 918 316 920
rect 324 918 346 920
rect 354 918 376 920
rect 384 918 406 920
rect 414 918 436 920
rect 444 918 466 920
rect 474 918 496 920
rect 504 918 526 920
rect 534 918 560 920
rect 42 910 46 918
rect 54 910 56 918
rect 64 910 66 918
rect 84 910 86 918
rect 94 910 96 918
rect 114 910 116 918
rect 124 910 126 918
rect 144 910 146 918
rect 154 910 156 918
rect 174 910 176 918
rect 184 910 186 918
rect 204 910 206 918
rect 214 910 216 918
rect 234 910 236 918
rect 244 910 246 918
rect 264 910 266 918
rect 274 910 276 918
rect 294 910 296 918
rect 304 910 306 918
rect 324 910 326 918
rect 334 910 336 918
rect 354 910 356 918
rect 364 910 366 918
rect 384 910 386 918
rect 394 910 396 918
rect 414 910 416 918
rect 424 910 426 918
rect 444 910 446 918
rect 454 910 456 918
rect 474 910 476 918
rect 484 910 486 918
rect 504 910 506 918
rect 514 910 516 918
rect 534 910 536 918
rect 544 910 546 918
rect 554 910 560 918
rect 42 908 76 910
rect 84 908 106 910
rect 114 908 136 910
rect 144 908 166 910
rect 174 908 196 910
rect 204 908 226 910
rect 234 908 256 910
rect 264 908 286 910
rect 294 908 316 910
rect 324 908 346 910
rect 354 908 376 910
rect 384 908 406 910
rect 414 908 436 910
rect 444 908 466 910
rect 474 908 496 910
rect 504 908 526 910
rect 534 908 560 910
rect 42 900 46 908
rect 54 900 56 908
rect 64 900 66 908
rect 74 900 76 908
rect 94 900 96 908
rect 104 900 106 908
rect 124 900 126 908
rect 134 900 136 908
rect 154 900 156 908
rect 164 900 166 908
rect 184 900 186 908
rect 194 900 196 908
rect 214 900 216 908
rect 224 900 226 908
rect 244 900 246 908
rect 254 900 256 908
rect 274 900 276 908
rect 284 900 286 908
rect 304 900 306 908
rect 314 900 316 908
rect 334 900 336 908
rect 344 900 346 908
rect 364 900 366 908
rect 374 900 376 908
rect 394 900 396 908
rect 404 900 406 908
rect 424 900 426 908
rect 434 900 436 908
rect 454 900 456 908
rect 464 900 466 908
rect 484 900 486 908
rect 494 900 496 908
rect 514 900 516 908
rect 524 900 526 908
rect 544 900 546 908
rect 554 900 560 908
rect 42 898 76 900
rect 84 898 106 900
rect 114 898 136 900
rect 144 898 166 900
rect 174 898 196 900
rect 204 898 226 900
rect 234 898 256 900
rect 264 898 286 900
rect 294 898 316 900
rect 324 898 346 900
rect 354 898 376 900
rect 384 898 406 900
rect 414 898 436 900
rect 444 898 466 900
rect 474 898 496 900
rect 504 898 526 900
rect 534 898 560 900
rect 42 890 46 898
rect 54 890 56 898
rect 64 890 66 898
rect 84 890 86 898
rect 94 890 96 898
rect 114 890 116 898
rect 124 890 126 898
rect 144 890 146 898
rect 154 890 156 898
rect 174 890 176 898
rect 184 890 186 898
rect 204 890 206 898
rect 214 890 216 898
rect 234 890 236 898
rect 244 890 246 898
rect 264 890 266 898
rect 274 890 276 898
rect 294 890 296 898
rect 304 890 306 898
rect 324 890 326 898
rect 334 890 336 898
rect 354 890 356 898
rect 364 890 366 898
rect 384 890 386 898
rect 394 890 396 898
rect 414 890 416 898
rect 424 890 426 898
rect 444 890 446 898
rect 454 890 456 898
rect 474 890 476 898
rect 484 890 486 898
rect 504 890 506 898
rect 514 890 516 898
rect 534 890 536 898
rect 544 890 546 898
rect 554 890 560 898
rect 42 888 76 890
rect 84 888 106 890
rect 114 888 136 890
rect 144 888 166 890
rect 174 888 196 890
rect 204 888 226 890
rect 234 888 256 890
rect 264 888 286 890
rect 294 888 316 890
rect 324 888 346 890
rect 354 888 376 890
rect 384 888 406 890
rect 414 888 436 890
rect 444 888 466 890
rect 474 888 496 890
rect 504 888 526 890
rect 534 888 560 890
rect 42 880 46 888
rect 54 880 56 888
rect 42 878 56 880
rect 64 880 66 888
rect 74 880 76 888
rect 64 878 76 880
rect 94 880 96 888
rect 104 880 106 888
rect 94 878 106 880
rect 124 880 126 888
rect 134 880 136 888
rect 124 878 136 880
rect 154 880 156 888
rect 164 880 166 888
rect 154 878 166 880
rect 184 880 186 888
rect 194 880 196 888
rect 184 878 196 880
rect 214 880 216 888
rect 224 880 226 888
rect 214 878 226 880
rect 244 880 246 888
rect 254 880 256 888
rect 244 878 256 880
rect 274 880 276 888
rect 284 880 286 888
rect 274 878 286 880
rect 304 880 306 888
rect 314 880 316 888
rect 304 878 316 880
rect 334 880 336 888
rect 344 880 346 888
rect 334 878 346 880
rect 364 880 366 888
rect 374 880 376 888
rect 364 878 376 880
rect 394 880 396 888
rect 404 880 406 888
rect 394 878 406 880
rect 424 880 426 888
rect 434 880 436 888
rect 424 878 436 880
rect 454 880 456 888
rect 464 880 466 888
rect 454 878 466 880
rect 484 880 486 888
rect 494 880 496 888
rect 484 878 496 880
rect 514 880 516 888
rect 524 880 526 888
rect 514 878 526 880
rect 544 880 546 888
rect 554 880 560 888
rect 544 878 560 880
rect 42 870 46 878
rect 554 870 560 878
rect 42 866 560 870
rect 0 838 21 840
rect 204 848 396 866
rect 0 836 198 838
rect 0 828 4 836
rect 12 828 14 836
rect 22 828 24 836
rect 42 828 44 836
rect 52 828 54 836
rect 72 828 74 836
rect 82 828 84 836
rect 102 828 104 836
rect 112 828 114 836
rect 132 828 134 836
rect 142 828 144 836
rect 162 828 164 836
rect 172 828 174 836
rect 182 828 184 836
rect 192 828 198 836
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 198 828
rect 0 818 4 826
rect 12 818 14 826
rect 22 818 24 826
rect 32 818 34 826
rect 52 818 54 826
rect 62 818 64 826
rect 82 818 84 826
rect 92 818 94 826
rect 112 818 114 826
rect 122 818 124 826
rect 142 818 144 826
rect 152 818 154 826
rect 172 818 174 826
rect 182 818 184 826
rect 192 818 198 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 198 818
rect 0 808 4 816
rect 12 808 14 816
rect 22 808 24 816
rect 42 808 44 816
rect 52 808 54 816
rect 72 808 74 816
rect 82 808 84 816
rect 102 808 104 816
rect 112 808 114 816
rect 132 808 134 816
rect 142 808 144 816
rect 162 808 164 816
rect 172 808 174 816
rect 182 808 184 816
rect 192 808 198 816
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 198 808
rect 0 798 4 806
rect 12 798 14 806
rect 22 798 24 806
rect 32 798 34 806
rect 52 798 54 806
rect 62 798 64 806
rect 82 798 84 806
rect 92 798 94 806
rect 112 798 114 806
rect 122 798 124 806
rect 142 798 144 806
rect 152 798 154 806
rect 172 798 174 806
rect 182 798 184 806
rect 192 798 198 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 198 798
rect 0 788 4 796
rect 12 788 14 796
rect 22 788 24 796
rect 42 788 44 796
rect 52 788 54 796
rect 72 788 74 796
rect 82 788 84 796
rect 102 788 104 796
rect 112 788 114 796
rect 132 788 134 796
rect 142 788 144 796
rect 162 788 164 796
rect 172 788 174 796
rect 182 788 184 796
rect 192 788 198 796
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 198 788
rect 0 778 4 786
rect 12 778 14 786
rect 22 778 24 786
rect 32 778 34 786
rect 52 778 54 786
rect 62 778 64 786
rect 82 778 84 786
rect 92 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 778 114 786
rect 122 778 124 786
rect 112 776 124 778
rect 142 778 144 786
rect 152 778 154 786
rect 142 776 154 778
rect 172 778 174 786
rect 182 778 184 786
rect 172 776 184 778
rect 0 768 4 776
rect 12 768 14 776
rect 22 768 24 776
rect 42 768 44 776
rect 52 768 54 776
rect 72 768 74 776
rect 82 768 84 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 4 766
rect 12 758 14 766
rect 22 758 24 766
rect 32 758 34 766
rect 52 758 54 766
rect 62 758 64 766
rect 82 758 84 766
rect 92 758 94 766
rect 112 766 124 768
rect 112 758 114 766
rect 122 758 124 766
rect 142 766 154 768
rect 142 758 144 766
rect 152 758 154 766
rect 172 766 184 768
rect 172 758 174 766
rect 182 758 184 766
rect 192 758 198 786
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 198 758
rect 0 748 4 756
rect 12 748 14 756
rect 22 748 24 756
rect 42 748 44 756
rect 52 748 54 756
rect 72 748 74 756
rect 82 748 84 756
rect 102 748 104 756
rect 112 748 114 756
rect 132 748 134 756
rect 142 748 144 756
rect 162 748 164 756
rect 172 748 174 756
rect 182 748 184 756
rect 192 748 198 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 198 748
rect 0 738 4 746
rect 12 738 14 746
rect 22 738 24 746
rect 32 738 34 746
rect 52 738 54 746
rect 62 738 64 746
rect 82 738 84 746
rect 92 738 94 746
rect 112 738 114 746
rect 122 738 124 746
rect 142 738 144 746
rect 152 738 154 746
rect 172 738 174 746
rect 182 738 184 746
rect 192 738 198 746
rect 0 737 198 738
rect 0 736 42 737
rect 0 728 4 736
rect 12 728 14 736
rect 22 728 24 736
rect 32 728 42 736
rect 0 727 42 728
rect 0 726 198 727
rect 0 718 4 726
rect 12 718 14 726
rect 22 718 24 726
rect 32 718 34 726
rect 52 718 54 726
rect 62 718 64 726
rect 82 718 84 726
rect 92 718 94 726
rect 112 718 114 726
rect 122 718 124 726
rect 142 718 144 726
rect 152 718 154 726
rect 172 718 174 726
rect 182 718 184 726
rect 192 718 198 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 198 718
rect 0 708 4 716
rect 12 708 14 716
rect 22 708 24 716
rect 42 708 44 716
rect 52 708 54 716
rect 72 708 74 716
rect 82 708 84 716
rect 102 708 104 716
rect 112 708 114 716
rect 132 708 134 716
rect 142 708 144 716
rect 162 708 164 716
rect 172 708 174 716
rect 182 708 184 716
rect 192 708 198 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 198 708
rect 0 698 4 706
rect 12 698 14 706
rect 22 698 24 706
rect 32 698 34 706
rect 52 698 54 706
rect 62 698 64 706
rect 82 698 84 706
rect 92 698 94 706
rect 112 698 114 706
rect 122 698 124 706
rect 142 698 144 706
rect 152 698 154 706
rect 172 698 174 706
rect 182 698 184 706
rect 192 698 198 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 198 698
rect 0 688 4 696
rect 12 688 14 696
rect 22 688 24 696
rect 42 688 44 696
rect 52 688 54 696
rect 72 688 74 696
rect 82 688 84 696
rect 102 688 104 696
rect 112 688 114 696
rect 132 688 134 696
rect 142 688 144 696
rect 162 688 164 696
rect 172 688 174 696
rect 182 688 184 696
rect 192 688 198 696
rect 204 682 280 848
rect 286 836 314 842
rect 294 828 296 836
rect 304 828 306 836
rect 286 826 314 828
rect 294 818 296 826
rect 304 818 306 826
rect 286 816 314 818
rect 294 808 296 816
rect 304 808 306 816
rect 286 806 314 808
rect 294 798 296 806
rect 304 798 306 806
rect 286 796 314 798
rect 294 788 296 796
rect 304 788 306 796
rect 286 786 314 788
rect 294 778 296 786
rect 304 778 306 786
rect 294 776 306 778
rect 286 766 296 768
rect 294 758 296 766
rect 304 766 314 768
rect 304 758 306 766
rect 286 756 314 758
rect 294 748 296 756
rect 304 748 306 756
rect 286 746 314 748
rect 294 738 296 746
rect 304 738 306 746
rect 286 736 314 738
rect 294 728 296 736
rect 304 728 306 736
rect 286 726 314 728
rect 294 718 296 726
rect 304 718 306 726
rect 286 716 314 718
rect 294 708 296 716
rect 286 706 296 708
rect 304 708 306 716
rect 304 706 314 708
rect 286 696 314 698
rect 320 682 396 848
rect 579 840 580 1319
rect 598 840 600 1338
rect 579 838 600 840
rect 402 836 600 838
rect 402 828 408 836
rect 416 828 418 836
rect 426 828 428 836
rect 436 828 438 836
rect 456 828 458 836
rect 466 828 468 836
rect 486 828 488 836
rect 496 828 498 836
rect 516 828 518 836
rect 526 828 528 836
rect 546 828 548 836
rect 556 828 558 836
rect 576 828 578 836
rect 586 828 588 836
rect 596 828 600 836
rect 402 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 402 818 408 826
rect 416 818 418 826
rect 426 818 428 826
rect 446 818 448 826
rect 456 818 458 826
rect 476 818 478 826
rect 486 818 488 826
rect 506 818 508 826
rect 516 818 518 826
rect 536 818 538 826
rect 546 818 548 826
rect 566 818 568 826
rect 576 818 578 826
rect 586 818 588 826
rect 596 818 600 826
rect 402 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 402 808 408 816
rect 416 808 418 816
rect 426 808 428 816
rect 436 808 438 816
rect 456 808 458 816
rect 466 808 468 816
rect 486 808 488 816
rect 496 808 498 816
rect 516 808 518 816
rect 526 808 528 816
rect 546 808 548 816
rect 556 808 558 816
rect 576 808 578 816
rect 586 808 588 816
rect 596 808 600 816
rect 402 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 402 798 408 806
rect 416 798 418 806
rect 426 798 428 806
rect 446 798 448 806
rect 456 798 458 806
rect 476 798 478 806
rect 486 798 488 806
rect 506 798 508 806
rect 516 798 518 806
rect 536 798 538 806
rect 546 798 548 806
rect 566 798 568 806
rect 576 798 578 806
rect 586 798 588 806
rect 596 798 600 806
rect 402 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 402 788 408 796
rect 416 788 418 796
rect 426 788 428 796
rect 436 788 438 796
rect 456 788 458 796
rect 466 788 468 796
rect 486 788 488 796
rect 496 788 498 796
rect 516 788 518 796
rect 526 788 528 796
rect 546 788 548 796
rect 556 788 558 796
rect 576 788 578 796
rect 586 788 588 796
rect 596 788 600 796
rect 402 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 402 758 408 786
rect 416 778 418 786
rect 426 778 428 786
rect 416 776 428 778
rect 446 778 448 786
rect 456 778 458 786
rect 446 776 458 778
rect 476 778 478 786
rect 486 778 488 786
rect 476 776 488 778
rect 506 778 508 786
rect 516 778 518 786
rect 536 778 538 786
rect 546 778 548 786
rect 566 778 568 786
rect 576 778 578 786
rect 586 778 588 786
rect 596 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 516 768 518 776
rect 526 768 528 776
rect 546 768 548 776
rect 556 768 558 776
rect 576 768 578 776
rect 586 768 588 776
rect 596 768 600 776
rect 416 766 428 768
rect 416 758 418 766
rect 426 758 428 766
rect 446 766 458 768
rect 446 758 448 766
rect 456 758 458 766
rect 476 766 488 768
rect 476 758 478 766
rect 486 758 488 766
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 508 766
rect 516 758 518 766
rect 536 758 538 766
rect 546 758 548 766
rect 566 758 568 766
rect 576 758 578 766
rect 586 758 588 766
rect 596 758 600 766
rect 402 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 402 748 408 756
rect 416 748 418 756
rect 426 748 428 756
rect 436 748 438 756
rect 456 748 458 756
rect 466 748 468 756
rect 486 748 488 756
rect 496 748 498 756
rect 516 748 518 756
rect 526 748 528 756
rect 546 748 548 756
rect 556 748 558 756
rect 576 748 578 756
rect 586 748 588 756
rect 596 748 600 756
rect 402 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 402 738 408 746
rect 416 738 418 746
rect 426 738 428 746
rect 446 738 448 746
rect 456 738 458 746
rect 476 738 478 746
rect 486 738 488 746
rect 506 738 508 746
rect 516 738 518 746
rect 536 738 538 746
rect 546 738 548 746
rect 566 738 568 746
rect 576 738 578 746
rect 586 738 588 746
rect 596 738 600 746
rect 560 736 600 738
rect 560 728 568 736
rect 576 728 578 736
rect 586 728 588 736
rect 596 728 600 736
rect 402 726 600 728
rect 402 718 408 726
rect 416 718 418 726
rect 426 718 428 726
rect 446 718 448 726
rect 456 718 458 726
rect 476 718 478 726
rect 486 718 488 726
rect 506 718 508 726
rect 516 718 518 726
rect 536 718 538 726
rect 546 718 548 726
rect 566 718 568 726
rect 576 718 578 726
rect 586 718 588 726
rect 596 718 600 726
rect 402 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 402 708 408 716
rect 416 708 418 716
rect 426 708 428 716
rect 436 708 438 716
rect 456 708 458 716
rect 466 708 468 716
rect 486 708 488 716
rect 496 708 498 716
rect 516 708 518 716
rect 526 708 528 716
rect 546 708 548 716
rect 556 708 558 716
rect 576 708 578 716
rect 586 708 588 716
rect 596 708 600 716
rect 402 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 402 698 408 706
rect 416 698 418 706
rect 426 698 428 706
rect 446 698 448 706
rect 456 698 458 706
rect 476 698 478 706
rect 486 698 488 706
rect 506 698 508 706
rect 516 698 518 706
rect 536 698 538 706
rect 546 698 548 706
rect 566 698 568 706
rect 576 698 578 706
rect 586 698 588 706
rect 596 698 600 706
rect 402 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 402 688 408 696
rect 416 688 418 696
rect 426 688 428 696
rect 436 688 438 696
rect 456 688 458 696
rect 466 688 468 696
rect 486 688 488 696
rect 496 688 498 696
rect 516 688 518 696
rect 526 688 528 696
rect 546 688 548 696
rect 556 688 558 696
rect 576 688 578 696
rect 586 688 588 696
rect 596 688 600 696
rect 204 652 396 682
rect 0 644 4 652
rect 12 644 14 652
rect 22 644 24 652
rect 42 644 44 652
rect 52 644 54 652
rect 72 644 74 652
rect 82 644 84 652
rect 102 644 104 652
rect 112 644 114 652
rect 132 644 134 652
rect 142 644 144 652
rect 162 644 164 652
rect 172 644 174 652
rect 192 644 194 652
rect 202 644 204 652
rect 222 644 224 652
rect 232 644 234 652
rect 242 644 244 652
rect 252 644 256 652
rect 264 644 266 652
rect 274 644 276 652
rect 294 644 296 652
rect 304 644 306 652
rect 324 644 326 652
rect 334 644 336 652
rect 344 644 348 652
rect 356 644 358 652
rect 366 644 368 652
rect 376 644 378 652
rect 396 644 398 652
rect 406 644 408 652
rect 426 644 428 652
rect 436 644 438 652
rect 456 644 458 652
rect 466 644 468 652
rect 486 644 488 652
rect 496 644 498 652
rect 516 644 518 652
rect 526 644 528 652
rect 546 644 548 652
rect 556 644 558 652
rect 576 644 578 652
rect 586 644 588 652
rect 596 644 600 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 192 642 214 644
rect 222 642 286 644
rect 294 642 316 644
rect 324 642 378 644
rect 386 642 408 644
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 0 634 4 642
rect 12 634 14 642
rect 22 634 24 642
rect 32 634 34 642
rect 52 634 54 642
rect 62 634 64 642
rect 82 634 84 642
rect 92 634 94 642
rect 112 634 114 642
rect 122 634 124 642
rect 142 634 144 642
rect 152 634 154 642
rect 172 634 174 642
rect 182 634 184 642
rect 202 634 204 642
rect 212 634 214 642
rect 232 634 234 642
rect 242 634 244 642
rect 252 634 256 642
rect 264 634 266 642
rect 274 634 276 642
rect 284 634 286 642
rect 304 634 306 642
rect 314 634 316 642
rect 334 634 336 642
rect 344 634 348 642
rect 356 634 358 642
rect 366 634 368 642
rect 386 634 388 642
rect 396 634 398 642
rect 416 634 418 642
rect 426 634 428 642
rect 446 634 448 642
rect 456 634 458 642
rect 476 634 478 642
rect 486 634 488 642
rect 506 634 508 642
rect 516 634 518 642
rect 536 634 538 642
rect 546 634 548 642
rect 566 634 568 642
rect 576 634 578 642
rect 586 634 588 642
rect 596 634 600 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 192 632 214 634
rect 222 632 286 634
rect 294 632 316 634
rect 324 632 378 634
rect 386 632 408 634
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 0 624 4 632
rect 12 624 14 632
rect 22 624 24 632
rect 42 624 44 632
rect 52 624 54 632
rect 72 624 74 632
rect 82 624 84 632
rect 102 624 104 632
rect 112 624 114 632
rect 132 624 134 632
rect 142 624 144 632
rect 162 624 164 632
rect 172 624 174 632
rect 192 624 194 632
rect 202 624 204 632
rect 222 624 224 632
rect 232 624 234 632
rect 242 624 244 632
rect 252 624 256 632
rect 264 624 266 632
rect 274 624 276 632
rect 294 624 296 632
rect 304 624 306 632
rect 324 624 326 632
rect 334 624 336 632
rect 344 624 348 632
rect 356 624 358 632
rect 366 624 368 632
rect 376 624 378 632
rect 396 624 398 632
rect 406 624 408 632
rect 426 624 428 632
rect 436 624 438 632
rect 456 624 458 632
rect 466 624 468 632
rect 486 624 488 632
rect 496 624 498 632
rect 516 624 518 632
rect 526 624 528 632
rect 546 624 548 632
rect 556 624 558 632
rect 576 624 578 632
rect 586 624 588 632
rect 596 624 600 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 192 622 214 624
rect 222 622 286 624
rect 294 622 316 624
rect 324 622 378 624
rect 386 622 408 624
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 0 614 4 622
rect 12 614 14 622
rect 22 614 24 622
rect 32 614 34 622
rect 52 614 54 622
rect 62 614 64 622
rect 82 614 84 622
rect 92 614 94 622
rect 112 614 114 622
rect 122 614 124 622
rect 142 614 144 622
rect 152 614 154 622
rect 172 614 174 622
rect 182 614 184 622
rect 202 614 204 622
rect 212 614 214 622
rect 232 614 234 622
rect 242 614 244 622
rect 252 614 256 622
rect 264 614 266 622
rect 274 614 276 622
rect 284 614 286 622
rect 304 614 306 622
rect 314 614 316 622
rect 334 614 336 622
rect 344 614 348 622
rect 356 614 358 622
rect 366 614 368 622
rect 386 614 388 622
rect 396 614 398 622
rect 416 614 418 622
rect 426 614 428 622
rect 446 614 448 622
rect 456 614 458 622
rect 476 614 478 622
rect 486 614 488 622
rect 506 614 508 622
rect 516 614 518 622
rect 536 614 538 622
rect 546 614 548 622
rect 566 614 568 622
rect 576 614 578 622
rect 586 614 588 622
rect 596 614 600 622
rect 0 612 214 614
rect 0 604 4 612
rect 12 604 14 612
rect 22 604 24 612
rect 32 604 40 612
rect 0 602 40 604
rect 204 602 214 612
rect 222 612 286 614
rect 294 612 316 614
rect 324 612 378 614
rect 222 604 224 612
rect 232 604 234 612
rect 242 604 244 612
rect 252 604 256 612
rect 264 604 266 612
rect 274 604 276 612
rect 294 604 296 612
rect 304 604 306 612
rect 324 604 326 612
rect 334 604 336 612
rect 344 604 348 612
rect 356 604 358 612
rect 366 604 368 612
rect 376 604 378 612
rect 222 602 286 604
rect 294 602 316 604
rect 324 602 378 604
rect 386 612 600 614
rect 386 602 396 612
rect 560 604 568 612
rect 576 604 578 612
rect 586 604 588 612
rect 596 604 600 612
rect 560 602 600 604
rect 0 594 4 602
rect 12 594 14 602
rect 22 594 24 602
rect 32 594 34 602
rect 52 594 54 602
rect 62 594 64 602
rect 82 594 84 602
rect 92 594 94 602
rect 112 594 114 602
rect 122 594 124 602
rect 142 594 144 602
rect 152 594 154 602
rect 172 594 174 602
rect 182 594 184 602
rect 202 594 204 602
rect 212 594 214 602
rect 232 594 234 602
rect 242 594 244 602
rect 252 594 256 602
rect 264 594 266 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 192 592 214 594
rect 222 592 266 594
rect 274 594 276 602
rect 284 594 286 602
rect 274 592 286 594
rect 304 594 306 602
rect 314 594 316 602
rect 304 592 316 594
rect 334 594 336 602
rect 344 594 348 602
rect 356 594 358 602
rect 366 594 368 602
rect 386 594 388 602
rect 396 594 398 602
rect 416 594 418 602
rect 426 594 428 602
rect 446 594 448 602
rect 456 594 458 602
rect 476 594 478 602
rect 486 594 488 602
rect 506 594 508 602
rect 516 594 518 602
rect 536 594 538 602
rect 546 594 548 602
rect 566 594 568 602
rect 576 594 578 602
rect 586 594 588 602
rect 596 594 600 602
rect 334 592 378 594
rect 386 592 408 594
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 0 584 4 592
rect 12 584 14 592
rect 22 584 24 592
rect 42 584 44 592
rect 52 584 54 592
rect 72 584 74 592
rect 82 584 84 592
rect 102 584 104 592
rect 112 584 114 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 584
rect 132 584 134 592
rect 142 584 144 592
rect 132 582 144 584
rect 162 584 164 592
rect 172 584 174 592
rect 162 582 174 584
rect 192 584 194 592
rect 202 584 204 592
rect 192 582 204 584
rect 222 584 224 592
rect 232 584 234 592
rect 222 582 234 584
rect 242 584 244 592
rect 252 584 256 592
rect 242 582 256 584
rect 0 574 4 582
rect 12 574 14 582
rect 22 574 24 582
rect 32 574 34 582
rect 52 574 54 582
rect 62 574 64 582
rect 82 574 84 582
rect 92 574 94 582
rect 252 574 256 582
rect 344 584 348 592
rect 356 584 358 592
rect 344 582 358 584
rect 366 584 368 592
rect 376 584 378 592
rect 366 582 378 584
rect 396 584 398 592
rect 406 584 408 592
rect 396 582 408 584
rect 426 584 428 592
rect 436 584 438 592
rect 426 582 438 584
rect 456 584 458 592
rect 466 584 468 592
rect 456 582 468 584
rect 486 584 488 592
rect 496 584 498 592
rect 516 584 518 592
rect 526 584 528 592
rect 546 584 548 592
rect 556 584 558 592
rect 576 584 578 592
rect 586 584 588 592
rect 596 584 600 592
rect 486 582 498 584
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 344 574 348 582
rect 506 574 508 582
rect 516 574 518 582
rect 536 574 538 582
rect 546 574 548 582
rect 566 574 568 582
rect 576 574 578 582
rect 586 574 588 582
rect 596 574 600 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 102 572 114 574
rect 0 564 4 572
rect 12 564 14 572
rect 22 564 24 572
rect 42 564 44 572
rect 52 564 54 572
rect 72 564 74 572
rect 82 564 84 572
rect 102 564 104 572
rect 112 564 114 572
rect 132 572 144 574
rect 132 564 134 572
rect 142 564 144 572
rect 162 572 174 574
rect 162 564 164 572
rect 172 564 174 572
rect 192 572 204 574
rect 192 564 194 572
rect 202 564 204 572
rect 222 572 234 574
rect 222 564 224 572
rect 232 564 234 572
rect 242 572 256 574
rect 242 564 244 572
rect 252 564 256 572
rect 264 572 276 574
rect 264 564 266 572
rect 274 564 276 572
rect 294 572 306 574
rect 294 564 296 572
rect 304 564 306 572
rect 324 572 336 574
rect 324 564 326 572
rect 334 564 336 572
rect 344 572 358 574
rect 344 564 348 572
rect 356 564 358 572
rect 366 572 378 574
rect 366 564 368 572
rect 376 564 378 572
rect 396 572 408 574
rect 396 564 398 572
rect 406 564 408 572
rect 426 572 438 574
rect 426 564 428 572
rect 436 564 438 572
rect 456 572 468 574
rect 456 564 458 572
rect 466 564 468 572
rect 486 572 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 486 564 488 572
rect 496 564 498 572
rect 516 564 518 572
rect 526 564 528 572
rect 546 564 548 572
rect 556 564 558 572
rect 576 564 578 572
rect 586 564 588 572
rect 596 564 600 572
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 192 562 214 564
rect 222 562 286 564
rect 294 562 316 564
rect 324 562 378 564
rect 386 562 408 564
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 0 554 4 562
rect 12 554 14 562
rect 22 554 24 562
rect 32 554 34 562
rect 52 554 54 562
rect 62 554 64 562
rect 82 554 84 562
rect 92 554 94 562
rect 112 554 114 562
rect 122 554 124 562
rect 142 554 144 562
rect 152 554 154 562
rect 172 554 174 562
rect 182 554 184 562
rect 202 554 204 562
rect 212 554 214 562
rect 232 554 234 562
rect 242 554 244 562
rect 252 554 256 562
rect 264 554 266 562
rect 274 554 276 562
rect 284 554 286 562
rect 304 554 306 562
rect 314 554 316 562
rect 334 554 336 562
rect 344 554 348 562
rect 356 554 358 562
rect 366 554 368 562
rect 386 554 388 562
rect 396 554 398 562
rect 416 554 418 562
rect 426 554 428 562
rect 446 554 448 562
rect 456 554 458 562
rect 476 554 478 562
rect 486 554 488 562
rect 506 554 508 562
rect 516 554 518 562
rect 536 554 538 562
rect 546 554 548 562
rect 566 554 568 562
rect 576 554 578 562
rect 586 554 588 562
rect 596 554 600 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 192 552 214 554
rect 222 552 286 554
rect 294 552 316 554
rect 324 552 378 554
rect 386 552 408 554
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 0 544 4 552
rect 12 544 14 552
rect 22 544 24 552
rect 42 544 44 552
rect 52 544 54 552
rect 72 544 74 552
rect 82 544 84 552
rect 102 544 104 552
rect 112 544 114 552
rect 132 544 134 552
rect 142 544 144 552
rect 162 544 164 552
rect 172 544 174 552
rect 192 544 194 552
rect 202 544 204 552
rect 222 544 224 552
rect 232 544 234 552
rect 242 544 244 552
rect 252 544 256 552
rect 264 544 266 552
rect 274 544 276 552
rect 294 544 296 552
rect 304 544 306 552
rect 324 544 326 552
rect 334 544 336 552
rect 344 544 348 552
rect 356 544 358 552
rect 366 544 368 552
rect 376 544 378 552
rect 396 544 398 552
rect 406 544 408 552
rect 426 544 428 552
rect 436 544 438 552
rect 456 544 458 552
rect 466 544 468 552
rect 486 544 488 552
rect 496 544 498 552
rect 516 544 518 552
rect 526 544 528 552
rect 546 544 548 552
rect 556 544 558 552
rect 576 544 578 552
rect 586 544 588 552
rect 596 544 600 552
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 192 542 214 544
rect 222 542 286 544
rect 294 542 316 544
rect 324 542 378 544
rect 386 542 408 544
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 0 534 4 542
rect 12 534 14 542
rect 22 534 24 542
rect 32 534 34 542
rect 52 534 54 542
rect 62 534 64 542
rect 82 534 84 542
rect 92 534 94 542
rect 112 534 114 542
rect 122 534 124 542
rect 142 534 144 542
rect 152 534 154 542
rect 172 534 174 542
rect 182 534 184 542
rect 202 534 204 542
rect 212 534 214 542
rect 232 534 234 542
rect 242 534 244 542
rect 252 534 256 542
rect 264 534 266 542
rect 274 534 276 542
rect 284 534 286 542
rect 304 534 306 542
rect 314 534 316 542
rect 334 534 336 542
rect 344 534 348 542
rect 356 534 358 542
rect 366 534 368 542
rect 386 534 388 542
rect 396 534 398 542
rect 416 534 418 542
rect 426 534 428 542
rect 446 534 448 542
rect 456 534 458 542
rect 476 534 478 542
rect 486 534 488 542
rect 506 534 508 542
rect 516 534 518 542
rect 536 534 538 542
rect 546 534 548 542
rect 566 534 568 542
rect 576 534 578 542
rect 586 534 588 542
rect 596 534 600 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 192 532 214 534
rect 222 532 286 534
rect 294 532 316 534
rect 324 532 378 534
rect 386 532 408 534
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 0 524 4 532
rect 12 524 14 532
rect 22 524 24 532
rect 42 524 44 532
rect 52 524 54 532
rect 72 524 74 532
rect 82 524 84 532
rect 102 524 104 532
rect 112 524 114 532
rect 132 524 134 532
rect 142 524 144 532
rect 162 524 164 532
rect 172 524 174 532
rect 192 524 194 532
rect 202 524 204 532
rect 222 524 224 532
rect 232 524 234 532
rect 242 524 244 532
rect 252 524 256 532
rect 264 524 266 532
rect 274 524 276 532
rect 294 524 296 532
rect 304 524 306 532
rect 324 524 326 532
rect 334 524 336 532
rect 344 524 348 532
rect 356 524 358 532
rect 366 524 368 532
rect 376 524 378 532
rect 396 524 398 532
rect 406 524 408 532
rect 426 524 428 532
rect 436 524 438 532
rect 456 524 458 532
rect 466 524 468 532
rect 486 524 488 532
rect 496 524 498 532
rect 516 524 518 532
rect 526 524 528 532
rect 546 524 548 532
rect 556 524 558 532
rect 576 524 578 532
rect 586 524 588 532
rect 596 524 600 532
rect 0 516 600 524
rect 0 8 4 516
rect 12 508 14 516
rect 22 508 24 516
rect 32 508 34 516
rect 42 508 44 516
rect 52 508 54 516
rect 62 508 64 516
rect 72 508 74 516
rect 82 508 84 516
rect 92 508 94 516
rect 102 508 104 516
rect 112 508 114 516
rect 122 508 124 516
rect 132 508 134 516
rect 142 508 144 516
rect 152 508 154 516
rect 162 508 164 516
rect 172 508 174 516
rect 182 508 184 516
rect 192 508 194 516
rect 202 508 204 516
rect 212 508 214 516
rect 222 508 224 516
rect 232 508 234 516
rect 242 508 244 516
rect 252 508 254 516
rect 262 508 264 516
rect 272 508 274 516
rect 282 508 284 516
rect 292 508 294 516
rect 302 508 308 516
rect 316 508 318 516
rect 326 508 328 516
rect 336 508 338 516
rect 346 508 348 516
rect 356 508 358 516
rect 366 508 368 516
rect 376 508 378 516
rect 386 508 388 516
rect 396 508 398 516
rect 406 508 408 516
rect 416 508 418 516
rect 426 508 428 516
rect 436 508 438 516
rect 446 508 448 516
rect 456 508 458 516
rect 466 508 468 516
rect 476 508 478 516
rect 486 508 488 516
rect 496 508 498 516
rect 506 508 508 516
rect 516 508 518 516
rect 526 508 528 516
rect 536 508 538 516
rect 546 508 548 516
rect 556 508 558 516
rect 566 508 568 516
rect 576 508 578 516
rect 12 506 588 508
rect 12 502 198 506
rect 12 14 16 502
rect 28 484 198 490
rect 28 456 38 484
rect 56 456 78 466
rect 196 456 198 484
rect 28 454 198 456
rect 28 446 38 454
rect 56 452 198 454
rect 56 446 82 452
rect 28 444 82 446
rect 190 444 198 452
rect 28 436 38 444
rect 56 436 198 444
rect 28 434 198 436
rect 28 426 38 434
rect 56 432 198 434
rect 56 426 64 432
rect 28 424 64 426
rect 28 416 38 424
rect 56 416 64 424
rect 28 414 64 416
rect 28 406 38 414
rect 56 406 64 414
rect 28 404 64 406
rect 28 396 38 404
rect 56 396 64 404
rect 28 394 64 396
rect 28 386 38 394
rect 56 386 64 394
rect 28 384 64 386
rect 28 376 38 384
rect 56 376 64 384
rect 28 374 64 376
rect 28 366 38 374
rect 56 366 64 374
rect 28 364 64 366
rect 28 356 38 364
rect 56 356 64 364
rect 28 354 64 356
rect 28 346 38 354
rect 56 346 64 354
rect 28 344 64 346
rect 28 336 38 344
rect 56 336 64 344
rect 28 334 64 336
rect 28 326 38 334
rect 56 326 64 334
rect 28 324 64 326
rect 28 316 38 324
rect 56 316 64 324
rect 28 314 64 316
rect 28 306 38 314
rect 56 306 64 314
rect 28 304 64 306
rect 28 296 38 304
rect 56 296 64 304
rect 28 294 64 296
rect 28 286 38 294
rect 56 286 64 294
rect 28 284 64 286
rect 28 276 38 284
rect 56 276 64 284
rect 28 274 64 276
rect 28 266 38 274
rect 56 266 64 274
rect 28 264 64 266
rect 28 256 38 264
rect 56 256 64 264
rect 28 254 64 256
rect 28 246 38 254
rect 56 246 64 254
rect 28 244 64 246
rect 28 236 38 244
rect 56 236 64 244
rect 28 234 64 236
rect 28 226 38 234
rect 56 226 64 234
rect 28 224 64 226
rect 28 216 38 224
rect 56 216 64 224
rect 28 214 64 216
rect 28 206 38 214
rect 56 206 64 214
rect 28 204 64 206
rect 28 196 38 204
rect 56 196 64 204
rect 28 194 64 196
rect 28 186 38 194
rect 56 186 64 194
rect 28 184 64 186
rect 28 176 38 184
rect 56 176 64 184
rect 28 174 64 176
rect 28 166 38 174
rect 56 166 64 174
rect 28 164 64 166
rect 28 156 38 164
rect 56 156 64 164
rect 28 154 64 156
rect 28 146 38 154
rect 56 146 64 154
rect 28 144 64 146
rect 28 136 38 144
rect 56 136 64 144
rect 28 134 64 136
rect 28 126 38 134
rect 56 126 64 134
rect 28 124 64 126
rect 28 116 38 124
rect 56 116 64 124
rect 28 114 64 116
rect 28 106 38 114
rect 56 106 64 114
rect 28 104 64 106
rect 28 96 38 104
rect 56 96 64 104
rect 28 94 64 96
rect 28 86 38 94
rect 56 86 64 94
rect 28 84 64 86
rect 72 428 198 432
rect 72 390 78 428
rect 196 420 198 428
rect 204 458 396 506
rect 402 502 588 506
rect 204 414 285 458
rect 72 386 106 390
rect 72 348 78 386
rect 112 398 285 414
rect 315 414 396 458
rect 402 484 572 490
rect 402 456 404 484
rect 522 456 544 466
rect 562 456 572 484
rect 402 454 572 456
rect 402 452 544 454
rect 402 444 410 452
rect 518 446 544 452
rect 562 446 572 454
rect 518 444 572 446
rect 402 436 544 444
rect 562 436 572 444
rect 402 434 572 436
rect 402 432 544 434
rect 402 428 528 432
rect 402 420 404 428
rect 315 398 488 414
rect 240 390 360 398
rect 112 386 488 390
rect 240 378 360 386
rect 112 362 488 378
rect 522 390 528 428
rect 494 386 528 390
rect 236 348 240 356
rect 72 332 240 348
rect 72 324 82 332
rect 72 320 240 324
rect 72 312 82 320
rect 72 296 240 312
rect 72 218 78 296
rect 236 288 240 296
rect 246 282 354 362
rect 360 348 364 356
rect 522 348 528 386
rect 360 332 528 348
rect 518 324 528 332
rect 360 320 528 324
rect 518 312 528 320
rect 360 296 528 312
rect 360 288 364 296
rect 112 274 488 282
rect 112 266 285 274
rect 240 248 285 266
rect 112 238 285 248
rect 315 266 488 274
rect 315 248 360 266
rect 315 238 488 248
rect 112 232 488 238
rect 236 218 240 226
rect 72 202 240 218
rect 72 194 82 202
rect 72 190 240 194
rect 72 182 82 190
rect 72 166 240 182
rect 72 88 78 166
rect 236 158 240 166
rect 246 152 354 232
rect 360 218 364 226
rect 522 218 528 296
rect 360 202 528 218
rect 518 194 528 202
rect 360 190 528 194
rect 518 182 528 190
rect 360 166 528 182
rect 360 158 364 166
rect 112 138 488 152
rect 112 136 285 138
rect 240 118 285 136
rect 315 136 488 138
rect 112 102 285 118
rect 196 88 198 96
rect 72 84 198 88
rect 28 76 38 84
rect 56 76 198 84
rect 28 74 198 76
rect 28 66 38 74
rect 56 72 198 74
rect 56 66 82 72
rect 28 64 82 66
rect 190 64 198 72
rect 28 56 38 64
rect 56 56 78 64
rect 196 56 198 64
rect 28 54 78 56
rect 28 46 38 54
rect 66 46 68 54
rect 76 46 78 54
rect 86 54 98 56
rect 86 46 88 54
rect 96 46 98 54
rect 106 54 118 56
rect 106 46 108 54
rect 116 46 118 54
rect 126 54 138 56
rect 126 46 128 54
rect 136 46 138 54
rect 146 54 158 56
rect 146 46 148 54
rect 156 46 158 54
rect 166 54 178 56
rect 166 46 168 54
rect 176 46 178 54
rect 186 54 198 56
rect 186 46 188 54
rect 196 46 198 54
rect 28 44 198 46
rect 28 36 38 44
rect 66 36 68 44
rect 76 36 78 44
rect 86 36 88 44
rect 96 36 98 44
rect 106 36 108 44
rect 116 36 118 44
rect 126 36 128 44
rect 136 36 138 44
rect 146 36 148 44
rect 156 36 158 44
rect 166 36 168 44
rect 176 36 178 44
rect 186 36 188 44
rect 196 36 198 44
rect 28 26 198 36
rect 204 54 285 102
rect 315 118 360 136
rect 315 102 488 118
rect 315 54 396 102
rect 12 12 198 14
rect 0 4 14 8
rect 182 4 198 12
rect 0 -2 198 4
rect 204 -2 396 54
rect 402 88 404 96
rect 522 88 528 166
rect 402 84 528 88
rect 536 426 544 432
rect 562 426 572 434
rect 536 424 572 426
rect 536 416 544 424
rect 562 416 572 424
rect 536 414 572 416
rect 536 406 544 414
rect 562 406 572 414
rect 536 404 572 406
rect 536 396 544 404
rect 562 396 572 404
rect 536 394 572 396
rect 536 386 544 394
rect 562 386 572 394
rect 536 384 572 386
rect 536 376 544 384
rect 562 376 572 384
rect 536 374 572 376
rect 536 366 544 374
rect 562 366 572 374
rect 536 364 572 366
rect 536 356 544 364
rect 562 356 572 364
rect 536 354 572 356
rect 536 346 544 354
rect 562 346 572 354
rect 536 344 572 346
rect 536 336 544 344
rect 562 336 572 344
rect 536 334 572 336
rect 536 326 544 334
rect 562 326 572 334
rect 536 324 572 326
rect 536 316 544 324
rect 562 316 572 324
rect 536 314 572 316
rect 536 306 544 314
rect 562 306 572 314
rect 536 304 572 306
rect 536 296 544 304
rect 562 296 572 304
rect 536 294 572 296
rect 536 286 544 294
rect 562 286 572 294
rect 536 284 572 286
rect 536 276 544 284
rect 562 276 572 284
rect 536 274 572 276
rect 536 266 544 274
rect 562 266 572 274
rect 536 264 572 266
rect 536 256 544 264
rect 562 256 572 264
rect 536 254 572 256
rect 536 246 544 254
rect 562 246 572 254
rect 536 244 572 246
rect 536 236 544 244
rect 562 236 572 244
rect 536 234 572 236
rect 536 226 544 234
rect 562 226 572 234
rect 536 224 572 226
rect 536 216 544 224
rect 562 216 572 224
rect 536 214 572 216
rect 536 206 544 214
rect 562 206 572 214
rect 536 204 572 206
rect 536 196 544 204
rect 562 196 572 204
rect 536 194 572 196
rect 536 186 544 194
rect 562 186 572 194
rect 536 184 572 186
rect 536 176 544 184
rect 562 176 572 184
rect 536 174 572 176
rect 536 166 544 174
rect 562 166 572 174
rect 536 164 572 166
rect 536 156 544 164
rect 562 156 572 164
rect 536 154 572 156
rect 536 146 544 154
rect 562 146 572 154
rect 536 144 572 146
rect 536 136 544 144
rect 562 136 572 144
rect 536 134 572 136
rect 536 126 544 134
rect 562 126 572 134
rect 536 124 572 126
rect 536 116 544 124
rect 562 116 572 124
rect 536 114 572 116
rect 536 106 544 114
rect 562 106 572 114
rect 536 104 572 106
rect 536 96 544 104
rect 562 96 572 104
rect 536 94 572 96
rect 536 86 544 94
rect 562 86 572 94
rect 536 84 572 86
rect 402 76 544 84
rect 562 76 572 84
rect 402 74 572 76
rect 402 72 544 74
rect 402 64 410 72
rect 518 66 544 72
rect 562 66 572 74
rect 518 64 572 66
rect 402 56 404 64
rect 522 56 544 64
rect 562 56 572 64
rect 402 54 414 56
rect 402 46 404 54
rect 412 46 414 54
rect 422 54 434 56
rect 422 46 424 54
rect 432 46 434 54
rect 442 54 454 56
rect 442 46 444 54
rect 452 46 454 54
rect 462 54 474 56
rect 462 46 464 54
rect 472 46 474 54
rect 482 54 494 56
rect 482 46 484 54
rect 492 46 494 54
rect 502 54 514 56
rect 502 46 504 54
rect 512 46 514 54
rect 522 54 572 56
rect 522 46 524 54
rect 532 46 534 54
rect 562 46 572 54
rect 402 44 572 46
rect 402 36 404 44
rect 412 36 414 44
rect 422 36 424 44
rect 432 36 434 44
rect 442 36 444 44
rect 452 36 454 44
rect 462 36 464 44
rect 472 36 474 44
rect 482 36 484 44
rect 492 36 494 44
rect 502 36 504 44
rect 512 36 514 44
rect 522 36 524 44
rect 532 36 534 44
rect 562 36 572 44
rect 402 26 572 36
rect 584 14 588 502
rect 402 12 588 14
rect 402 4 408 12
rect 596 8 600 516
rect 586 4 600 8
rect 402 -2 600 4
<< m2contact >>
rect 56 1290 64 1298
rect 86 1290 94 1298
rect 116 1290 124 1298
rect 146 1290 154 1298
rect 176 1290 184 1298
rect 206 1290 214 1298
rect 236 1290 244 1298
rect 266 1290 274 1298
rect 296 1290 304 1298
rect 326 1290 334 1298
rect 356 1290 364 1298
rect 386 1290 394 1298
rect 416 1290 424 1298
rect 446 1290 454 1298
rect 476 1290 484 1298
rect 506 1290 514 1298
rect 536 1290 544 1298
rect 46 1280 54 1288
rect 66 1280 74 1288
rect 96 1280 104 1288
rect 126 1280 134 1288
rect 156 1280 164 1288
rect 186 1280 194 1288
rect 216 1280 224 1288
rect 246 1280 254 1288
rect 276 1280 284 1288
rect 306 1280 314 1288
rect 336 1280 344 1288
rect 366 1280 374 1288
rect 396 1280 404 1288
rect 426 1280 434 1288
rect 456 1280 464 1288
rect 486 1280 494 1288
rect 516 1280 524 1288
rect 546 1280 554 1288
rect 56 1270 64 1278
rect 86 1270 94 1278
rect 116 1270 124 1278
rect 146 1270 154 1278
rect 176 1270 184 1278
rect 206 1270 214 1278
rect 236 1270 244 1278
rect 266 1270 274 1278
rect 296 1270 304 1278
rect 326 1270 334 1278
rect 356 1270 364 1278
rect 386 1270 394 1278
rect 416 1270 424 1278
rect 446 1270 454 1278
rect 476 1270 484 1278
rect 506 1270 514 1278
rect 536 1270 544 1278
rect 46 1260 54 1268
rect 66 1260 74 1268
rect 96 1260 104 1268
rect 126 1260 134 1268
rect 156 1260 164 1268
rect 186 1260 194 1268
rect 216 1260 224 1268
rect 246 1260 254 1268
rect 276 1260 284 1268
rect 306 1260 314 1268
rect 336 1260 344 1268
rect 366 1260 374 1268
rect 396 1260 404 1268
rect 426 1260 434 1268
rect 456 1260 464 1268
rect 486 1260 494 1268
rect 516 1260 524 1268
rect 546 1260 554 1268
rect 56 1250 64 1258
rect 86 1250 94 1258
rect 116 1250 124 1258
rect 146 1250 154 1258
rect 176 1250 184 1258
rect 206 1250 214 1258
rect 236 1250 244 1258
rect 266 1250 274 1258
rect 296 1250 304 1258
rect 326 1250 334 1258
rect 356 1250 364 1258
rect 386 1250 394 1258
rect 416 1250 424 1258
rect 446 1250 454 1258
rect 476 1250 484 1258
rect 506 1250 514 1258
rect 536 1250 544 1258
rect 46 1240 54 1248
rect 66 1240 74 1248
rect 96 1240 104 1248
rect 126 1240 134 1248
rect 156 1240 164 1248
rect 186 1240 194 1248
rect 216 1240 224 1248
rect 246 1240 254 1248
rect 276 1240 284 1248
rect 306 1240 314 1248
rect 336 1240 344 1248
rect 366 1240 374 1248
rect 396 1240 404 1248
rect 426 1240 434 1248
rect 456 1240 464 1248
rect 486 1240 494 1248
rect 516 1240 524 1248
rect 546 1240 554 1248
rect 56 1230 64 1238
rect 86 1230 94 1238
rect 116 1230 124 1238
rect 146 1230 154 1238
rect 176 1230 184 1238
rect 206 1230 214 1238
rect 236 1230 244 1238
rect 266 1230 274 1238
rect 296 1230 304 1238
rect 326 1230 334 1238
rect 356 1230 364 1238
rect 386 1230 394 1238
rect 416 1230 424 1238
rect 446 1230 454 1238
rect 476 1230 484 1238
rect 506 1230 514 1238
rect 536 1230 544 1238
rect 46 1220 54 1228
rect 66 1220 74 1228
rect 96 1220 104 1228
rect 126 1220 134 1228
rect 156 1220 164 1228
rect 186 1220 194 1228
rect 216 1220 224 1228
rect 246 1220 254 1228
rect 276 1220 284 1228
rect 306 1220 314 1228
rect 336 1220 344 1228
rect 366 1220 374 1228
rect 396 1220 404 1228
rect 426 1220 434 1228
rect 456 1220 464 1228
rect 486 1220 494 1228
rect 516 1220 524 1228
rect 546 1220 554 1228
rect 56 1210 64 1218
rect 86 1210 94 1218
rect 116 1210 124 1218
rect 146 1210 154 1218
rect 176 1210 184 1218
rect 206 1210 214 1218
rect 236 1210 244 1218
rect 266 1210 274 1218
rect 296 1210 304 1218
rect 326 1210 334 1218
rect 356 1210 364 1218
rect 386 1210 394 1218
rect 416 1210 424 1218
rect 446 1210 454 1218
rect 476 1210 484 1218
rect 506 1210 514 1218
rect 536 1210 544 1218
rect 46 1200 54 1208
rect 66 1200 74 1208
rect 96 1200 104 1208
rect 126 1200 134 1208
rect 156 1200 164 1208
rect 186 1200 194 1208
rect 216 1200 224 1208
rect 246 1200 254 1208
rect 276 1200 284 1208
rect 306 1200 314 1208
rect 336 1200 344 1208
rect 366 1200 374 1208
rect 396 1200 404 1208
rect 426 1200 434 1208
rect 456 1200 464 1208
rect 486 1200 494 1208
rect 516 1200 524 1208
rect 546 1200 554 1208
rect 56 1190 64 1198
rect 86 1190 94 1198
rect 116 1190 124 1198
rect 146 1190 154 1198
rect 176 1190 184 1198
rect 206 1190 214 1198
rect 236 1190 244 1198
rect 266 1190 274 1198
rect 296 1190 304 1198
rect 326 1190 334 1198
rect 356 1190 364 1198
rect 386 1190 394 1198
rect 416 1190 424 1198
rect 446 1190 454 1198
rect 476 1190 484 1198
rect 506 1190 514 1198
rect 536 1190 544 1198
rect 46 1180 54 1188
rect 66 1180 74 1188
rect 516 1180 524 1188
rect 546 1180 554 1188
rect 56 1170 64 1178
rect 86 1170 94 1178
rect 116 1170 124 1178
rect 146 1170 154 1178
rect 176 1170 184 1178
rect 206 1170 214 1178
rect 236 1170 244 1178
rect 266 1170 274 1178
rect 296 1170 304 1178
rect 326 1170 334 1178
rect 356 1170 364 1178
rect 386 1170 394 1178
rect 416 1170 424 1178
rect 446 1170 454 1178
rect 476 1170 484 1178
rect 506 1170 514 1178
rect 536 1170 544 1178
rect 46 1160 54 1168
rect 66 1160 74 1168
rect 96 1160 104 1168
rect 126 1160 134 1168
rect 156 1160 164 1168
rect 186 1160 194 1168
rect 216 1160 224 1168
rect 246 1160 254 1168
rect 276 1160 284 1168
rect 306 1160 314 1168
rect 336 1160 344 1168
rect 366 1160 374 1168
rect 396 1160 404 1168
rect 426 1160 434 1168
rect 456 1160 464 1168
rect 486 1160 494 1168
rect 516 1160 524 1168
rect 546 1160 554 1168
rect 56 1150 64 1158
rect 86 1150 94 1158
rect 116 1150 124 1158
rect 146 1150 154 1158
rect 176 1150 184 1158
rect 206 1150 214 1158
rect 236 1150 244 1158
rect 266 1150 274 1158
rect 296 1150 304 1158
rect 326 1150 334 1158
rect 356 1150 364 1158
rect 386 1150 394 1158
rect 416 1150 424 1158
rect 446 1150 454 1158
rect 476 1150 484 1158
rect 506 1150 514 1158
rect 536 1150 544 1158
rect 46 1140 54 1148
rect 66 1140 74 1148
rect 96 1140 104 1148
rect 126 1140 134 1148
rect 156 1140 164 1148
rect 186 1140 194 1148
rect 216 1140 224 1148
rect 246 1140 254 1148
rect 276 1140 284 1148
rect 306 1140 314 1148
rect 336 1140 344 1148
rect 366 1140 374 1148
rect 396 1140 404 1148
rect 426 1140 434 1148
rect 456 1140 464 1148
rect 486 1140 494 1148
rect 516 1140 524 1148
rect 546 1140 554 1148
rect 56 1130 64 1138
rect 86 1130 94 1138
rect 116 1130 124 1138
rect 146 1130 154 1138
rect 176 1130 184 1138
rect 206 1130 214 1138
rect 236 1130 244 1138
rect 266 1130 274 1138
rect 296 1130 304 1138
rect 326 1130 334 1138
rect 356 1130 364 1138
rect 386 1130 394 1138
rect 416 1130 424 1138
rect 446 1130 454 1138
rect 476 1130 484 1138
rect 506 1130 514 1138
rect 536 1130 544 1138
rect 46 1120 54 1128
rect 66 1120 74 1128
rect 96 1120 104 1128
rect 126 1120 134 1128
rect 156 1120 164 1128
rect 186 1120 194 1128
rect 216 1120 224 1128
rect 246 1120 254 1128
rect 276 1120 284 1128
rect 306 1120 314 1128
rect 336 1120 344 1128
rect 366 1120 374 1128
rect 396 1120 404 1128
rect 426 1120 434 1128
rect 456 1120 464 1128
rect 486 1120 494 1128
rect 56 1110 64 1118
rect 76 1110 84 1118
rect 46 1100 54 1108
rect 66 1100 74 1108
rect 96 1100 104 1108
rect 126 1100 134 1108
rect 156 1100 164 1108
rect 186 1100 194 1108
rect 216 1100 224 1108
rect 246 1100 254 1108
rect 276 1100 284 1108
rect 306 1100 314 1108
rect 336 1100 344 1108
rect 366 1100 374 1108
rect 396 1100 404 1108
rect 426 1100 434 1108
rect 456 1100 464 1108
rect 486 1100 494 1108
rect 516 1100 524 1128
rect 546 1120 554 1128
rect 536 1110 544 1118
rect 546 1100 554 1108
rect 56 1090 64 1098
rect 86 1090 94 1098
rect 116 1090 124 1098
rect 146 1090 154 1098
rect 176 1090 184 1098
rect 206 1090 214 1098
rect 236 1090 244 1098
rect 266 1090 274 1098
rect 296 1090 304 1098
rect 326 1090 334 1098
rect 356 1090 364 1098
rect 386 1090 394 1098
rect 416 1090 424 1098
rect 446 1090 454 1098
rect 476 1090 484 1098
rect 506 1090 514 1098
rect 536 1090 544 1098
rect 46 1080 54 1088
rect 66 1080 74 1088
rect 96 1080 104 1088
rect 126 1080 134 1088
rect 156 1080 164 1088
rect 186 1080 194 1088
rect 216 1080 224 1088
rect 246 1080 254 1088
rect 276 1080 284 1088
rect 306 1080 314 1088
rect 336 1080 344 1088
rect 366 1080 374 1088
rect 396 1080 404 1088
rect 426 1080 434 1088
rect 456 1080 464 1088
rect 486 1080 494 1088
rect 516 1080 524 1088
rect 546 1080 554 1088
rect 56 1070 64 1078
rect 86 1070 94 1078
rect 116 1070 124 1078
rect 146 1070 154 1078
rect 176 1070 184 1078
rect 206 1070 214 1078
rect 236 1070 244 1078
rect 266 1070 274 1078
rect 296 1070 304 1078
rect 326 1070 334 1078
rect 356 1070 364 1078
rect 386 1070 394 1078
rect 416 1070 424 1078
rect 446 1070 454 1078
rect 476 1070 484 1078
rect 506 1070 514 1078
rect 536 1070 544 1078
rect 46 1060 54 1068
rect 66 1060 74 1068
rect 96 1060 104 1068
rect 126 1060 134 1068
rect 156 1060 164 1068
rect 186 1060 194 1068
rect 216 1060 224 1068
rect 246 1060 254 1068
rect 276 1060 284 1068
rect 306 1060 314 1068
rect 336 1060 344 1068
rect 366 1060 374 1068
rect 396 1060 404 1068
rect 426 1060 434 1068
rect 456 1060 464 1068
rect 486 1060 494 1068
rect 516 1060 524 1068
rect 546 1060 554 1068
rect 56 1050 64 1058
rect 86 1050 94 1058
rect 116 1050 124 1058
rect 146 1050 154 1058
rect 176 1050 184 1058
rect 206 1050 214 1058
rect 236 1050 244 1058
rect 266 1050 274 1058
rect 296 1050 304 1058
rect 326 1050 334 1058
rect 356 1050 364 1058
rect 386 1050 394 1058
rect 416 1050 424 1058
rect 446 1050 454 1058
rect 476 1050 484 1058
rect 506 1050 514 1058
rect 536 1050 544 1058
rect 46 1040 54 1048
rect 66 1040 74 1048
rect 96 1040 104 1048
rect 126 1040 134 1048
rect 156 1040 164 1048
rect 186 1040 194 1048
rect 216 1040 224 1048
rect 246 1040 254 1048
rect 276 1040 284 1048
rect 306 1040 314 1048
rect 336 1040 344 1048
rect 366 1040 374 1048
rect 396 1040 404 1048
rect 426 1040 434 1048
rect 456 1040 464 1048
rect 486 1040 494 1048
rect 56 1030 64 1038
rect 86 1030 94 1038
rect 46 1020 54 1028
rect 66 1020 74 1028
rect 96 1020 104 1028
rect 126 1020 134 1028
rect 156 1020 164 1028
rect 186 1020 194 1028
rect 216 1020 224 1028
rect 246 1020 254 1028
rect 276 1020 284 1028
rect 306 1020 314 1028
rect 336 1020 344 1028
rect 366 1020 374 1028
rect 396 1020 404 1028
rect 426 1020 434 1028
rect 456 1020 464 1028
rect 486 1020 494 1028
rect 516 1020 524 1048
rect 546 1040 554 1048
rect 536 1030 544 1038
rect 546 1020 554 1028
rect 56 1010 64 1018
rect 86 1010 94 1018
rect 116 1010 124 1018
rect 146 1010 154 1018
rect 176 1010 184 1018
rect 206 1010 214 1018
rect 236 1010 244 1018
rect 266 1010 274 1018
rect 296 1010 304 1018
rect 326 1010 334 1018
rect 356 1010 364 1018
rect 386 1010 394 1018
rect 416 1010 424 1018
rect 446 1010 454 1018
rect 476 1010 484 1018
rect 506 1010 514 1018
rect 536 1010 544 1018
rect 46 1000 54 1008
rect 66 1000 74 1008
rect 96 1000 104 1008
rect 126 1000 134 1008
rect 156 1000 164 1008
rect 186 1000 194 1008
rect 216 1000 224 1008
rect 246 1000 254 1008
rect 276 1000 284 1008
rect 306 1000 314 1008
rect 336 1000 344 1008
rect 366 1000 374 1008
rect 396 1000 404 1008
rect 426 1000 434 1008
rect 456 1000 464 1008
rect 486 1000 494 1008
rect 516 1000 524 1008
rect 546 1000 554 1008
rect 56 990 64 998
rect 86 990 94 998
rect 116 990 124 998
rect 146 990 154 998
rect 176 990 184 998
rect 206 990 214 998
rect 236 990 244 998
rect 266 990 274 998
rect 296 990 304 998
rect 326 990 334 998
rect 356 990 364 998
rect 386 990 394 998
rect 416 990 424 998
rect 446 990 454 998
rect 476 990 484 998
rect 506 990 514 998
rect 536 990 544 998
rect 46 980 54 988
rect 66 980 74 988
rect 96 980 104 988
rect 126 980 134 988
rect 156 980 164 988
rect 186 980 194 988
rect 216 980 224 988
rect 246 980 254 988
rect 276 980 284 988
rect 306 980 314 988
rect 336 980 344 988
rect 366 980 374 988
rect 396 980 404 988
rect 426 980 434 988
rect 456 980 464 988
rect 486 980 494 988
rect 516 980 524 988
rect 546 980 554 988
rect 56 970 64 978
rect 86 970 94 978
rect 116 970 124 978
rect 146 970 154 978
rect 176 970 184 978
rect 206 970 214 978
rect 236 970 244 978
rect 266 970 274 978
rect 296 970 304 978
rect 326 970 334 978
rect 356 970 364 978
rect 386 970 394 978
rect 416 970 424 978
rect 446 970 454 978
rect 476 970 484 978
rect 506 970 514 978
rect 536 970 544 978
rect 46 960 54 968
rect 546 960 554 968
rect 56 950 64 958
rect 86 950 94 958
rect 116 950 124 958
rect 146 950 154 958
rect 176 950 184 958
rect 206 950 214 958
rect 236 950 244 958
rect 266 950 274 958
rect 296 950 304 958
rect 326 950 334 958
rect 356 950 364 958
rect 386 950 394 958
rect 416 950 424 958
rect 446 950 454 958
rect 476 950 484 958
rect 506 950 514 958
rect 536 950 544 958
rect 46 940 54 948
rect 66 940 74 948
rect 96 940 104 948
rect 126 940 134 948
rect 156 940 164 948
rect 186 940 194 948
rect 216 940 224 948
rect 246 940 254 948
rect 276 940 284 948
rect 306 940 314 948
rect 336 940 344 948
rect 366 940 374 948
rect 396 940 404 948
rect 426 940 434 948
rect 456 940 464 948
rect 486 940 494 948
rect 516 940 524 948
rect 546 940 554 948
rect 56 930 64 938
rect 86 930 94 938
rect 116 930 124 938
rect 146 930 154 938
rect 176 930 184 938
rect 206 930 214 938
rect 236 930 244 938
rect 266 930 274 938
rect 296 930 304 938
rect 326 930 334 938
rect 356 930 364 938
rect 386 930 394 938
rect 416 930 424 938
rect 446 930 454 938
rect 476 930 484 938
rect 506 930 514 938
rect 536 930 544 938
rect 46 920 54 928
rect 66 920 74 928
rect 96 920 104 928
rect 126 920 134 928
rect 156 920 164 928
rect 186 920 194 928
rect 216 920 224 928
rect 246 920 254 928
rect 276 920 284 928
rect 306 920 314 928
rect 336 920 344 928
rect 366 920 374 928
rect 396 920 404 928
rect 426 920 434 928
rect 456 920 464 928
rect 486 920 494 928
rect 516 920 524 928
rect 546 920 554 928
rect 56 910 64 918
rect 86 910 94 918
rect 116 910 124 918
rect 146 910 154 918
rect 176 910 184 918
rect 206 910 214 918
rect 236 910 244 918
rect 266 910 274 918
rect 296 910 304 918
rect 326 910 334 918
rect 356 910 364 918
rect 386 910 394 918
rect 416 910 424 918
rect 446 910 454 918
rect 476 910 484 918
rect 506 910 514 918
rect 536 910 544 918
rect 46 900 54 908
rect 66 900 74 908
rect 96 900 104 908
rect 126 900 134 908
rect 156 900 164 908
rect 186 900 194 908
rect 216 900 224 908
rect 246 900 254 908
rect 276 900 284 908
rect 306 900 314 908
rect 336 900 344 908
rect 366 900 374 908
rect 396 900 404 908
rect 426 900 434 908
rect 456 900 464 908
rect 486 900 494 908
rect 516 900 524 908
rect 546 900 554 908
rect 56 890 64 898
rect 86 890 94 898
rect 116 890 124 898
rect 146 890 154 898
rect 176 890 184 898
rect 206 890 214 898
rect 236 890 244 898
rect 266 890 274 898
rect 296 890 304 898
rect 326 890 334 898
rect 356 890 364 898
rect 386 890 394 898
rect 416 890 424 898
rect 446 890 454 898
rect 476 890 484 898
rect 506 890 514 898
rect 536 890 544 898
rect 46 880 54 888
rect 66 880 74 888
rect 96 880 104 888
rect 126 880 134 888
rect 156 880 164 888
rect 186 880 194 888
rect 216 880 224 888
rect 246 880 254 888
rect 276 880 284 888
rect 306 880 314 888
rect 336 880 344 888
rect 366 880 374 888
rect 396 880 404 888
rect 426 880 434 888
rect 456 880 464 888
rect 486 880 494 888
rect 516 880 524 888
rect 546 880 554 888
rect 14 828 22 836
rect 44 828 52 836
rect 74 828 82 836
rect 104 828 112 836
rect 134 828 142 836
rect 164 828 172 836
rect 184 828 192 836
rect 4 818 12 826
rect 24 818 32 826
rect 54 818 62 826
rect 84 818 92 826
rect 114 818 122 826
rect 144 818 152 826
rect 174 818 182 826
rect 14 808 22 816
rect 44 808 52 816
rect 74 808 82 816
rect 104 808 112 816
rect 134 808 142 816
rect 164 808 172 816
rect 184 808 192 816
rect 4 798 12 806
rect 24 798 32 806
rect 54 798 62 806
rect 84 798 92 806
rect 114 798 122 806
rect 144 798 152 806
rect 174 798 182 806
rect 14 788 22 796
rect 44 788 52 796
rect 74 788 82 796
rect 104 788 112 796
rect 134 788 142 796
rect 164 788 172 796
rect 184 788 192 796
rect 4 778 12 786
rect 24 778 32 786
rect 54 778 62 786
rect 84 778 92 786
rect 114 778 122 786
rect 144 778 152 786
rect 174 778 182 786
rect 14 768 22 776
rect 44 768 52 776
rect 74 768 82 776
rect 4 758 12 766
rect 24 758 32 766
rect 54 758 62 766
rect 84 758 92 766
rect 114 758 122 766
rect 144 758 152 766
rect 174 758 182 766
rect 14 748 22 756
rect 44 748 52 756
rect 74 748 82 756
rect 104 748 112 756
rect 134 748 142 756
rect 164 748 172 756
rect 184 748 192 756
rect 4 738 12 746
rect 24 738 32 746
rect 54 738 62 746
rect 84 738 92 746
rect 114 738 122 746
rect 144 738 152 746
rect 174 738 182 746
rect 14 728 22 736
rect 4 718 12 726
rect 24 718 32 726
rect 54 718 62 726
rect 84 718 92 726
rect 114 718 122 726
rect 144 718 152 726
rect 174 718 182 726
rect 14 708 22 716
rect 44 708 52 716
rect 74 708 82 716
rect 104 708 112 716
rect 134 708 142 716
rect 164 708 172 716
rect 184 708 192 716
rect 4 698 12 706
rect 24 698 32 706
rect 54 698 62 706
rect 84 698 92 706
rect 114 698 122 706
rect 144 698 152 706
rect 174 698 182 706
rect 14 688 22 696
rect 44 688 52 696
rect 74 688 82 696
rect 104 688 112 696
rect 134 688 142 696
rect 164 688 172 696
rect 184 688 192 696
rect 286 828 294 836
rect 306 828 314 836
rect 296 818 304 826
rect 286 808 294 816
rect 306 808 314 816
rect 296 798 304 806
rect 286 788 294 796
rect 306 788 314 796
rect 296 778 304 786
rect 286 758 294 766
rect 306 758 314 766
rect 296 748 304 756
rect 286 738 294 746
rect 306 738 314 746
rect 296 728 304 736
rect 286 718 294 726
rect 306 718 314 726
rect 296 706 304 716
rect 286 698 314 706
rect 408 828 416 836
rect 428 828 436 836
rect 458 828 466 836
rect 488 828 496 836
rect 518 828 526 836
rect 548 828 556 836
rect 578 828 586 836
rect 418 818 426 826
rect 448 818 456 826
rect 478 818 486 826
rect 508 818 516 826
rect 538 818 546 826
rect 568 818 576 826
rect 588 818 596 826
rect 408 808 416 816
rect 428 808 436 816
rect 458 808 466 816
rect 488 808 496 816
rect 518 808 526 816
rect 548 808 556 816
rect 578 808 586 816
rect 418 798 426 806
rect 448 798 456 806
rect 478 798 486 806
rect 508 798 516 806
rect 538 798 546 806
rect 568 798 576 806
rect 588 798 596 806
rect 408 788 416 796
rect 428 788 436 796
rect 458 788 466 796
rect 488 788 496 796
rect 518 788 526 796
rect 548 788 556 796
rect 578 788 586 796
rect 418 778 426 786
rect 448 778 456 786
rect 478 778 486 786
rect 508 778 516 786
rect 538 778 546 786
rect 568 778 576 786
rect 588 778 596 786
rect 518 768 526 776
rect 548 768 556 776
rect 578 768 586 776
rect 418 758 426 766
rect 448 758 456 766
rect 478 758 486 766
rect 508 758 516 766
rect 538 758 546 766
rect 568 758 576 766
rect 588 758 596 766
rect 408 748 416 756
rect 428 748 436 756
rect 458 748 466 756
rect 488 748 496 756
rect 518 748 526 756
rect 548 748 556 756
rect 578 748 586 756
rect 418 738 426 746
rect 448 738 456 746
rect 478 738 486 746
rect 508 738 516 746
rect 538 738 546 746
rect 568 738 576 746
rect 588 738 596 746
rect 578 728 586 736
rect 418 718 426 726
rect 448 718 456 726
rect 478 718 486 726
rect 508 718 516 726
rect 538 718 546 726
rect 568 718 576 726
rect 588 718 596 726
rect 408 708 416 716
rect 428 708 436 716
rect 458 708 466 716
rect 488 708 496 716
rect 518 708 526 716
rect 548 708 556 716
rect 578 708 586 716
rect 418 698 426 706
rect 448 698 456 706
rect 478 698 486 706
rect 508 698 516 706
rect 538 698 546 706
rect 568 698 576 706
rect 588 698 596 706
rect 408 688 416 696
rect 428 688 436 696
rect 458 688 466 696
rect 488 688 496 696
rect 518 688 526 696
rect 548 688 556 696
rect 578 688 586 696
rect 14 644 22 652
rect 44 644 52 652
rect 74 644 82 652
rect 104 644 112 652
rect 134 644 142 652
rect 164 644 172 652
rect 194 644 202 652
rect 224 644 232 652
rect 244 644 252 652
rect 266 644 274 652
rect 296 644 304 652
rect 326 644 334 652
rect 348 644 356 652
rect 368 644 376 652
rect 398 644 406 652
rect 428 644 436 652
rect 458 644 466 652
rect 488 644 496 652
rect 518 644 526 652
rect 548 644 556 652
rect 578 644 586 652
rect 4 634 12 642
rect 24 634 32 642
rect 54 634 62 642
rect 84 634 92 642
rect 114 634 122 642
rect 144 634 152 642
rect 174 634 182 642
rect 204 634 212 642
rect 234 634 242 642
rect 256 634 264 642
rect 276 634 284 642
rect 306 634 314 642
rect 336 634 344 642
rect 358 634 366 642
rect 388 634 396 642
rect 418 634 426 642
rect 448 634 456 642
rect 478 634 486 642
rect 508 634 516 642
rect 538 634 546 642
rect 568 634 576 642
rect 588 634 596 642
rect 14 624 22 632
rect 44 624 52 632
rect 74 624 82 632
rect 104 624 112 632
rect 134 624 142 632
rect 164 624 172 632
rect 194 624 202 632
rect 224 624 232 632
rect 244 624 252 632
rect 266 624 274 632
rect 296 624 304 632
rect 326 624 334 632
rect 348 624 356 632
rect 368 624 376 632
rect 398 624 406 632
rect 428 624 436 632
rect 458 624 466 632
rect 488 624 496 632
rect 518 624 526 632
rect 548 624 556 632
rect 578 624 586 632
rect 4 614 12 622
rect 24 614 32 622
rect 54 614 62 622
rect 84 614 92 622
rect 114 614 122 622
rect 144 614 152 622
rect 174 614 182 622
rect 204 614 212 622
rect 234 614 242 622
rect 256 614 264 622
rect 276 614 284 622
rect 306 614 314 622
rect 336 614 344 622
rect 358 614 366 622
rect 388 614 396 622
rect 418 614 426 622
rect 448 614 456 622
rect 478 614 486 622
rect 508 614 516 622
rect 538 614 546 622
rect 568 614 576 622
rect 588 614 596 622
rect 14 604 22 612
rect 224 604 232 612
rect 244 604 252 612
rect 266 604 274 612
rect 296 604 304 612
rect 326 604 334 612
rect 348 604 356 612
rect 368 604 376 612
rect 578 604 586 612
rect 4 594 12 602
rect 24 594 32 602
rect 54 594 62 602
rect 84 594 92 602
rect 114 594 122 602
rect 144 594 152 602
rect 174 594 182 602
rect 204 594 212 602
rect 234 594 242 602
rect 256 594 264 602
rect 276 594 284 602
rect 306 594 314 602
rect 336 594 344 602
rect 358 594 366 602
rect 388 594 396 602
rect 418 594 426 602
rect 448 594 456 602
rect 478 594 486 602
rect 508 594 516 602
rect 538 594 546 602
rect 568 594 576 602
rect 588 594 596 602
rect 14 584 22 592
rect 44 584 52 592
rect 74 584 82 592
rect 104 584 112 592
rect 134 584 142 592
rect 164 584 172 592
rect 194 584 202 592
rect 224 584 232 592
rect 244 584 252 592
rect 4 574 12 582
rect 24 574 32 582
rect 54 574 62 582
rect 84 574 92 582
rect 348 584 356 592
rect 368 584 376 592
rect 398 584 406 592
rect 428 584 436 592
rect 458 584 466 592
rect 488 584 496 592
rect 518 584 526 592
rect 548 584 556 592
rect 578 584 586 592
rect 508 574 516 582
rect 538 574 546 582
rect 568 574 576 582
rect 588 574 596 582
rect 14 564 22 572
rect 44 564 52 572
rect 74 564 82 572
rect 104 564 112 572
rect 134 564 142 572
rect 164 564 172 572
rect 194 564 202 572
rect 224 564 232 572
rect 244 564 252 572
rect 266 564 274 572
rect 296 564 304 572
rect 326 564 334 572
rect 348 564 356 572
rect 368 564 376 572
rect 398 564 406 572
rect 428 564 436 572
rect 458 564 466 572
rect 488 564 496 572
rect 518 564 526 572
rect 548 564 556 572
rect 578 564 586 572
rect 4 554 12 562
rect 24 554 32 562
rect 54 554 62 562
rect 84 554 92 562
rect 114 554 122 562
rect 144 554 152 562
rect 174 554 182 562
rect 204 554 212 562
rect 234 554 242 562
rect 256 554 264 562
rect 276 554 284 562
rect 306 554 314 562
rect 336 554 344 562
rect 358 554 366 562
rect 388 554 396 562
rect 418 554 426 562
rect 448 554 456 562
rect 478 554 486 562
rect 508 554 516 562
rect 538 554 546 562
rect 568 554 576 562
rect 588 554 596 562
rect 14 544 22 552
rect 44 544 52 552
rect 74 544 82 552
rect 104 544 112 552
rect 134 544 142 552
rect 164 544 172 552
rect 194 544 202 552
rect 224 544 232 552
rect 244 544 252 552
rect 266 544 274 552
rect 296 544 304 552
rect 326 544 334 552
rect 348 544 356 552
rect 368 544 376 552
rect 398 544 406 552
rect 428 544 436 552
rect 458 544 466 552
rect 488 544 496 552
rect 518 544 526 552
rect 548 544 556 552
rect 578 544 586 552
rect 4 534 12 542
rect 24 534 32 542
rect 54 534 62 542
rect 84 534 92 542
rect 114 534 122 542
rect 144 534 152 542
rect 174 534 182 542
rect 204 534 212 542
rect 234 534 242 542
rect 256 534 264 542
rect 276 534 284 542
rect 306 534 314 542
rect 336 534 344 542
rect 358 534 366 542
rect 388 534 396 542
rect 418 534 426 542
rect 448 534 456 542
rect 478 534 486 542
rect 508 534 516 542
rect 538 534 546 542
rect 568 534 576 542
rect 588 534 596 542
rect 14 524 22 532
rect 44 524 52 532
rect 74 524 82 532
rect 104 524 112 532
rect 134 524 142 532
rect 164 524 172 532
rect 194 524 202 532
rect 224 524 232 532
rect 244 524 252 532
rect 266 524 274 532
rect 296 524 304 532
rect 326 524 334 532
rect 348 524 356 532
rect 368 524 376 532
rect 398 524 406 532
rect 428 524 436 532
rect 458 524 466 532
rect 488 524 496 532
rect 518 524 526 532
rect 548 524 556 532
rect 578 524 586 532
rect 14 508 22 516
rect 34 508 42 516
rect 54 508 62 516
rect 74 508 82 516
rect 94 508 102 516
rect 114 508 122 516
rect 134 508 142 516
rect 154 508 162 516
rect 174 508 182 516
rect 194 508 202 516
rect 214 508 222 516
rect 234 508 242 516
rect 254 508 262 516
rect 274 508 282 516
rect 294 508 302 516
rect 308 508 316 516
rect 328 508 336 516
rect 348 508 356 516
rect 368 508 376 516
rect 388 508 396 516
rect 408 508 416 516
rect 428 508 436 516
rect 448 508 456 516
rect 468 508 476 516
rect 488 508 496 516
rect 508 508 516 516
rect 528 508 536 516
rect 548 508 556 516
rect 568 508 576 516
rect 38 446 56 454
rect 38 426 56 434
rect 38 406 56 414
rect 38 386 56 394
rect 38 366 56 374
rect 38 346 56 354
rect 38 326 56 334
rect 38 306 56 314
rect 38 286 56 294
rect 38 266 56 274
rect 38 246 56 254
rect 38 226 56 234
rect 38 206 56 214
rect 38 186 56 194
rect 38 166 56 174
rect 38 146 56 154
rect 38 126 56 134
rect 38 106 56 114
rect 38 86 56 94
rect 78 420 196 428
rect 78 390 106 420
rect 78 356 106 386
rect 291 444 309 452
rect 291 428 309 436
rect 291 412 309 420
rect 544 446 562 454
rect 404 420 522 428
rect 494 390 522 420
rect 78 348 236 356
rect 78 288 236 296
rect 78 226 106 288
rect 494 356 522 386
rect 364 348 522 356
rect 364 288 522 296
rect 291 252 309 260
rect 78 218 236 226
rect 78 158 236 166
rect 78 96 106 158
rect 494 226 522 288
rect 364 218 522 226
rect 364 158 522 166
rect 78 88 196 96
rect 38 66 56 74
rect 78 56 196 64
rect 38 46 66 54
rect 78 46 86 56
rect 98 46 106 56
rect 118 46 126 56
rect 138 46 146 56
rect 158 46 166 56
rect 178 46 186 56
rect 68 36 76 44
rect 88 36 96 44
rect 108 36 116 44
rect 128 36 136 44
rect 148 36 156 44
rect 168 36 176 44
rect 188 36 196 44
rect 291 124 309 132
rect 291 108 309 116
rect 291 92 309 100
rect 291 76 309 84
rect 291 60 309 68
rect 494 96 522 158
rect 404 88 522 96
rect 544 426 562 434
rect 544 406 562 414
rect 544 386 562 394
rect 544 366 562 374
rect 544 346 562 354
rect 544 326 562 334
rect 544 306 562 314
rect 544 286 562 294
rect 544 266 562 274
rect 544 246 562 254
rect 544 226 562 234
rect 544 206 562 214
rect 544 186 562 194
rect 544 166 562 174
rect 544 146 562 154
rect 544 126 562 134
rect 544 106 562 114
rect 544 86 562 94
rect 544 66 562 74
rect 404 56 522 64
rect 414 46 422 56
rect 434 46 442 56
rect 454 46 462 56
rect 474 46 482 56
rect 494 46 502 56
rect 514 46 522 56
rect 534 46 562 54
rect 404 36 412 44
rect 424 36 432 44
rect 444 36 452 44
rect 464 36 472 44
rect 484 36 492 44
rect 504 36 512 44
rect 524 36 532 44
<< metal2 >>
rect 0 1298 600 1340
rect 0 1290 56 1298
rect 64 1290 86 1298
rect 94 1290 116 1298
rect 124 1290 146 1298
rect 154 1290 176 1298
rect 184 1290 206 1298
rect 214 1290 236 1298
rect 244 1290 266 1298
rect 274 1290 296 1298
rect 304 1290 326 1298
rect 334 1290 356 1298
rect 364 1290 386 1298
rect 394 1290 416 1298
rect 424 1290 446 1298
rect 454 1290 476 1298
rect 484 1290 506 1298
rect 514 1290 536 1298
rect 544 1290 600 1298
rect 0 1288 600 1290
rect 0 1280 46 1288
rect 54 1280 66 1288
rect 74 1280 96 1288
rect 104 1280 126 1288
rect 134 1280 156 1288
rect 164 1280 186 1288
rect 194 1280 216 1288
rect 224 1280 246 1288
rect 254 1280 276 1288
rect 284 1280 306 1288
rect 314 1280 336 1288
rect 344 1280 366 1288
rect 374 1280 396 1288
rect 404 1280 426 1288
rect 434 1280 456 1288
rect 464 1280 486 1288
rect 494 1280 516 1288
rect 524 1280 546 1288
rect 554 1280 600 1288
rect 0 1278 600 1280
rect 0 1270 56 1278
rect 64 1270 86 1278
rect 94 1270 116 1278
rect 124 1270 146 1278
rect 154 1270 176 1278
rect 184 1270 206 1278
rect 214 1270 236 1278
rect 244 1270 266 1278
rect 274 1270 296 1278
rect 304 1270 326 1278
rect 334 1270 356 1278
rect 364 1270 386 1278
rect 394 1270 416 1278
rect 424 1270 446 1278
rect 454 1270 476 1278
rect 484 1270 506 1278
rect 514 1270 536 1278
rect 544 1270 600 1278
rect 0 1268 600 1270
rect 0 1260 46 1268
rect 54 1260 66 1268
rect 74 1260 96 1268
rect 104 1260 126 1268
rect 134 1260 156 1268
rect 164 1260 186 1268
rect 194 1260 216 1268
rect 224 1260 246 1268
rect 254 1260 276 1268
rect 284 1260 306 1268
rect 314 1260 336 1268
rect 344 1260 366 1268
rect 374 1260 396 1268
rect 404 1260 426 1268
rect 434 1260 456 1268
rect 464 1260 486 1268
rect 494 1260 516 1268
rect 524 1260 546 1268
rect 554 1260 600 1268
rect 0 1258 600 1260
rect 0 1250 56 1258
rect 64 1250 86 1258
rect 94 1250 116 1258
rect 124 1250 146 1258
rect 154 1250 176 1258
rect 184 1250 206 1258
rect 214 1250 236 1258
rect 244 1250 266 1258
rect 274 1250 296 1258
rect 304 1250 326 1258
rect 334 1250 356 1258
rect 364 1250 386 1258
rect 394 1250 416 1258
rect 424 1250 446 1258
rect 454 1250 476 1258
rect 484 1250 506 1258
rect 514 1250 536 1258
rect 544 1250 600 1258
rect 0 1248 600 1250
rect 0 1240 46 1248
rect 54 1240 66 1248
rect 74 1240 96 1248
rect 104 1240 126 1248
rect 134 1240 156 1248
rect 164 1240 186 1248
rect 194 1240 216 1248
rect 224 1240 246 1248
rect 254 1240 276 1248
rect 284 1240 306 1248
rect 314 1240 336 1248
rect 344 1240 366 1248
rect 374 1240 396 1248
rect 404 1240 426 1248
rect 434 1240 456 1248
rect 464 1240 486 1248
rect 494 1240 516 1248
rect 524 1240 546 1248
rect 554 1240 600 1248
rect 0 1238 600 1240
rect 0 1230 56 1238
rect 64 1230 86 1238
rect 94 1230 116 1238
rect 124 1230 146 1238
rect 154 1230 176 1238
rect 184 1230 206 1238
rect 214 1230 236 1238
rect 244 1230 266 1238
rect 274 1230 296 1238
rect 304 1230 326 1238
rect 334 1230 356 1238
rect 364 1230 386 1238
rect 394 1230 416 1238
rect 424 1230 446 1238
rect 454 1230 476 1238
rect 484 1230 506 1238
rect 514 1230 536 1238
rect 544 1230 600 1238
rect 0 1228 600 1230
rect 0 1220 46 1228
rect 54 1220 66 1228
rect 74 1220 96 1228
rect 104 1220 126 1228
rect 134 1220 156 1228
rect 164 1220 186 1228
rect 194 1220 216 1228
rect 224 1220 246 1228
rect 254 1220 276 1228
rect 284 1220 306 1228
rect 314 1220 336 1228
rect 344 1220 366 1228
rect 374 1220 396 1228
rect 404 1220 426 1228
rect 434 1220 456 1228
rect 464 1220 486 1228
rect 494 1220 516 1228
rect 524 1220 546 1228
rect 554 1220 600 1228
rect 0 1218 600 1220
rect 0 1210 56 1218
rect 64 1210 86 1218
rect 94 1210 116 1218
rect 124 1210 146 1218
rect 154 1210 176 1218
rect 184 1210 206 1218
rect 214 1210 236 1218
rect 244 1210 266 1218
rect 274 1210 296 1218
rect 304 1210 326 1218
rect 334 1210 356 1218
rect 364 1210 386 1218
rect 394 1210 416 1218
rect 424 1210 446 1218
rect 454 1210 476 1218
rect 484 1210 506 1218
rect 514 1210 536 1218
rect 544 1210 600 1218
rect 0 1208 600 1210
rect 0 1200 46 1208
rect 54 1200 66 1208
rect 74 1200 96 1208
rect 104 1200 126 1208
rect 134 1200 156 1208
rect 164 1200 186 1208
rect 194 1200 216 1208
rect 224 1200 246 1208
rect 254 1200 276 1208
rect 284 1200 306 1208
rect 314 1200 336 1208
rect 344 1200 366 1208
rect 374 1200 396 1208
rect 404 1200 426 1208
rect 434 1200 456 1208
rect 464 1200 486 1208
rect 494 1200 516 1208
rect 524 1200 546 1208
rect 554 1200 600 1208
rect 0 1198 600 1200
rect 0 1190 56 1198
rect 64 1190 86 1198
rect 94 1190 116 1198
rect 124 1190 146 1198
rect 154 1190 176 1198
rect 184 1190 206 1198
rect 214 1190 236 1198
rect 244 1190 266 1198
rect 274 1190 296 1198
rect 304 1190 326 1198
rect 334 1190 356 1198
rect 364 1190 386 1198
rect 394 1190 416 1198
rect 424 1190 446 1198
rect 454 1190 476 1198
rect 484 1190 506 1198
rect 514 1190 536 1198
rect 544 1190 600 1198
rect 0 1188 100 1190
rect 0 1180 46 1188
rect 54 1180 66 1188
rect 74 1180 100 1188
rect 500 1188 600 1190
rect 500 1180 516 1188
rect 524 1180 546 1188
rect 554 1180 600 1188
rect 0 1178 600 1180
rect 0 1170 56 1178
rect 64 1170 86 1178
rect 94 1170 116 1178
rect 124 1170 146 1178
rect 154 1170 176 1178
rect 184 1170 206 1178
rect 214 1170 236 1178
rect 244 1170 266 1178
rect 274 1170 296 1178
rect 304 1170 326 1178
rect 334 1170 356 1178
rect 364 1170 386 1178
rect 394 1170 416 1178
rect 424 1170 446 1178
rect 454 1170 476 1178
rect 484 1170 506 1178
rect 514 1170 536 1178
rect 544 1170 600 1178
rect 0 1168 600 1170
rect 0 1160 46 1168
rect 54 1160 66 1168
rect 74 1160 96 1168
rect 104 1160 126 1168
rect 134 1160 156 1168
rect 164 1160 186 1168
rect 194 1160 216 1168
rect 224 1160 246 1168
rect 254 1160 276 1168
rect 284 1160 306 1168
rect 314 1160 336 1168
rect 344 1160 366 1168
rect 374 1160 396 1168
rect 404 1160 426 1168
rect 434 1160 456 1168
rect 464 1160 486 1168
rect 494 1160 516 1168
rect 524 1160 546 1168
rect 554 1160 600 1168
rect 0 1158 600 1160
rect 0 1150 56 1158
rect 64 1150 86 1158
rect 94 1150 116 1158
rect 124 1150 146 1158
rect 154 1150 176 1158
rect 184 1150 206 1158
rect 214 1150 236 1158
rect 244 1150 266 1158
rect 274 1150 296 1158
rect 304 1150 326 1158
rect 334 1150 356 1158
rect 364 1150 386 1158
rect 394 1150 416 1158
rect 424 1150 446 1158
rect 454 1150 476 1158
rect 484 1150 506 1158
rect 514 1150 536 1158
rect 544 1150 600 1158
rect 0 1148 600 1150
rect 0 1140 46 1148
rect 54 1140 66 1148
rect 74 1140 96 1148
rect 104 1140 126 1148
rect 134 1140 156 1148
rect 164 1140 186 1148
rect 194 1140 216 1148
rect 224 1140 246 1148
rect 254 1140 276 1148
rect 284 1140 306 1148
rect 314 1140 336 1148
rect 344 1140 366 1148
rect 374 1140 396 1148
rect 404 1140 426 1148
rect 434 1140 456 1148
rect 464 1140 486 1148
rect 494 1140 516 1148
rect 524 1140 546 1148
rect 554 1140 600 1148
rect 0 1138 600 1140
rect 0 1130 56 1138
rect 64 1130 86 1138
rect 94 1130 116 1138
rect 124 1130 146 1138
rect 154 1130 176 1138
rect 184 1130 206 1138
rect 214 1130 236 1138
rect 244 1130 266 1138
rect 274 1130 296 1138
rect 304 1130 326 1138
rect 334 1130 356 1138
rect 364 1130 386 1138
rect 394 1130 416 1138
rect 424 1130 446 1138
rect 454 1130 476 1138
rect 484 1130 506 1138
rect 514 1130 536 1138
rect 544 1130 600 1138
rect 0 1128 600 1130
rect 0 1120 46 1128
rect 54 1120 66 1128
rect 74 1120 96 1128
rect 104 1120 126 1128
rect 134 1120 156 1128
rect 164 1120 186 1128
rect 194 1120 216 1128
rect 224 1120 246 1128
rect 254 1120 276 1128
rect 284 1120 306 1128
rect 314 1120 336 1128
rect 344 1120 366 1128
rect 374 1120 396 1128
rect 404 1120 426 1128
rect 434 1120 456 1128
rect 464 1120 486 1128
rect 494 1120 516 1128
rect 0 1118 516 1120
rect 0 1110 56 1118
rect 64 1110 76 1118
rect 84 1110 516 1118
rect 0 1108 516 1110
rect 0 1100 46 1108
rect 54 1100 66 1108
rect 74 1100 96 1108
rect 104 1100 126 1108
rect 134 1100 156 1108
rect 164 1100 186 1108
rect 194 1100 216 1108
rect 224 1100 246 1108
rect 254 1100 276 1108
rect 284 1100 306 1108
rect 314 1100 336 1108
rect 344 1100 366 1108
rect 374 1100 396 1108
rect 404 1100 426 1108
rect 434 1100 456 1108
rect 464 1100 486 1108
rect 494 1100 516 1108
rect 524 1120 546 1128
rect 554 1120 600 1128
rect 524 1118 600 1120
rect 524 1110 536 1118
rect 544 1110 600 1118
rect 524 1108 600 1110
rect 524 1100 546 1108
rect 554 1100 600 1108
rect 0 1098 600 1100
rect 0 1090 56 1098
rect 64 1090 86 1098
rect 94 1090 116 1098
rect 124 1090 146 1098
rect 154 1090 176 1098
rect 184 1090 206 1098
rect 214 1090 236 1098
rect 244 1090 266 1098
rect 274 1090 296 1098
rect 304 1090 326 1098
rect 334 1090 356 1098
rect 364 1090 386 1098
rect 394 1090 416 1098
rect 424 1090 446 1098
rect 454 1090 476 1098
rect 484 1090 506 1098
rect 514 1090 536 1098
rect 544 1090 600 1098
rect 0 1088 600 1090
rect 0 1080 46 1088
rect 54 1080 66 1088
rect 74 1080 96 1088
rect 104 1080 126 1088
rect 134 1080 156 1088
rect 164 1080 186 1088
rect 194 1080 216 1088
rect 224 1080 246 1088
rect 254 1080 276 1088
rect 284 1080 306 1088
rect 314 1080 336 1088
rect 344 1080 366 1088
rect 374 1080 396 1088
rect 404 1080 426 1088
rect 434 1080 456 1088
rect 464 1080 486 1088
rect 494 1080 516 1088
rect 524 1080 546 1088
rect 554 1080 600 1088
rect 0 1078 600 1080
rect 0 1070 56 1078
rect 64 1070 86 1078
rect 94 1070 116 1078
rect 124 1070 146 1078
rect 154 1070 176 1078
rect 184 1070 206 1078
rect 214 1070 236 1078
rect 244 1070 266 1078
rect 274 1070 296 1078
rect 304 1070 326 1078
rect 334 1070 356 1078
rect 364 1070 386 1078
rect 394 1070 416 1078
rect 424 1070 446 1078
rect 454 1070 476 1078
rect 484 1070 506 1078
rect 514 1070 536 1078
rect 544 1070 600 1078
rect 0 1068 600 1070
rect 0 1060 46 1068
rect 54 1060 66 1068
rect 74 1060 96 1068
rect 104 1060 126 1068
rect 134 1060 156 1068
rect 164 1060 186 1068
rect 194 1060 216 1068
rect 224 1060 246 1068
rect 254 1060 276 1068
rect 284 1060 306 1068
rect 314 1060 336 1068
rect 344 1060 366 1068
rect 374 1060 396 1068
rect 404 1060 426 1068
rect 434 1060 456 1068
rect 464 1060 486 1068
rect 494 1060 516 1068
rect 524 1060 546 1068
rect 554 1060 600 1068
rect 0 1058 600 1060
rect 0 1050 56 1058
rect 64 1050 86 1058
rect 94 1050 116 1058
rect 124 1050 146 1058
rect 154 1050 176 1058
rect 184 1050 206 1058
rect 214 1050 236 1058
rect 244 1050 266 1058
rect 274 1050 296 1058
rect 304 1050 326 1058
rect 334 1050 356 1058
rect 364 1050 386 1058
rect 394 1050 416 1058
rect 424 1050 446 1058
rect 454 1050 476 1058
rect 484 1050 506 1058
rect 514 1050 536 1058
rect 544 1050 600 1058
rect 0 1048 600 1050
rect 0 1040 46 1048
rect 54 1040 66 1048
rect 74 1040 96 1048
rect 104 1040 126 1048
rect 134 1040 156 1048
rect 164 1040 186 1048
rect 194 1040 216 1048
rect 224 1040 246 1048
rect 254 1040 276 1048
rect 284 1040 306 1048
rect 314 1040 336 1048
rect 344 1040 366 1048
rect 374 1040 396 1048
rect 404 1040 426 1048
rect 434 1040 456 1048
rect 464 1040 486 1048
rect 494 1040 516 1048
rect 0 1038 100 1040
rect 0 1030 56 1038
rect 64 1030 86 1038
rect 94 1030 100 1038
rect 500 1030 516 1040
rect 0 1028 516 1030
rect 0 1020 46 1028
rect 54 1020 66 1028
rect 74 1020 96 1028
rect 104 1020 126 1028
rect 134 1020 156 1028
rect 164 1020 186 1028
rect 194 1020 216 1028
rect 224 1020 246 1028
rect 254 1020 276 1028
rect 284 1020 306 1028
rect 314 1020 336 1028
rect 344 1020 366 1028
rect 374 1020 396 1028
rect 404 1020 426 1028
rect 434 1020 456 1028
rect 464 1020 486 1028
rect 494 1020 516 1028
rect 524 1040 546 1048
rect 554 1040 600 1048
rect 524 1038 600 1040
rect 524 1030 536 1038
rect 544 1030 600 1038
rect 524 1028 600 1030
rect 524 1020 546 1028
rect 554 1020 600 1028
rect 0 1018 600 1020
rect 0 1010 56 1018
rect 64 1010 86 1018
rect 94 1010 116 1018
rect 124 1010 146 1018
rect 154 1010 176 1018
rect 184 1010 206 1018
rect 214 1010 236 1018
rect 244 1010 266 1018
rect 274 1010 296 1018
rect 304 1010 326 1018
rect 334 1010 356 1018
rect 364 1010 386 1018
rect 394 1010 416 1018
rect 424 1010 446 1018
rect 454 1010 476 1018
rect 484 1010 506 1018
rect 514 1010 536 1018
rect 544 1010 600 1018
rect 0 1008 600 1010
rect 0 1000 46 1008
rect 54 1000 66 1008
rect 74 1000 96 1008
rect 104 1000 126 1008
rect 134 1000 156 1008
rect 164 1000 186 1008
rect 194 1000 216 1008
rect 224 1000 246 1008
rect 254 1000 276 1008
rect 284 1000 306 1008
rect 314 1000 336 1008
rect 344 1000 366 1008
rect 374 1000 396 1008
rect 404 1000 426 1008
rect 434 1000 456 1008
rect 464 1000 486 1008
rect 494 1000 516 1008
rect 524 1000 546 1008
rect 554 1000 600 1008
rect 0 998 600 1000
rect 0 990 56 998
rect 64 990 86 998
rect 94 990 116 998
rect 124 990 146 998
rect 154 990 176 998
rect 184 990 206 998
rect 214 990 236 998
rect 244 990 266 998
rect 274 990 296 998
rect 304 990 326 998
rect 334 990 356 998
rect 364 990 386 998
rect 394 990 416 998
rect 424 990 446 998
rect 454 990 476 998
rect 484 990 506 998
rect 514 990 536 998
rect 544 990 600 998
rect 0 988 600 990
rect 0 980 46 988
rect 54 980 66 988
rect 74 980 96 988
rect 104 980 126 988
rect 134 980 156 988
rect 164 980 186 988
rect 194 980 216 988
rect 224 980 246 988
rect 254 980 276 988
rect 284 980 306 988
rect 314 980 336 988
rect 344 980 366 988
rect 374 980 396 988
rect 404 980 426 988
rect 434 980 456 988
rect 464 980 486 988
rect 494 980 516 988
rect 524 980 546 988
rect 554 980 600 988
rect 0 978 600 980
rect 0 970 56 978
rect 64 970 86 978
rect 94 970 116 978
rect 124 970 146 978
rect 154 970 176 978
rect 184 970 206 978
rect 214 970 236 978
rect 244 970 266 978
rect 274 970 296 978
rect 304 970 326 978
rect 334 970 356 978
rect 364 970 386 978
rect 394 970 416 978
rect 424 970 446 978
rect 454 970 476 978
rect 484 970 506 978
rect 514 970 536 978
rect 544 970 600 978
rect 0 968 600 970
rect 0 960 46 968
rect 54 960 546 968
rect 554 960 600 968
rect 0 958 600 960
rect 0 950 56 958
rect 64 950 86 958
rect 94 950 116 958
rect 124 950 146 958
rect 154 950 176 958
rect 184 950 206 958
rect 214 950 236 958
rect 244 950 266 958
rect 274 950 296 958
rect 304 950 326 958
rect 334 950 356 958
rect 364 950 386 958
rect 394 950 416 958
rect 424 950 446 958
rect 454 950 476 958
rect 484 950 506 958
rect 514 950 536 958
rect 544 950 600 958
rect 0 948 600 950
rect 0 940 46 948
rect 54 940 66 948
rect 74 940 96 948
rect 104 940 126 948
rect 134 940 156 948
rect 164 940 186 948
rect 194 940 216 948
rect 224 940 246 948
rect 254 940 276 948
rect 284 940 306 948
rect 314 940 336 948
rect 344 940 366 948
rect 374 940 396 948
rect 404 940 426 948
rect 434 940 456 948
rect 464 940 486 948
rect 494 940 516 948
rect 524 940 546 948
rect 554 940 600 948
rect 0 938 600 940
rect 0 930 56 938
rect 64 930 86 938
rect 94 930 116 938
rect 124 930 146 938
rect 154 930 176 938
rect 184 930 206 938
rect 214 930 236 938
rect 244 930 266 938
rect 274 930 296 938
rect 304 930 326 938
rect 334 930 356 938
rect 364 930 386 938
rect 394 930 416 938
rect 424 930 446 938
rect 454 930 476 938
rect 484 930 506 938
rect 514 930 536 938
rect 544 930 600 938
rect 0 928 600 930
rect 0 920 46 928
rect 54 920 66 928
rect 74 920 96 928
rect 104 920 126 928
rect 134 920 156 928
rect 164 920 186 928
rect 194 920 216 928
rect 224 920 246 928
rect 254 920 276 928
rect 284 920 306 928
rect 314 920 336 928
rect 344 920 366 928
rect 374 920 396 928
rect 404 920 426 928
rect 434 920 456 928
rect 464 920 486 928
rect 494 920 516 928
rect 524 920 546 928
rect 554 920 600 928
rect 0 918 600 920
rect 0 910 56 918
rect 64 910 86 918
rect 94 910 116 918
rect 124 910 146 918
rect 154 910 176 918
rect 184 910 206 918
rect 214 910 236 918
rect 244 910 266 918
rect 274 910 296 918
rect 304 910 326 918
rect 334 910 356 918
rect 364 910 386 918
rect 394 910 416 918
rect 424 910 446 918
rect 454 910 476 918
rect 484 910 506 918
rect 514 910 536 918
rect 544 910 600 918
rect 0 908 600 910
rect 0 900 46 908
rect 54 900 66 908
rect 74 900 96 908
rect 104 900 126 908
rect 134 900 156 908
rect 164 900 186 908
rect 194 900 216 908
rect 224 900 246 908
rect 254 900 276 908
rect 284 900 306 908
rect 314 900 336 908
rect 344 900 366 908
rect 374 900 396 908
rect 404 900 426 908
rect 434 900 456 908
rect 464 900 486 908
rect 494 900 516 908
rect 524 900 546 908
rect 554 900 600 908
rect 0 898 600 900
rect 0 890 56 898
rect 64 890 86 898
rect 94 890 116 898
rect 124 890 146 898
rect 154 890 176 898
rect 184 890 206 898
rect 214 890 236 898
rect 244 890 266 898
rect 274 890 296 898
rect 304 890 326 898
rect 334 890 356 898
rect 364 890 386 898
rect 394 890 416 898
rect 424 890 446 898
rect 454 890 476 898
rect 484 890 506 898
rect 514 890 536 898
rect 544 890 600 898
rect 0 888 600 890
rect 0 880 46 888
rect 54 880 66 888
rect 74 880 96 888
rect 104 880 126 888
rect 134 880 156 888
rect 164 880 186 888
rect 194 880 216 888
rect 224 880 246 888
rect 254 880 276 888
rect 284 880 306 888
rect 314 880 336 888
rect 344 880 366 888
rect 374 880 396 888
rect 404 880 426 888
rect 434 880 456 888
rect 464 880 486 888
rect 494 880 516 888
rect 524 880 546 888
rect 554 880 600 888
rect 0 836 600 848
rect 0 828 14 836
rect 22 828 44 836
rect 52 828 74 836
rect 82 828 104 836
rect 112 828 134 836
rect 142 828 164 836
rect 172 828 184 836
rect 192 828 286 836
rect 294 828 306 836
rect 314 828 408 836
rect 416 828 428 836
rect 436 828 458 836
rect 466 828 488 836
rect 496 828 518 836
rect 526 828 548 836
rect 556 828 578 836
rect 586 828 600 836
rect 0 826 600 828
rect 0 818 4 826
rect 12 818 24 826
rect 32 818 54 826
rect 62 818 84 826
rect 92 818 114 826
rect 122 818 144 826
rect 152 818 174 826
rect 182 818 296 826
rect 304 818 418 826
rect 426 818 448 826
rect 456 818 478 826
rect 486 818 508 826
rect 516 818 538 826
rect 546 818 568 826
rect 576 818 588 826
rect 596 818 600 826
rect 0 816 600 818
rect 0 808 14 816
rect 22 808 44 816
rect 52 808 74 816
rect 82 808 104 816
rect 112 808 134 816
rect 142 808 164 816
rect 172 808 184 816
rect 192 808 286 816
rect 294 808 306 816
rect 314 808 408 816
rect 416 808 428 816
rect 436 808 458 816
rect 466 808 488 816
rect 496 808 518 816
rect 526 808 548 816
rect 556 808 578 816
rect 586 808 600 816
rect 0 806 600 808
rect 0 798 4 806
rect 12 798 24 806
rect 32 798 54 806
rect 62 798 84 806
rect 92 798 114 806
rect 122 798 144 806
rect 152 798 174 806
rect 182 798 296 806
rect 304 798 418 806
rect 426 798 448 806
rect 456 798 478 806
rect 486 798 508 806
rect 516 798 538 806
rect 546 798 568 806
rect 576 798 588 806
rect 596 798 600 806
rect 0 796 600 798
rect 0 788 14 796
rect 22 788 44 796
rect 52 788 74 796
rect 82 788 104 796
rect 112 788 134 796
rect 142 788 164 796
rect 172 788 184 796
rect 192 788 286 796
rect 294 788 306 796
rect 314 788 408 796
rect 416 788 428 796
rect 436 788 458 796
rect 466 788 488 796
rect 496 788 518 796
rect 526 788 548 796
rect 556 788 578 796
rect 586 788 600 796
rect 0 786 600 788
rect 0 778 4 786
rect 12 778 24 786
rect 32 778 54 786
rect 62 778 84 786
rect 92 778 114 786
rect 122 778 144 786
rect 152 778 174 786
rect 182 778 296 786
rect 304 778 418 786
rect 426 778 448 786
rect 456 778 478 786
rect 486 778 508 786
rect 516 778 538 786
rect 546 778 568 786
rect 576 778 588 786
rect 596 778 600 786
rect 0 776 100 778
rect 0 768 14 776
rect 22 768 44 776
rect 52 768 74 776
rect 82 768 100 776
rect 500 776 600 778
rect 500 768 518 776
rect 526 768 548 776
rect 556 768 578 776
rect 586 768 600 776
rect 0 766 600 768
rect 0 758 4 766
rect 12 758 24 766
rect 32 758 54 766
rect 62 758 84 766
rect 92 758 114 766
rect 122 758 144 766
rect 152 758 174 766
rect 182 758 286 766
rect 294 758 306 766
rect 314 758 418 766
rect 426 758 448 766
rect 456 758 478 766
rect 486 758 508 766
rect 516 758 538 766
rect 546 758 568 766
rect 576 758 588 766
rect 596 758 600 766
rect 0 756 600 758
rect 0 748 14 756
rect 22 748 44 756
rect 52 748 74 756
rect 82 748 104 756
rect 112 748 134 756
rect 142 748 164 756
rect 172 748 184 756
rect 192 748 296 756
rect 304 748 408 756
rect 416 748 428 756
rect 436 748 458 756
rect 466 748 488 756
rect 496 748 518 756
rect 526 748 548 756
rect 556 748 578 756
rect 586 748 600 756
rect 0 746 600 748
rect 0 738 4 746
rect 12 738 24 746
rect 32 738 54 746
rect 62 738 84 746
rect 92 738 114 746
rect 122 738 144 746
rect 152 738 174 746
rect 182 738 286 746
rect 294 738 306 746
rect 314 738 418 746
rect 426 738 448 746
rect 456 738 478 746
rect 486 738 508 746
rect 516 738 538 746
rect 546 738 568 746
rect 576 738 588 746
rect 596 738 600 746
rect 0 736 600 738
rect 0 728 14 736
rect 22 728 296 736
rect 304 728 578 736
rect 586 728 600 736
rect 0 726 600 728
rect 0 718 4 726
rect 12 718 24 726
rect 32 718 54 726
rect 62 718 84 726
rect 92 718 114 726
rect 122 718 144 726
rect 152 718 174 726
rect 182 718 286 726
rect 294 718 306 726
rect 314 718 418 726
rect 426 718 448 726
rect 456 718 478 726
rect 486 718 508 726
rect 516 718 538 726
rect 546 718 568 726
rect 576 718 588 726
rect 596 718 600 726
rect 0 716 600 718
rect 0 708 14 716
rect 22 708 44 716
rect 52 708 74 716
rect 82 708 104 716
rect 112 708 134 716
rect 142 708 164 716
rect 172 708 184 716
rect 192 708 296 716
rect 0 706 296 708
rect 304 708 408 716
rect 416 708 428 716
rect 436 708 458 716
rect 466 708 488 716
rect 496 708 518 716
rect 526 708 548 716
rect 556 708 578 716
rect 586 708 600 716
rect 304 706 600 708
rect 0 698 4 706
rect 12 698 24 706
rect 32 698 54 706
rect 62 698 84 706
rect 92 698 114 706
rect 122 698 144 706
rect 152 698 174 706
rect 182 698 286 706
rect 314 698 418 706
rect 426 698 448 706
rect 456 698 478 706
rect 486 698 508 706
rect 516 698 538 706
rect 546 698 568 706
rect 576 698 588 706
rect 596 698 600 706
rect 0 696 600 698
rect 0 688 14 696
rect 22 688 44 696
rect 52 688 74 696
rect 82 688 104 696
rect 112 688 134 696
rect 142 688 164 696
rect 172 688 184 696
rect 192 688 408 696
rect 416 688 428 696
rect 436 688 458 696
rect 466 688 488 696
rect 496 688 518 696
rect 526 688 548 696
rect 556 688 578 696
rect 586 688 600 696
rect 0 644 14 652
rect 22 644 44 652
rect 52 644 74 652
rect 82 644 104 652
rect 112 644 134 652
rect 142 644 164 652
rect 172 644 194 652
rect 202 644 224 652
rect 232 644 244 652
rect 252 644 266 652
rect 274 644 296 652
rect 304 644 326 652
rect 334 644 348 652
rect 356 644 368 652
rect 376 644 398 652
rect 406 644 428 652
rect 436 644 458 652
rect 466 644 488 652
rect 496 644 518 652
rect 526 644 548 652
rect 556 644 578 652
rect 586 644 600 652
rect 0 642 600 644
rect 0 634 4 642
rect 12 634 24 642
rect 32 634 54 642
rect 62 634 84 642
rect 92 634 114 642
rect 122 634 144 642
rect 152 634 174 642
rect 182 634 204 642
rect 212 634 234 642
rect 242 634 256 642
rect 264 634 276 642
rect 284 634 306 642
rect 314 634 336 642
rect 344 634 358 642
rect 366 634 388 642
rect 396 634 418 642
rect 426 634 448 642
rect 456 634 478 642
rect 486 634 508 642
rect 516 634 538 642
rect 546 634 568 642
rect 576 634 588 642
rect 596 634 600 642
rect 0 632 600 634
rect 0 624 14 632
rect 22 624 44 632
rect 52 624 74 632
rect 82 624 104 632
rect 112 624 134 632
rect 142 624 164 632
rect 172 624 194 632
rect 202 624 224 632
rect 232 624 244 632
rect 252 624 266 632
rect 274 624 296 632
rect 304 624 326 632
rect 334 624 348 632
rect 356 624 368 632
rect 376 624 398 632
rect 406 624 428 632
rect 436 624 458 632
rect 466 624 488 632
rect 496 624 518 632
rect 526 624 548 632
rect 556 624 578 632
rect 586 624 600 632
rect 0 622 600 624
rect 0 614 4 622
rect 12 614 24 622
rect 32 614 54 622
rect 62 614 84 622
rect 92 614 114 622
rect 122 614 144 622
rect 152 614 174 622
rect 182 614 204 622
rect 212 614 234 622
rect 242 614 256 622
rect 264 614 276 622
rect 284 614 306 622
rect 314 614 336 622
rect 344 614 358 622
rect 366 614 388 622
rect 396 614 418 622
rect 426 614 448 622
rect 456 614 478 622
rect 486 614 508 622
rect 516 614 538 622
rect 546 614 568 622
rect 576 614 588 622
rect 596 614 600 622
rect 0 612 600 614
rect 0 604 14 612
rect 22 604 224 612
rect 232 604 244 612
rect 252 604 266 612
rect 274 604 296 612
rect 304 604 326 612
rect 334 604 348 612
rect 356 604 368 612
rect 376 604 578 612
rect 586 604 600 612
rect 0 602 600 604
rect 0 594 4 602
rect 12 594 24 602
rect 32 594 54 602
rect 62 594 84 602
rect 92 594 114 602
rect 122 594 144 602
rect 152 594 174 602
rect 182 594 204 602
rect 212 594 234 602
rect 242 594 256 602
rect 264 594 276 602
rect 284 594 306 602
rect 314 594 336 602
rect 344 594 358 602
rect 366 594 388 602
rect 396 594 418 602
rect 426 594 448 602
rect 456 594 478 602
rect 486 594 508 602
rect 516 594 538 602
rect 546 594 568 602
rect 576 594 588 602
rect 596 594 600 602
rect 0 592 600 594
rect 0 584 14 592
rect 22 584 44 592
rect 52 584 74 592
rect 82 584 104 592
rect 112 584 134 592
rect 142 584 164 592
rect 172 584 194 592
rect 202 584 224 592
rect 232 584 244 592
rect 252 584 348 592
rect 356 584 368 592
rect 376 584 398 592
rect 406 584 428 592
rect 436 584 458 592
rect 466 584 488 592
rect 496 584 518 592
rect 526 584 548 592
rect 556 584 578 592
rect 586 584 600 592
rect 0 582 600 584
rect 0 574 4 582
rect 12 574 24 582
rect 32 574 54 582
rect 62 574 84 582
rect 92 574 100 582
rect 0 572 100 574
rect 500 574 508 582
rect 516 574 538 582
rect 546 574 568 582
rect 576 574 588 582
rect 596 574 600 582
rect 500 572 600 574
rect 0 564 14 572
rect 22 564 44 572
rect 52 564 74 572
rect 82 564 104 572
rect 112 564 134 572
rect 142 564 164 572
rect 172 564 194 572
rect 202 564 224 572
rect 232 564 244 572
rect 252 564 266 572
rect 274 564 296 572
rect 304 564 326 572
rect 334 564 348 572
rect 356 564 368 572
rect 376 564 398 572
rect 406 564 428 572
rect 436 564 458 572
rect 466 564 488 572
rect 496 564 518 572
rect 526 564 548 572
rect 556 564 578 572
rect 586 564 600 572
rect 0 562 600 564
rect 0 554 4 562
rect 12 554 24 562
rect 32 554 54 562
rect 62 554 84 562
rect 92 554 114 562
rect 122 554 144 562
rect 152 554 174 562
rect 182 554 204 562
rect 212 554 234 562
rect 242 554 256 562
rect 264 554 276 562
rect 284 554 306 562
rect 314 554 336 562
rect 344 554 358 562
rect 366 554 388 562
rect 396 554 418 562
rect 426 554 448 562
rect 456 554 478 562
rect 486 554 508 562
rect 516 554 538 562
rect 546 554 568 562
rect 576 554 588 562
rect 596 554 600 562
rect 0 552 600 554
rect 0 544 14 552
rect 22 544 44 552
rect 52 544 74 552
rect 82 544 104 552
rect 112 544 134 552
rect 142 544 164 552
rect 172 544 194 552
rect 202 544 224 552
rect 232 544 244 552
rect 252 544 266 552
rect 274 544 296 552
rect 304 544 326 552
rect 334 544 348 552
rect 356 544 368 552
rect 376 544 398 552
rect 406 544 428 552
rect 436 544 458 552
rect 466 544 488 552
rect 496 544 518 552
rect 526 544 548 552
rect 556 544 578 552
rect 586 544 600 552
rect 0 542 600 544
rect 0 534 4 542
rect 12 534 24 542
rect 32 534 54 542
rect 62 534 84 542
rect 92 534 114 542
rect 122 534 144 542
rect 152 534 174 542
rect 182 534 204 542
rect 212 534 234 542
rect 242 534 256 542
rect 264 534 276 542
rect 284 534 306 542
rect 314 534 336 542
rect 344 534 358 542
rect 366 534 388 542
rect 396 534 418 542
rect 426 534 448 542
rect 456 534 478 542
rect 486 534 508 542
rect 516 534 538 542
rect 546 534 568 542
rect 576 534 588 542
rect 596 534 600 542
rect 0 532 600 534
rect 0 524 14 532
rect 22 524 44 532
rect 52 524 74 532
rect 82 524 104 532
rect 112 524 134 532
rect 142 524 164 532
rect 172 524 194 532
rect 202 524 224 532
rect 232 524 244 532
rect 252 524 266 532
rect 274 524 296 532
rect 304 524 326 532
rect 334 524 348 532
rect 356 524 368 532
rect 376 524 398 532
rect 406 524 428 532
rect 436 524 458 532
rect 466 524 488 532
rect 496 524 518 532
rect 526 524 548 532
rect 556 524 578 532
rect 586 524 600 532
rect 0 516 600 524
rect 0 508 14 516
rect 22 508 34 516
rect 42 508 54 516
rect 62 508 74 516
rect 82 508 94 516
rect 102 508 114 516
rect 122 508 134 516
rect 142 508 154 516
rect 162 508 174 516
rect 182 508 194 516
rect 202 508 214 516
rect 222 508 234 516
rect 242 508 254 516
rect 262 508 274 516
rect 282 508 294 516
rect 302 508 308 516
rect 316 508 328 516
rect 336 508 348 516
rect 356 508 368 516
rect 376 508 388 516
rect 396 508 408 516
rect 416 508 428 516
rect 436 508 448 516
rect 456 508 468 516
rect 476 508 488 516
rect 496 508 508 516
rect 516 508 528 516
rect 536 508 548 516
rect 556 508 568 516
rect 576 508 600 516
rect 0 492 600 508
rect 0 454 600 458
rect 0 446 38 454
rect 56 452 544 454
rect 56 446 291 452
rect 0 444 291 446
rect 309 446 544 452
rect 562 446 600 454
rect 309 444 600 446
rect 0 436 600 444
rect 0 434 291 436
rect 0 426 38 434
rect 56 428 291 434
rect 309 434 600 436
rect 309 428 544 434
rect 56 426 78 428
rect 0 414 78 426
rect 196 420 404 428
rect 522 426 544 428
rect 562 426 600 434
rect 0 406 38 414
rect 56 406 78 414
rect 0 394 78 406
rect 0 386 38 394
rect 56 390 78 394
rect 106 412 291 420
rect 309 412 494 420
rect 106 390 494 412
rect 522 414 600 426
rect 522 406 544 414
rect 562 406 600 414
rect 522 394 600 406
rect 522 390 544 394
rect 56 386 544 390
rect 562 386 600 394
rect 0 374 78 386
rect 0 366 38 374
rect 56 366 78 374
rect 0 354 78 366
rect 106 356 494 386
rect 522 374 600 386
rect 522 366 544 374
rect 562 366 600 374
rect 0 346 38 354
rect 56 348 78 354
rect 236 348 364 356
rect 522 354 600 366
rect 522 348 544 354
rect 56 346 544 348
rect 562 346 600 354
rect 0 334 600 346
rect 0 326 38 334
rect 56 326 544 334
rect 562 326 600 334
rect 0 314 600 326
rect 0 306 38 314
rect 56 308 544 314
rect 56 306 100 308
rect 0 298 100 306
rect 500 306 544 308
rect 562 306 600 314
rect 500 298 600 306
rect 0 296 600 298
rect 0 294 78 296
rect 0 286 38 294
rect 56 286 78 294
rect 236 288 364 296
rect 522 294 600 296
rect 0 274 78 286
rect 0 266 38 274
rect 56 266 78 274
rect 0 254 78 266
rect 0 246 38 254
rect 56 246 78 254
rect 0 234 78 246
rect 0 226 38 234
rect 56 226 78 234
rect 106 260 494 288
rect 106 252 291 260
rect 309 252 494 260
rect 106 226 494 252
rect 522 286 544 294
rect 562 286 600 294
rect 522 274 600 286
rect 522 266 544 274
rect 562 266 600 274
rect 522 254 600 266
rect 522 246 544 254
rect 562 246 600 254
rect 522 234 600 246
rect 522 226 544 234
rect 562 226 600 234
rect 0 218 78 226
rect 236 218 364 226
rect 522 218 600 226
rect 0 214 600 218
rect 0 206 38 214
rect 56 206 544 214
rect 562 206 600 214
rect 0 194 600 206
rect 0 186 38 194
rect 56 186 544 194
rect 562 186 600 194
rect 0 174 600 186
rect 0 166 38 174
rect 56 166 544 174
rect 562 166 600 174
rect 0 154 78 166
rect 236 158 364 166
rect 0 146 38 154
rect 56 146 78 154
rect 0 134 78 146
rect 0 126 38 134
rect 56 126 78 134
rect 0 114 78 126
rect 0 106 38 114
rect 56 106 78 114
rect 0 94 78 106
rect 106 132 494 148
rect 106 124 291 132
rect 309 124 494 132
rect 106 116 494 124
rect 106 108 291 116
rect 309 108 494 116
rect 106 100 494 108
rect 106 96 291 100
rect 0 86 38 94
rect 56 88 78 94
rect 196 92 291 96
rect 309 96 494 100
rect 522 154 600 166
rect 522 146 544 154
rect 562 146 600 154
rect 522 134 600 146
rect 522 126 544 134
rect 562 126 600 134
rect 522 114 600 126
rect 522 106 544 114
rect 562 106 600 114
rect 309 92 404 96
rect 196 88 404 92
rect 522 94 600 106
rect 522 88 544 94
rect 56 86 544 88
rect 562 86 600 94
rect 0 84 600 86
rect 0 76 291 84
rect 309 76 600 84
rect 0 74 600 76
rect 0 66 38 74
rect 56 68 544 74
rect 56 66 291 68
rect 0 64 291 66
rect 0 54 78 64
rect 196 60 291 64
rect 309 66 544 68
rect 562 66 600 74
rect 309 64 600 66
rect 309 60 404 64
rect 196 56 404 60
rect 0 46 38 54
rect 66 46 78 54
rect 86 46 98 56
rect 106 46 118 56
rect 126 46 138 56
rect 146 46 158 56
rect 166 46 178 56
rect 186 46 414 56
rect 422 46 434 56
rect 442 46 454 56
rect 462 46 474 56
rect 482 46 494 56
rect 502 46 514 56
rect 522 54 600 64
rect 522 46 534 54
rect 562 46 600 54
rect 0 44 600 46
rect 0 36 68 44
rect 76 36 88 44
rect 96 36 108 44
rect 116 36 128 44
rect 136 36 148 44
rect 156 36 168 44
rect 176 36 188 44
rect 196 36 404 44
rect 412 36 424 44
rect 432 36 444 44
rect 452 36 464 44
rect 472 36 484 44
rect 492 36 504 44
rect 512 36 524 44
rect 532 36 600 44
rect 0 13 600 36
rect 0 -2 196 13
rect 404 -2 600 13
use PadBox  PadBox_0
timestamp 1570494029
transform 1 0 40 0 1 1480
box 0 0 520 520
<< labels >>
flabel nwell 600 -6 600 -6 6 FreeSans 16 0 0 0 VddNW
flabel nwell 0 -6 0 -6 4 FreeSans 16 0 0 0 VddNW
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 VddAct
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 VddAct
flabel psubstratepdiff 0 686 0 686 4 FreeSans 16 0 0 0 GndAct
flabel psubstratepdiff 600 686 600 686 6 FreeSans 16 0 0 0 GndAct
flabel metal1 204 -2 204 -2 4 FreeSans 64 0 0 0 Vdd
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 688 600 688 6 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 688 0 688 4 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 880 0 880 4 FreeSans 16 0 0 0 VddM2A
flabel metal2 600 880 600 880 6 FreeSans 16 0 0 0 VddM2A
flabel metal2 0 492 0 492 4 FreeSans 16 0 0 0 VddM2B
flabel metal2 600 492 600 492 6 FreeSans 16 0 0 0 VddM2B
<< properties >>
string path 220.500 2556.000 238.500 2556.000 238.500 2601.000 220.500 2601.000 220.500 2556.000 
<< end >>
