magic
tech amic5n
timestamp 1608317706
<< poly2cap >>
rect 810 240 1470 840
<< poly2capcontact >>
rect 1115 605 1165 655
<< polysilicon >>
rect 660 60 1620 1050
<< polycontact >>
rect 695 95 745 145
<< metal1 >>
rect 1080 570 1200 690
rect 660 60 780 180
<< labels >>
flabel metal1 s 690 90 690 90 2 FreeSans 400 0 0 0 a1
flabel metal1 s 1110 600 1110 600 2 FreeSans 400 0 0 0 b1
<< checkpaint >>
rect -10 -10 1630 1060
<< end >>
