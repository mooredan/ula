magic
tech amic5n
timestamp 1625766115
<< nwell >>
rect -150 550 4780 1495
<< ntransistor >>
rect 265 95 325 375
rect 455 95 515 375
rect 645 95 705 375
rect 795 95 855 375
rect 1065 95 1125 375
rect 1215 95 1275 375
rect 1410 95 1470 375
rect 1530 95 1590 375
rect 1845 95 1905 375
rect 2370 95 2430 375
rect 2975 95 3035 375
rect 3165 95 3225 375
rect 3565 95 3625 375
rect 3725 95 3785 375
rect 4135 95 4195 375
rect 4325 95 4385 375
<< ptransistor >>
rect 265 865 325 1345
rect 455 865 515 1345
rect 645 865 705 1345
rect 825 865 885 1345
rect 1065 865 1125 1345
rect 1215 865 1275 1345
rect 1410 865 1470 1345
rect 1530 865 1590 1345
rect 1845 865 1905 1345
rect 2975 865 3035 1345
rect 3165 865 3225 1345
rect 3565 865 3625 1345
rect 3725 865 3785 1345
rect 3860 865 3920 1345
rect 4135 865 4195 1345
rect 4325 865 4385 1345
<< nselect >>
rect 10 835 145 1440
rect 2025 835 2145 1440
rect 4505 835 4640 1440
rect -10 320 4660 430
rect 145 45 2555 320
rect 245 0 2555 45
rect 2690 0 4505 320
<< pselect >>
rect 145 835 2025 1440
rect 2145 835 4505 1440
rect 10 45 145 320
rect 2555 0 2690 320
rect 4505 0 4640 320
<< ndiffusion >>
rect 145 345 265 375
rect 145 295 175 345
rect 225 295 265 345
rect 145 175 265 295
rect 145 125 175 175
rect 225 125 265 175
rect 145 95 265 125
rect 325 345 455 375
rect 325 295 365 345
rect 415 295 455 345
rect 325 175 455 295
rect 325 125 365 175
rect 415 125 455 175
rect 325 95 455 125
rect 515 345 645 375
rect 515 295 555 345
rect 605 295 645 345
rect 515 175 645 295
rect 515 125 555 175
rect 605 125 645 175
rect 515 95 645 125
rect 705 95 795 375
rect 855 345 1065 375
rect 855 295 950 345
rect 1000 295 1065 345
rect 855 200 1065 295
rect 855 150 950 200
rect 1000 150 1065 200
rect 855 95 1065 150
rect 1125 95 1215 375
rect 1275 345 1410 375
rect 1275 295 1320 345
rect 1370 295 1410 345
rect 1275 175 1410 295
rect 1275 125 1320 175
rect 1370 125 1410 175
rect 1275 95 1410 125
rect 1470 95 1530 375
rect 1590 345 1845 375
rect 1590 295 1730 345
rect 1780 295 1845 345
rect 1590 95 1845 295
rect 1905 345 2025 375
rect 1905 295 1945 345
rect 1995 295 2025 345
rect 1905 95 2025 295
rect 2250 345 2370 375
rect 2250 295 2280 345
rect 2330 295 2370 345
rect 2250 185 2370 295
rect 2250 135 2280 185
rect 2330 135 2370 185
rect 2250 95 2370 135
rect 2430 345 2555 375
rect 2430 295 2470 345
rect 2520 295 2555 345
rect 2790 345 2975 375
rect 2430 175 2555 295
rect 2430 125 2470 175
rect 2520 125 2555 175
rect 2430 95 2555 125
rect 2790 295 2820 345
rect 2870 295 2975 345
rect 2790 185 2975 295
rect 2790 135 2820 185
rect 2870 135 2975 185
rect 2790 95 2975 135
rect 3035 345 3165 375
rect 3035 295 3075 345
rect 3125 295 3165 345
rect 3035 175 3165 295
rect 3035 125 3075 175
rect 3125 125 3165 175
rect 3035 95 3165 125
rect 3225 345 3355 375
rect 3225 295 3275 345
rect 3325 295 3355 345
rect 3225 175 3355 295
rect 3225 125 3275 175
rect 3325 125 3355 175
rect 3225 95 3355 125
rect 3445 345 3565 375
rect 3445 295 3475 345
rect 3525 295 3565 345
rect 3445 95 3565 295
rect 3625 95 3725 375
rect 3785 345 4135 375
rect 3785 295 4035 345
rect 4085 295 4135 345
rect 3785 175 4135 295
rect 3785 125 4035 175
rect 4085 125 4135 175
rect 3785 95 4135 125
rect 4195 345 4325 375
rect 4195 295 4235 345
rect 4285 295 4325 345
rect 4195 175 4325 295
rect 4195 125 4235 175
rect 4285 125 4325 175
rect 4195 95 4325 125
rect 4385 345 4505 375
rect 4385 295 4425 345
rect 4475 295 4505 345
rect 4385 175 4505 295
rect 4385 125 4425 175
rect 4475 125 4505 175
rect 4385 95 4505 125
<< pdiffusion >>
rect 145 1315 265 1345
rect 145 1265 175 1315
rect 225 1265 265 1315
rect 145 1195 265 1265
rect 145 1145 175 1195
rect 225 1145 265 1195
rect 145 1070 265 1145
rect 145 1020 175 1070
rect 225 1020 265 1070
rect 145 945 265 1020
rect 145 895 175 945
rect 225 895 265 945
rect 145 865 265 895
rect 325 1315 455 1345
rect 325 1265 365 1315
rect 415 1265 455 1315
rect 325 1195 455 1265
rect 325 1145 365 1195
rect 415 1145 455 1195
rect 325 1070 455 1145
rect 325 1020 365 1070
rect 415 1020 455 1070
rect 325 945 455 1020
rect 325 895 365 945
rect 415 895 455 945
rect 325 865 455 895
rect 515 1315 645 1345
rect 515 1265 555 1315
rect 605 1265 645 1315
rect 515 1200 645 1265
rect 515 1150 555 1200
rect 605 1150 645 1200
rect 515 1085 645 1150
rect 515 1035 555 1085
rect 605 1035 645 1085
rect 515 975 645 1035
rect 515 925 555 975
rect 605 925 645 975
rect 515 865 645 925
rect 705 865 825 1345
rect 885 1315 1065 1345
rect 885 1265 945 1315
rect 995 1265 1065 1315
rect 885 1195 1065 1265
rect 885 1145 945 1195
rect 995 1145 1065 1195
rect 885 1080 1065 1145
rect 885 1030 945 1080
rect 995 1030 1065 1080
rect 885 945 1065 1030
rect 885 895 945 945
rect 995 895 1065 945
rect 885 865 1065 895
rect 1125 865 1215 1345
rect 1275 1315 1410 1345
rect 1275 1265 1320 1315
rect 1370 1265 1410 1315
rect 1275 1200 1410 1265
rect 1275 1150 1320 1200
rect 1370 1150 1410 1200
rect 1275 1085 1410 1150
rect 1275 1035 1320 1085
rect 1370 1035 1410 1085
rect 1275 975 1410 1035
rect 1275 925 1320 975
rect 1370 925 1410 975
rect 1275 865 1410 925
rect 1470 865 1530 1345
rect 1590 1315 1845 1345
rect 1590 1265 1730 1315
rect 1780 1265 1845 1315
rect 1590 1195 1845 1265
rect 1590 1145 1730 1195
rect 1780 1145 1845 1195
rect 1590 1070 1845 1145
rect 1590 1020 1730 1070
rect 1780 1020 1845 1070
rect 1590 945 1845 1020
rect 1590 895 1730 945
rect 1780 895 1845 945
rect 1590 865 1845 895
rect 1905 1315 2025 1345
rect 1905 1265 1945 1315
rect 1995 1265 2025 1315
rect 1905 1195 2025 1265
rect 1905 1145 1945 1195
rect 1995 1145 2025 1195
rect 1905 1070 2025 1145
rect 1905 1020 1945 1070
rect 1995 1020 2025 1070
rect 1905 945 2025 1020
rect 1905 895 1945 945
rect 1995 895 2025 945
rect 1905 865 2025 895
rect 2790 1240 2975 1345
rect 2790 1190 2820 1240
rect 2870 1190 2975 1240
rect 2790 1125 2975 1190
rect 2790 1075 2820 1125
rect 2870 1075 2975 1125
rect 2790 1015 2975 1075
rect 2790 965 2820 1015
rect 2870 965 2975 1015
rect 2790 865 2975 965
rect 3035 1315 3165 1345
rect 3035 1265 3075 1315
rect 3125 1265 3165 1315
rect 3035 1200 3165 1265
rect 3035 1150 3075 1200
rect 3125 1150 3165 1200
rect 3035 1085 3165 1150
rect 3035 1035 3075 1085
rect 3125 1035 3165 1085
rect 3035 975 3165 1035
rect 3035 925 3075 975
rect 3125 925 3165 975
rect 3035 865 3165 925
rect 3225 1315 3355 1345
rect 3225 1265 3275 1315
rect 3325 1265 3355 1315
rect 3225 1195 3355 1265
rect 3225 1145 3275 1195
rect 3325 1145 3355 1195
rect 3225 1070 3355 1145
rect 3225 1020 3275 1070
rect 3325 1020 3355 1070
rect 3225 945 3355 1020
rect 3225 895 3275 945
rect 3325 895 3355 945
rect 3225 865 3355 895
rect 3445 1315 3565 1345
rect 3445 1265 3475 1315
rect 3525 1265 3565 1315
rect 3445 1195 3565 1265
rect 3445 1145 3475 1195
rect 3525 1145 3565 1195
rect 3445 1070 3565 1145
rect 3445 1020 3475 1070
rect 3525 1020 3565 1070
rect 3445 865 3565 1020
rect 3625 865 3725 1345
rect 3785 865 3860 1345
rect 3920 1315 4135 1345
rect 3920 1265 4030 1315
rect 4080 1265 4135 1315
rect 3920 1195 4135 1265
rect 3920 1145 4030 1195
rect 4080 1145 4135 1195
rect 3920 1070 4135 1145
rect 3920 1020 4030 1070
rect 4080 1020 4135 1070
rect 3920 945 4135 1020
rect 3920 895 4030 945
rect 4080 895 4135 945
rect 3920 865 4135 895
rect 4195 1315 4325 1345
rect 4195 1265 4235 1315
rect 4285 1265 4325 1315
rect 4195 1195 4325 1265
rect 4195 1145 4235 1195
rect 4285 1145 4325 1195
rect 4195 1070 4325 1145
rect 4195 1020 4235 1070
rect 4285 1020 4325 1070
rect 4195 945 4325 1020
rect 4195 895 4235 945
rect 4285 895 4325 945
rect 4195 865 4325 895
rect 4385 1315 4505 1345
rect 4385 1265 4425 1315
rect 4475 1265 4505 1315
rect 4385 1195 4505 1265
rect 4385 1145 4425 1195
rect 4475 1145 4505 1195
rect 4385 1070 4505 1145
rect 4385 1020 4425 1070
rect 4475 1020 4505 1070
rect 4385 945 4505 1020
rect 4385 895 4425 945
rect 4475 895 4505 945
rect 4385 865 4505 895
<< psubstratepdiff >>
rect 45 290 145 320
rect 45 240 75 290
rect 125 240 145 290
rect 45 175 145 240
rect 45 125 75 175
rect 125 125 145 175
rect 45 95 145 125
rect 2555 290 2655 320
rect 2555 240 2575 290
rect 2625 240 2655 290
rect 2555 175 2655 240
rect 2555 125 2575 175
rect 2625 125 2655 175
rect 2555 95 2655 125
rect 4505 290 4605 320
rect 4505 240 4525 290
rect 4575 240 4605 290
rect 4505 175 4605 240
rect 4505 125 4525 175
rect 4575 125 4605 175
rect 4505 95 4605 125
<< nsubstratendiff >>
rect 45 1315 145 1345
rect 45 1265 75 1315
rect 125 1265 145 1315
rect 45 1195 145 1265
rect 45 1145 75 1195
rect 125 1145 145 1195
rect 45 1070 145 1145
rect 45 1020 75 1070
rect 125 1020 145 1070
rect 45 945 145 1020
rect 45 895 75 945
rect 125 895 145 945
rect 45 865 145 895
rect 2025 1315 2125 1345
rect 2025 1265 2045 1315
rect 2095 1265 2125 1315
rect 2025 1195 2125 1265
rect 2025 1145 2045 1195
rect 2095 1145 2125 1195
rect 2025 1070 2125 1145
rect 2025 1020 2045 1070
rect 2095 1020 2125 1070
rect 2025 865 2125 1020
rect 4505 1315 4605 1345
rect 4505 1265 4525 1315
rect 4575 1265 4605 1315
rect 4505 1195 4605 1265
rect 4505 1145 4525 1195
rect 4575 1145 4605 1195
rect 4505 1070 4605 1145
rect 4505 1020 4525 1070
rect 4575 1020 4605 1070
rect 4505 945 4605 1020
rect 4505 895 4525 945
rect 4575 895 4605 945
rect 4505 865 4605 895
<< nsubstratencontact >>
rect 75 1265 125 1315
rect 75 1145 125 1195
rect 75 1020 125 1070
rect 75 895 125 945
rect 2045 1265 2095 1315
rect 2045 1145 2095 1195
rect 2045 1020 2095 1070
rect 4525 1265 4575 1315
rect 4525 1145 4575 1195
rect 4525 1020 4575 1070
rect 4525 895 4575 945
<< psubstratepcontact >>
rect 75 240 125 290
rect 75 125 125 175
rect 2575 240 2625 290
rect 2575 125 2625 175
rect 4525 240 4575 290
rect 4525 125 4575 175
<< ndcontact >>
rect 175 295 225 345
rect 175 125 225 175
rect 365 295 415 345
rect 365 125 415 175
rect 555 295 605 345
rect 555 125 605 175
rect 950 295 1000 345
rect 950 150 1000 200
rect 1320 295 1370 345
rect 1320 125 1370 175
rect 1730 295 1780 345
rect 1945 295 1995 345
rect 2280 295 2330 345
rect 2280 135 2330 185
rect 2470 295 2520 345
rect 2470 125 2520 175
rect 2820 295 2870 345
rect 2820 135 2870 185
rect 3075 295 3125 345
rect 3075 125 3125 175
rect 3275 295 3325 345
rect 3275 125 3325 175
rect 3475 295 3525 345
rect 4035 295 4085 345
rect 4035 125 4085 175
rect 4235 295 4285 345
rect 4235 125 4285 175
rect 4425 295 4475 345
rect 4425 125 4475 175
<< pdcontact >>
rect 175 1265 225 1315
rect 175 1145 225 1195
rect 175 1020 225 1070
rect 175 895 225 945
rect 365 1265 415 1315
rect 365 1145 415 1195
rect 365 1020 415 1070
rect 365 895 415 945
rect 555 1265 605 1315
rect 555 1150 605 1200
rect 555 1035 605 1085
rect 555 925 605 975
rect 945 1265 995 1315
rect 945 1145 995 1195
rect 945 1030 995 1080
rect 945 895 995 945
rect 1320 1265 1370 1315
rect 1320 1150 1370 1200
rect 1320 1035 1370 1085
rect 1320 925 1370 975
rect 1730 1265 1780 1315
rect 1730 1145 1780 1195
rect 1730 1020 1780 1070
rect 1730 895 1780 945
rect 1945 1265 1995 1315
rect 1945 1145 1995 1195
rect 1945 1020 1995 1070
rect 1945 895 1995 945
rect 2820 1190 2870 1240
rect 2820 1075 2870 1125
rect 2820 965 2870 1015
rect 3075 1265 3125 1315
rect 3075 1150 3125 1200
rect 3075 1035 3125 1085
rect 3075 925 3125 975
rect 3275 1265 3325 1315
rect 3275 1145 3325 1195
rect 3275 1020 3325 1070
rect 3275 895 3325 945
rect 3475 1265 3525 1315
rect 3475 1145 3525 1195
rect 3475 1020 3525 1070
rect 4030 1265 4080 1315
rect 4030 1145 4080 1195
rect 4030 1020 4080 1070
rect 4030 895 4080 945
rect 4235 1265 4285 1315
rect 4235 1145 4285 1195
rect 4235 1020 4285 1070
rect 4235 895 4285 945
rect 4425 1265 4475 1315
rect 4425 1145 4475 1195
rect 4425 1020 4475 1070
rect 4425 895 4475 945
<< polysilicon >>
rect 265 1345 325 1410
rect 455 1345 515 1410
rect 645 1345 705 1410
rect 825 1345 885 1410
rect 1065 1345 1125 1410
rect 1215 1345 1275 1410
rect 1410 1345 1470 1410
rect 1530 1345 1590 1410
rect 1845 1345 1905 1410
rect 2975 1345 3035 1410
rect 3165 1345 3225 1410
rect 3565 1345 3625 1410
rect 3725 1345 3785 1410
rect 3860 1345 3920 1410
rect 4135 1345 4195 1410
rect 4325 1345 4385 1410
rect 265 845 325 865
rect 455 845 515 865
rect 645 845 705 865
rect 825 845 885 865
rect 265 785 515 845
rect 615 825 705 845
rect 265 525 325 785
rect 615 775 635 825
rect 685 775 705 825
rect 615 755 705 775
rect 765 825 885 845
rect 765 775 785 825
rect 835 775 885 825
rect 765 755 885 775
rect 265 505 585 525
rect 265 455 515 505
rect 565 455 585 505
rect 265 435 585 455
rect 265 375 325 435
rect 455 375 515 435
rect 645 375 705 755
rect 1065 685 1125 865
rect 1050 665 1140 685
rect 1050 655 1070 665
rect 795 615 1070 655
rect 1120 615 1140 665
rect 795 595 1140 615
rect 795 375 855 595
rect 1215 525 1275 865
rect 1410 845 1470 865
rect 1335 825 1470 845
rect 1335 775 1355 825
rect 1405 775 1470 825
rect 1335 755 1470 775
rect 1530 845 1590 865
rect 1530 825 1620 845
rect 1530 775 1550 825
rect 1600 775 1620 825
rect 1530 755 1620 775
rect 1050 505 1140 525
rect 1050 455 1070 505
rect 1120 455 1140 505
rect 1050 435 1140 455
rect 1200 505 1290 525
rect 1200 455 1220 505
rect 1270 455 1290 505
rect 1200 435 1290 455
rect 1065 375 1125 435
rect 1215 375 1275 435
rect 1410 375 1470 755
rect 1845 685 1905 865
rect 2975 845 3035 865
rect 3165 845 3225 865
rect 2940 825 3035 845
rect 2940 775 2965 825
rect 3015 775 3035 825
rect 2940 755 3035 775
rect 3105 825 3225 845
rect 3105 775 3125 825
rect 3175 775 3225 825
rect 3105 755 3225 775
rect 3565 845 3625 865
rect 3565 825 3665 845
rect 3565 775 3595 825
rect 3645 775 3665 825
rect 3565 755 3665 775
rect 1830 665 1920 685
rect 1830 615 1850 665
rect 1900 615 1920 665
rect 1830 595 1920 615
rect 1530 505 1620 525
rect 1530 455 1550 505
rect 1600 455 1620 505
rect 1530 435 1620 455
rect 1830 505 1920 525
rect 1830 455 1850 505
rect 1900 455 1920 505
rect 1830 435 1920 455
rect 2370 505 2490 525
rect 2370 455 2420 505
rect 2470 455 2490 505
rect 2370 435 2490 455
rect 1530 375 1590 435
rect 1845 375 1905 435
rect 2370 375 2430 435
rect 2975 375 3035 755
rect 3165 375 3225 755
rect 3725 685 3785 865
rect 3860 845 3920 865
rect 4135 845 4195 865
rect 4325 845 4385 865
rect 3860 825 3950 845
rect 3860 775 3880 825
rect 3930 775 3950 825
rect 3860 755 3950 775
rect 4135 785 4385 845
rect 4135 685 4195 785
rect 3565 665 3655 685
rect 3565 615 3585 665
rect 3635 615 3655 665
rect 3565 595 3655 615
rect 3725 665 4195 685
rect 3725 615 3760 665
rect 3810 615 4085 665
rect 4135 615 4195 665
rect 3725 595 4195 615
rect 3565 375 3625 595
rect 3725 375 3785 595
rect 4135 455 4195 595
rect 4135 395 4385 455
rect 4135 375 4195 395
rect 4325 375 4385 395
rect 265 30 325 95
rect 455 30 515 95
rect 645 30 705 95
rect 795 30 855 95
rect 1065 30 1125 95
rect 1215 30 1275 95
rect 1410 30 1470 95
rect 1530 30 1590 95
rect 1845 30 1905 95
rect 2370 30 2430 95
rect 2975 30 3035 95
rect 3165 30 3225 95
rect 3565 30 3625 95
rect 3725 30 3785 95
rect 4135 30 4195 95
rect 4325 30 4385 95
<< polycontact >>
rect 635 775 685 825
rect 785 775 835 825
rect 515 455 565 505
rect 1070 615 1120 665
rect 1355 775 1405 825
rect 1550 775 1600 825
rect 1070 455 1120 505
rect 1220 455 1270 505
rect 2965 775 3015 825
rect 3125 775 3175 825
rect 3595 775 3645 825
rect 1850 615 1900 665
rect 1550 455 1600 505
rect 1850 455 1900 505
rect 2420 455 2470 505
rect 3880 775 3930 825
rect 3585 615 3635 665
rect 3760 615 3810 665
rect 4085 615 4135 665
<< metal1 >>
rect 0 1395 4650 1485
rect 55 1315 245 1395
rect 55 1265 75 1315
rect 125 1265 175 1315
rect 225 1265 245 1315
rect 55 1195 245 1265
rect 55 1145 75 1195
rect 125 1145 175 1195
rect 225 1145 245 1195
rect 55 1070 245 1145
rect 55 1020 75 1070
rect 125 1020 175 1070
rect 225 1020 245 1070
rect 55 945 245 1020
rect 55 895 75 945
rect 125 895 175 945
rect 225 895 245 945
rect 55 875 245 895
rect 345 1315 435 1335
rect 345 1265 365 1315
rect 415 1265 435 1315
rect 345 1195 435 1265
rect 345 1145 365 1195
rect 415 1145 435 1195
rect 345 1070 435 1145
rect 345 1020 365 1070
rect 415 1020 435 1070
rect 345 945 435 1020
rect 345 895 365 945
rect 415 895 435 945
rect 535 1315 625 1395
rect 535 1265 555 1315
rect 605 1265 625 1315
rect 535 1200 625 1265
rect 535 1150 555 1200
rect 605 1150 625 1200
rect 535 1085 625 1150
rect 535 1035 555 1085
rect 605 1035 625 1085
rect 535 975 625 1035
rect 535 925 555 975
rect 605 925 625 975
rect 535 905 625 925
rect 915 1315 1020 1335
rect 915 1265 945 1315
rect 995 1265 1020 1315
rect 915 1195 1020 1265
rect 915 1145 945 1195
rect 995 1145 1020 1195
rect 915 1080 1020 1145
rect 915 1030 945 1080
rect 995 1030 1020 1080
rect 915 945 1020 1030
rect 345 685 435 895
rect 915 895 945 945
rect 995 895 1020 945
rect 1300 1315 1390 1395
rect 1300 1265 1320 1315
rect 1370 1265 1390 1315
rect 1300 1200 1390 1265
rect 1300 1150 1320 1200
rect 1370 1150 1390 1200
rect 1680 1315 1800 1335
rect 1680 1265 1730 1315
rect 1780 1265 1800 1315
rect 1680 1195 1800 1265
rect 1300 1085 1390 1150
rect 1300 1035 1320 1085
rect 1370 1035 1390 1085
rect 1300 975 1390 1035
rect 1300 925 1320 975
rect 1370 925 1390 975
rect 1300 905 1390 925
rect 1530 1145 1620 1165
rect 1530 1095 1550 1145
rect 1600 1095 1620 1145
rect 915 845 1020 895
rect 505 825 705 845
rect 505 775 635 825
rect 685 775 705 825
rect 505 755 705 775
rect 765 825 855 845
rect 765 775 785 825
rect 835 775 855 825
rect 345 665 545 685
rect 345 615 365 665
rect 415 615 475 665
rect 525 615 545 665
rect 345 595 545 615
rect 145 345 245 365
rect 145 310 175 345
rect 55 295 175 310
rect 225 295 245 345
rect 55 290 245 295
rect 55 240 75 290
rect 125 240 245 290
rect 55 175 245 240
rect 55 125 75 175
rect 125 125 175 175
rect 225 125 245 175
rect 55 45 245 125
rect 345 345 435 595
rect 765 525 855 775
rect 495 505 855 525
rect 495 455 515 505
rect 565 455 645 505
rect 695 455 785 505
rect 835 455 855 505
rect 495 435 855 455
rect 915 825 1425 845
rect 915 775 1355 825
rect 1405 775 1425 825
rect 915 755 1425 775
rect 1530 825 1620 1095
rect 1530 775 1550 825
rect 1600 775 1620 825
rect 1530 755 1620 775
rect 1680 1145 1730 1195
rect 1780 1145 1800 1195
rect 1680 1070 1800 1145
rect 1680 1020 1730 1070
rect 1780 1020 1800 1070
rect 1680 945 1800 1020
rect 1680 895 1730 945
rect 1780 895 1800 945
rect 1680 865 1800 895
rect 1925 1315 2115 1335
rect 1925 1265 1945 1315
rect 1995 1265 2045 1315
rect 2095 1265 2115 1315
rect 3055 1315 3145 1395
rect 1925 1195 2115 1265
rect 1925 1145 1945 1195
rect 1995 1145 2045 1195
rect 2095 1145 2115 1195
rect 1925 1070 2115 1145
rect 1925 1020 1945 1070
rect 1995 1020 2045 1070
rect 2095 1020 2115 1070
rect 1925 985 2115 1020
rect 2800 1240 2890 1270
rect 2800 1190 2820 1240
rect 2870 1190 2890 1240
rect 2800 1145 2890 1190
rect 2800 1075 2820 1145
rect 2870 1075 2890 1145
rect 2800 1015 2890 1075
rect 1925 945 2000 985
rect 1925 895 1945 945
rect 1995 935 2000 945
rect 2050 935 2115 985
rect 1995 915 2115 935
rect 2260 985 2350 1005
rect 2260 935 2280 985
rect 2330 935 2350 985
rect 2260 915 2350 935
rect 2800 965 2820 1015
rect 2870 965 2890 1015
rect 2800 920 2890 965
rect 3055 1265 3075 1315
rect 3125 1265 3145 1315
rect 3055 1200 3145 1265
rect 3055 1150 3075 1200
rect 3125 1150 3145 1200
rect 3055 1085 3145 1150
rect 3055 1035 3075 1085
rect 3125 1035 3145 1085
rect 3055 975 3145 1035
rect 3055 925 3075 975
rect 3125 925 3145 975
rect 1995 895 2060 915
rect 1925 865 2060 895
rect 915 365 990 755
rect 1680 685 1770 865
rect 1050 665 1250 685
rect 1050 615 1070 665
rect 1120 615 1180 665
rect 1230 615 1250 665
rect 1050 595 1250 615
rect 1310 595 1770 685
rect 1830 665 1920 685
rect 1830 615 1850 665
rect 1900 615 1920 665
rect 1830 595 1920 615
rect 1310 525 1400 595
rect 1050 505 1140 525
rect 1050 455 1070 505
rect 1120 455 1140 505
rect 1050 435 1140 455
rect 1200 505 1400 525
rect 1200 455 1220 505
rect 1270 455 1400 505
rect 1200 435 1400 455
rect 1530 505 1620 525
rect 1530 455 1550 505
rect 1600 455 1620 505
rect 345 295 365 345
rect 415 295 435 345
rect 345 175 435 295
rect 345 125 365 175
rect 415 125 435 175
rect 345 105 435 125
rect 535 345 625 365
rect 535 295 555 345
rect 605 295 625 345
rect 535 175 625 295
rect 535 125 555 175
rect 605 125 625 175
rect 535 45 625 125
rect 915 345 1035 365
rect 915 295 950 345
rect 1000 295 1035 345
rect 915 200 1035 295
rect 915 150 950 200
rect 1000 150 1035 200
rect 915 105 1035 150
rect 1300 345 1390 365
rect 1300 295 1320 345
rect 1370 295 1390 345
rect 1300 175 1390 295
rect 1300 125 1320 175
rect 1370 125 1390 175
rect 1300 45 1390 125
rect 1530 210 1620 455
rect 1680 375 1770 595
rect 1830 505 1920 525
rect 1830 455 1850 505
rect 1900 455 1920 505
rect 1830 435 1920 455
rect 1980 375 2060 865
rect 2120 825 2210 845
rect 2120 775 2140 825
rect 2190 775 2210 825
rect 2120 755 2210 775
rect 1680 345 1800 375
rect 1680 295 1730 345
rect 1780 295 1800 345
rect 1680 275 1800 295
rect 1925 345 2060 375
rect 1925 295 1945 345
rect 1995 295 2060 345
rect 1925 275 2060 295
rect 2130 210 2200 755
rect 2270 375 2340 915
rect 2800 525 2865 920
rect 3055 905 3145 925
rect 3255 1315 3355 1335
rect 3255 1265 3275 1315
rect 3325 1265 3355 1315
rect 3255 1195 3355 1265
rect 3255 1145 3275 1195
rect 3325 1145 3355 1195
rect 3255 1070 3355 1145
rect 3255 1020 3275 1070
rect 3325 1020 3355 1070
rect 3255 945 3355 1020
rect 3255 895 3275 945
rect 3325 895 3355 945
rect 3255 865 3355 895
rect 2940 825 3035 845
rect 2940 775 2965 825
rect 3015 775 3035 825
rect 2940 755 3035 775
rect 3105 825 3195 845
rect 3105 775 3125 825
rect 3175 775 3195 825
rect 3105 755 3195 775
rect 2400 505 2865 525
rect 2400 455 2420 505
rect 2470 455 2865 505
rect 2400 435 2865 455
rect 2800 375 2865 435
rect 3265 375 3355 865
rect 1530 120 2200 210
rect 2260 345 2350 375
rect 2260 295 2280 345
rect 2330 295 2350 345
rect 2260 185 2350 295
rect 2260 135 2280 185
rect 2330 135 2350 185
rect 2260 105 2350 135
rect 2450 345 2540 365
rect 2450 295 2470 345
rect 2520 310 2540 345
rect 2800 345 2890 375
rect 2520 295 2645 310
rect 2450 290 2645 295
rect 2450 240 2575 290
rect 2625 240 2645 290
rect 2450 175 2645 240
rect 2450 125 2470 175
rect 2520 125 2575 175
rect 2625 125 2645 175
rect 2450 45 2645 125
rect 2800 295 2820 345
rect 2870 295 2890 345
rect 2800 185 2890 295
rect 2800 135 2820 185
rect 2870 135 2890 185
rect 2800 105 2890 135
rect 3055 345 3145 365
rect 3055 295 3075 345
rect 3125 295 3145 345
rect 3055 175 3145 295
rect 3055 125 3075 175
rect 3125 125 3145 175
rect 3055 45 3145 125
rect 3255 345 3355 375
rect 3255 295 3275 345
rect 3325 295 3355 345
rect 3255 195 3355 295
rect 3415 1315 3545 1335
rect 3415 1265 3475 1315
rect 3525 1265 3545 1315
rect 3415 1195 3545 1265
rect 3415 1145 3475 1195
rect 3525 1145 3545 1195
rect 4010 1315 4100 1395
rect 4010 1265 4030 1315
rect 4080 1265 4100 1315
rect 4010 1195 4100 1265
rect 3415 1070 3545 1145
rect 3415 1020 3475 1070
rect 3525 1020 3545 1070
rect 3415 925 3545 1020
rect 3860 1145 3950 1165
rect 3860 1095 3880 1145
rect 3930 1095 3950 1145
rect 3415 825 3505 925
rect 3415 775 3435 825
rect 3485 775 3505 825
rect 3415 375 3505 775
rect 3565 825 3665 845
rect 3565 775 3595 825
rect 3645 775 3665 825
rect 3565 755 3665 775
rect 3860 825 3950 1095
rect 4010 1145 4030 1195
rect 4080 1145 4100 1195
rect 4010 1070 4100 1145
rect 4010 1020 4030 1070
rect 4080 1020 4100 1070
rect 4010 945 4100 1020
rect 4010 895 4030 945
rect 4080 895 4100 945
rect 4010 875 4100 895
rect 4215 1315 4305 1335
rect 4215 1265 4235 1315
rect 4285 1265 4305 1315
rect 4215 1195 4305 1265
rect 4215 1145 4235 1195
rect 4285 1145 4305 1195
rect 4215 1070 4305 1145
rect 4215 1020 4235 1070
rect 4285 1020 4305 1070
rect 4215 945 4305 1020
rect 4215 895 4235 945
rect 4285 895 4305 945
rect 3860 775 3880 825
rect 3930 775 3950 825
rect 3860 755 3950 775
rect 3565 665 3655 685
rect 3565 615 3585 665
rect 3635 615 3655 665
rect 3565 595 3655 615
rect 3725 665 4155 685
rect 3725 615 3760 665
rect 3810 615 4085 665
rect 4135 615 4155 665
rect 3725 595 4155 615
rect 3415 345 3545 375
rect 3415 295 3475 345
rect 3525 295 3545 345
rect 3415 275 3545 295
rect 3860 195 3950 595
rect 3255 175 3950 195
rect 3255 125 3275 175
rect 3325 125 3950 175
rect 3255 105 3950 125
rect 4015 345 4105 365
rect 4015 295 4035 345
rect 4085 295 4105 345
rect 4015 175 4105 295
rect 4015 125 4035 175
rect 4085 125 4105 175
rect 4015 45 4105 125
rect 4215 345 4305 895
rect 4405 1315 4595 1395
rect 4405 1265 4425 1315
rect 4475 1265 4525 1315
rect 4575 1265 4595 1315
rect 4405 1195 4595 1265
rect 4405 1145 4425 1195
rect 4475 1145 4525 1195
rect 4575 1145 4595 1195
rect 4405 1070 4595 1145
rect 4405 1020 4425 1070
rect 4475 1020 4525 1070
rect 4575 1020 4595 1070
rect 4405 945 4595 1020
rect 4405 895 4425 945
rect 4475 895 4525 945
rect 4575 895 4595 945
rect 4405 875 4595 895
rect 4215 295 4235 345
rect 4285 295 4305 345
rect 4215 175 4305 295
rect 4215 125 4235 175
rect 4285 125 4305 175
rect 4215 105 4305 125
rect 4405 345 4505 365
rect 4405 295 4425 345
rect 4475 310 4505 345
rect 4475 295 4595 310
rect 4405 290 4595 295
rect 4405 240 4525 290
rect 4575 240 4595 290
rect 4405 175 4595 240
rect 4405 125 4425 175
rect 4475 125 4525 175
rect 4575 125 4595 175
rect 4405 45 4595 125
rect 0 -45 4650 45
<< via1 >>
rect 1550 1095 1600 1145
rect 365 615 415 665
rect 475 615 525 665
rect 515 455 565 505
rect 645 455 695 505
rect 785 455 835 505
rect 2820 1125 2870 1145
rect 2820 1095 2870 1125
rect 2000 935 2050 985
rect 2280 935 2330 985
rect 1070 615 1120 665
rect 1180 615 1230 665
rect 1850 615 1900 665
rect 1070 455 1120 505
rect 1850 455 1900 505
rect 2140 775 2190 825
rect 2965 775 3015 825
rect 3125 775 3175 825
rect 3880 1095 3930 1145
rect 3435 775 3485 825
rect 3595 775 3645 825
rect 3585 615 3635 665
<< metal2 >>
rect 1530 1145 3950 1165
rect 1530 1095 1550 1145
rect 1600 1095 2820 1145
rect 2870 1095 3880 1145
rect 3930 1095 3950 1145
rect 1530 1075 3950 1095
rect 1980 985 3195 1005
rect 1980 935 2000 985
rect 2050 935 2280 985
rect 2330 935 3195 985
rect 1980 915 3195 935
rect 3105 845 3195 915
rect 2120 825 3035 845
rect 2120 775 2140 825
rect 2190 775 2965 825
rect 3015 775 3035 825
rect 2120 755 3035 775
rect 3105 825 3505 845
rect 3105 775 3125 825
rect 3175 775 3435 825
rect 3485 775 3505 825
rect 3105 755 3505 775
rect 3575 825 3815 845
rect 3575 775 3595 825
rect 3645 775 3815 825
rect 3575 755 3815 775
rect 345 665 3655 685
rect 345 615 365 665
rect 415 615 475 665
rect 525 615 1070 665
rect 1120 615 1180 665
rect 1230 615 1850 665
rect 1900 615 3585 665
rect 3635 615 3655 665
rect 345 595 3655 615
rect 3725 525 3815 755
rect 495 505 3815 525
rect 495 455 515 505
rect 565 455 645 505
rect 695 455 785 505
rect 835 455 1070 505
rect 1120 455 1850 505
rect 1900 455 3815 505
rect 495 435 3815 455
<< labels >>
flabel ndiffusion s 1155 195 1155 195 2 FreeSans 400 0 0 0 x6
flabel ndiffusion 735 195 735 195 2 FreeSans 400 0 0 0 x5
flabel metal1 s 945 165 945 165 2 FreeSans 400 0 0 0 nmas
flabel metal1 360 610 360 610 2 FreeSans 400 0 0 0 nck
flabel metal1 s 515 800 515 800 2 FreeSans 400 0 0 0 d
port 1 s
flabel metal1 s 555 1395 555 1395 2 FreeSans 400 0 0 0 vdd
port 3 n
flabel pdiffusion s 1155 1065 1155 1065 2 FreeSans 400 0 0 0 x2
flabel pdiffusion s 765 1065 765 1065 2 FreeSans 400 0 0 0 x1
flabel metal1 s 1215 770 1215 770 2 FreeSans 400 0 0 0 nmas
flabel metal1 s 1050 465 1050 465 2 FreeSans 400 0 0 0 ck
port 2 ne
flabel metal1 s 945 925 945 925 2 FreeSans 400 0 0 0 nmas
flabel metal1 s 1740 1065 1740 1065 2 FreeSans 400 0 0 0 mas
flabel metal1 s 1725 285 1725 285 2 FreeSans 400 0 0 0 mas
flabel metal1 s 1986 770 1986 770 8 FreeSans 400 180 0 0 slv
flabel metal1 s 1986 940 1986 940 8 FreeSans 400 180 0 0 slv
flabel metal1 s 175 15 175 15 2 FreeSans 400 0 0 0 vss
port 4 s
flabel nwell s 2895 600 2895 600 2 FreeSans 400 0 0 0 vdd
flabel pdiffusion s 3655 1185 3655 1185 2 FreeSans 400 0 0 0 x4
flabel metal1 s 3795 640 3795 640 2 FreeSans 400 0 0 0 nslv
flabel ndiffusion s 3640 150 3640 150 2 FreeSans 400 0 0 0 x8
flabel metal1 s 4235 710 4235 710 2 FreeSans 400 0 0 0 q
port 0 e
<< properties >>
string LEFclass CORE
string LEFsite core
string FIXED_BBOX 0 0 3150 1440
string LEFsymmetry X Y
<< end >>
