magic
tech scmos
timestamp 1511733589
<< nwell >>
rect -1 24 52 65
<< nselect >>
rect 6 46 32 61
rect 6 2 27 19
rect 34 2 48 19
<< pselect >>
rect 32 46 48 61
rect 6 30 48 46
rect 32 28 48 30
rect 27 2 34 19
<< ntransistor >>
rect 13 4 15 17
rect 18 4 20 17
rect 39 4 41 17
<< ptransistor >>
rect 13 32 15 43
rect 21 32 23 43
rect 39 30 41 59
<< ndiffusion >>
rect 8 4 13 17
rect 15 4 18 17
rect 20 4 25 17
rect 34 4 39 17
rect 41 4 46 17
<< pdiffusion >>
rect 8 32 13 43
rect 15 32 21 43
rect 23 32 28 43
rect 34 30 39 59
rect 41 30 46 59
<< psubstratepdiff >>
rect 29 4 34 17
<< nsubstratendiff >>
rect 15 47 21 58
<< polysilicon >>
rect 39 59 41 61
rect 13 43 15 45
rect 21 43 23 45
rect 13 24 15 32
rect 8 18 15 24
rect 21 24 23 32
rect 39 24 41 30
rect 21 20 28 24
rect 13 17 15 18
rect 18 18 28 20
rect 34 18 41 24
rect 18 17 20 18
rect 39 17 41 18
rect 13 2 15 4
rect 18 2 20 4
rect 39 2 41 4
<< genericcontact >>
rect 17 55 19 57
rect 35 55 37 57
rect 43 53 45 55
rect 35 50 37 52
rect 35 44 37 46
rect 43 44 45 46
rect 9 39 11 41
rect 17 40 19 42
rect 25 39 27 41
rect 35 39 37 41
rect 43 38 45 40
rect 9 34 11 36
rect 17 34 19 36
rect 25 34 27 36
rect 35 34 37 36
rect 43 32 45 34
rect 10 20 12 22
rect 24 20 26 22
rect 36 20 38 22
rect 9 13 11 15
rect 22 13 24 15
rect 30 13 32 15
rect 35 13 37 15
rect 43 13 45 15
rect 9 6 11 8
rect 22 7 24 9
rect 43 7 45 9
rect 30 5 32 7
rect 35 5 37 7
<< metal1 >>
rect 5 60 46 63
rect 8 33 12 60
rect 16 54 20 60
rect 16 30 20 43
rect 24 33 28 60
rect 34 33 38 60
rect 16 26 39 30
rect 9 19 13 23
rect 16 16 20 26
rect 23 19 31 23
rect 35 19 39 26
rect 8 3 12 16
rect 16 12 25 16
rect 21 6 25 12
rect 29 3 38 16
rect 42 6 46 57
rect 5 0 46 3
<< bb >>
rect 0 0 51 63
<< labels >>
rlabel metal1 42 6 46 57 0 z
port 1 e
rlabel metal1 9 19 13 23 0 a
port 2 nw
rlabel metal1 23 19 31 23 0 b
port 3 nsew
rlabel metal1 5 60 46 63 0 Vdd
port 4 new
rlabel metal1 5 0 46 3 0 Gnd
port 5 sew
rlabel ndiffusion 16 8 16 8 2 x1
rlabel nwell 3 25 3 25 2 Vdd
<< end >>
