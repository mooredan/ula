magic
tech amic5n
timestamp 1624361752
<< nwell >>
rect -130 550 580 1495
<< ntransistor >>
rect 225 95 285 400
<< ptransistor >>
rect 225 705 285 1345
<< nselect >>
rect -10 0 460 430
<< pselect >>
rect -10 670 460 1440
<< ndiffusion >>
rect 105 370 225 400
rect 105 320 135 370
rect 185 320 225 370
rect 105 175 225 320
rect 105 125 135 175
rect 185 125 225 175
rect 105 95 225 125
rect 285 370 405 400
rect 285 320 325 370
rect 375 320 405 370
rect 285 175 405 320
rect 285 125 325 175
rect 375 125 405 175
rect 285 95 405 125
<< pdiffusion >>
rect 105 1315 225 1345
rect 105 1265 135 1315
rect 185 1265 225 1315
rect 105 1215 225 1265
rect 105 1165 135 1215
rect 185 1165 225 1215
rect 105 1115 225 1165
rect 105 1065 135 1115
rect 185 1065 225 1115
rect 105 1015 225 1065
rect 105 965 135 1015
rect 185 965 225 1015
rect 105 915 225 965
rect 105 865 135 915
rect 185 865 225 915
rect 105 815 225 865
rect 105 765 135 815
rect 185 765 225 815
rect 105 705 225 765
rect 285 1315 405 1345
rect 285 1265 325 1315
rect 375 1265 405 1315
rect 285 1185 405 1265
rect 285 1135 325 1185
rect 375 1135 405 1185
rect 285 1085 405 1135
rect 285 1035 325 1085
rect 375 1035 405 1085
rect 285 985 405 1035
rect 285 935 325 985
rect 375 935 405 985
rect 285 885 405 935
rect 285 835 325 885
rect 375 835 405 885
rect 285 785 405 835
rect 285 735 325 785
rect 375 735 405 785
rect 285 705 405 735
<< ndcontact >>
rect 135 320 185 370
rect 135 125 185 175
rect 325 320 375 370
rect 325 125 375 175
<< pdcontact >>
rect 135 1265 185 1315
rect 135 1165 185 1215
rect 135 1065 185 1115
rect 135 965 185 1015
rect 135 865 185 915
rect 135 765 185 815
rect 325 1265 375 1315
rect 325 1135 375 1185
rect 325 1035 375 1085
rect 325 935 375 985
rect 325 835 375 885
rect 325 735 375 785
<< polysilicon >>
rect 225 1345 285 1410
rect 225 685 285 705
rect 115 665 285 685
rect 115 615 135 665
rect 185 615 285 665
rect 115 595 285 615
rect 225 400 285 595
rect 225 30 285 95
<< polycontact >>
rect 135 615 185 665
<< metal1 >>
rect 0 1395 450 1485
rect 115 1315 205 1395
rect 115 1265 135 1315
rect 185 1265 205 1315
rect 115 1215 205 1265
rect 115 1165 135 1215
rect 185 1165 205 1215
rect 115 1115 205 1165
rect 115 1065 135 1115
rect 185 1065 205 1115
rect 115 1015 205 1065
rect 115 965 135 1015
rect 185 965 205 1015
rect 115 915 205 965
rect 115 865 135 915
rect 185 865 205 915
rect 115 815 205 865
rect 115 765 135 815
rect 185 765 205 815
rect 115 745 205 765
rect 305 1315 395 1335
rect 305 1265 325 1315
rect 375 1265 395 1315
rect 305 1185 395 1265
rect 305 1135 325 1185
rect 375 1135 395 1185
rect 305 1085 395 1135
rect 305 1035 325 1085
rect 375 1035 395 1085
rect 305 985 395 1035
rect 305 935 325 985
rect 375 935 395 985
rect 305 885 395 935
rect 305 835 325 885
rect 375 835 395 885
rect 305 785 395 835
rect 305 735 325 785
rect 375 735 395 785
rect 305 685 395 735
rect 115 665 395 685
rect 115 615 135 665
rect 185 615 395 665
rect 115 595 395 615
rect 115 370 205 390
rect 115 320 135 370
rect 185 320 205 370
rect 115 175 205 320
rect 115 125 135 175
rect 185 125 205 175
rect 115 45 205 125
rect 305 370 395 525
rect 305 320 325 370
rect 375 320 395 370
rect 305 175 395 320
rect 305 125 325 175
rect 375 125 395 175
rect 305 105 395 125
rect 0 -45 450 45
<< labels >>
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 1 ne
flabel nwell 395 600 395 600 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 335 470 335 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 2 ne
<< properties >>
string FIXED_BBOX 0 0 450 1440
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
<< end >>
