magic
tech scmos
magscale 1 2
timestamp 1570494029
<< error_p >>
rect 12 1316 14 1324
rect 20 1316 22 1318
rect 8 1314 10 1316
rect 14 1314 16 1316
rect 18 1314 22 1316
rect 10 1312 14 1314
rect 562 1302 564 1304
rect 36 1300 38 1302
rect 564 1300 566 1302
rect 34 1298 36 1300
rect 58 1282 60 1284
rect 60 1280 62 1282
rect 102 1105 104 1107
rect 100 1103 102 1105
rect 404 781 415 782
rect 586 703 598 705
rect 588 701 590 703
rect 94 700 96 701
rect 126 700 128 701
rect 132 700 134 701
rect 158 700 160 701
rect 164 700 166 701
rect 222 700 224 701
rect 228 700 230 701
rect 588 697 590 699
rect 590 695 592 697
rect 549 683 550 684
rect 555 670 556 671
rect 588 656 590 658
rect 590 654 592 656
rect 580 543 590 544
rect 580 541 592 543
rect 588 539 590 541
rect 588 536 590 538
rect 158 533 160 535
rect 164 533 166 535
rect 392 533 394 535
rect 482 533 484 535
rect 488 533 490 535
rect 578 534 580 535
rect 586 534 588 536
rect 578 533 590 534
rect 580 531 592 533
rect 588 529 590 531
rect 588 526 590 528
rect 586 524 588 526
rect 580 521 582 523
rect 216 518 218 520
rect 482 519 484 521
rect 488 519 490 521
rect 578 519 580 521
rect 218 516 220 518
rect 480 517 482 519
rect 490 517 492 519
rect 208 514 220 516
rect 216 512 218 514
rect 216 508 218 510
rect 214 506 216 508
rect 590 502 592 504
rect 588 500 590 502
rect 106 468 108 470
rect 126 468 128 470
rect 136 468 138 470
rect 156 468 158 470
rect 166 468 168 470
rect 186 468 188 470
rect 196 468 198 470
rect 216 468 218 470
rect 226 468 228 470
rect 234 468 236 476
rect 382 468 384 470
rect 392 468 394 470
rect 412 468 414 470
rect 422 468 424 470
rect 442 468 444 470
rect 452 468 454 470
rect 472 468 474 470
rect 482 468 484 470
rect 52 466 54 468
rect 108 466 110 468
rect 124 466 126 468
rect 138 466 140 468
rect 154 466 156 468
rect 168 466 170 468
rect 184 466 186 468
rect 198 466 200 468
rect 214 466 216 468
rect 228 466 230 468
rect 232 466 236 468
rect 380 466 382 468
rect 394 466 396 468
rect 410 466 412 468
rect 424 466 426 468
rect 440 466 442 468
rect 454 466 456 468
rect 470 466 472 468
rect 484 466 486 468
rect 50 464 52 466
rect 234 464 236 466
rect 68 60 78 64
rect 68 58 80 60
rect 76 56 78 58
rect 74 54 76 56
rect 68 50 78 54
rect 68 48 80 50
rect 76 46 78 48
rect 74 44 76 46
rect 68 40 78 44
rect 68 38 80 40
rect 76 36 78 38
rect 74 34 76 36
rect 578 14 580 22
rect 586 14 590 16
rect 580 12 582 14
rect 584 12 588 14
rect 590 12 592 14
rect 10 10 22 12
rect 46 10 58 12
rect 72 10 84 12
rect 106 10 118 12
rect 474 10 486 12
rect 528 10 540 12
rect 578 10 580 12
rect 12 8 14 10
rect 54 8 56 10
rect 74 8 76 10
rect 114 8 116 10
rect 476 8 478 10
rect 536 8 538 10
rect 12 4 14 6
rect 54 4 56 6
rect 74 4 76 6
rect 114 4 116 6
rect 476 4 478 6
rect 536 4 538 6
rect 14 2 16 4
rect 52 2 54 4
rect 76 2 78 4
rect 112 2 114 4
rect 478 2 480 4
rect 534 2 536 4
<< error_s >>
rect 110 1598 118 1600
rect 134 1598 142 1600
rect 158 1598 166 1600
rect 182 1598 190 1600
rect 206 1598 214 1600
rect 230 1598 238 1600
rect 254 1598 262 1600
rect 278 1598 286 1600
rect 302 1598 310 1600
rect 326 1598 334 1600
rect 350 1598 358 1600
rect 374 1598 382 1600
rect 398 1598 406 1600
rect 422 1598 430 1600
rect 446 1598 454 1600
rect 470 1598 478 1600
rect 494 1598 502 1600
rect 98 1592 106 1594
rect 98 1588 100 1592
rect 104 1588 106 1592
rect 98 1586 106 1588
rect 122 1592 130 1594
rect 122 1588 124 1592
rect 128 1588 130 1592
rect 122 1586 130 1588
rect 146 1592 154 1594
rect 146 1588 148 1592
rect 152 1588 154 1592
rect 146 1586 154 1588
rect 170 1592 178 1594
rect 170 1588 172 1592
rect 176 1588 178 1592
rect 170 1586 178 1588
rect 194 1592 202 1594
rect 194 1588 196 1592
rect 200 1588 202 1592
rect 194 1586 202 1588
rect 218 1592 226 1594
rect 218 1588 220 1592
rect 224 1588 226 1592
rect 218 1586 226 1588
rect 242 1592 250 1594
rect 242 1588 244 1592
rect 248 1588 250 1592
rect 242 1586 250 1588
rect 266 1592 274 1594
rect 266 1588 268 1592
rect 272 1588 274 1592
rect 266 1586 274 1588
rect 290 1592 298 1594
rect 290 1588 292 1592
rect 296 1588 298 1592
rect 290 1586 298 1588
rect 314 1592 322 1594
rect 314 1588 316 1592
rect 320 1588 322 1592
rect 314 1586 322 1588
rect 338 1592 346 1594
rect 338 1588 340 1592
rect 344 1588 346 1592
rect 338 1586 346 1588
rect 362 1592 370 1594
rect 362 1588 364 1592
rect 368 1588 370 1592
rect 362 1586 370 1588
rect 386 1592 394 1594
rect 386 1588 388 1592
rect 392 1588 394 1592
rect 386 1586 394 1588
rect 410 1592 418 1594
rect 410 1588 412 1592
rect 416 1588 418 1592
rect 410 1586 418 1588
rect 434 1592 442 1594
rect 434 1588 436 1592
rect 440 1588 442 1592
rect 434 1586 442 1588
rect 458 1592 466 1594
rect 458 1588 460 1592
rect 464 1588 466 1592
rect 458 1586 466 1588
rect 482 1592 490 1594
rect 482 1588 484 1592
rect 488 1588 490 1592
rect 482 1586 490 1588
rect 110 1580 118 1582
rect 110 1576 112 1580
rect 116 1576 118 1580
rect 110 1574 118 1576
rect 134 1580 142 1582
rect 134 1576 136 1580
rect 140 1576 142 1580
rect 134 1574 142 1576
rect 158 1580 166 1582
rect 158 1576 160 1580
rect 164 1576 166 1580
rect 158 1574 166 1576
rect 182 1580 190 1582
rect 182 1576 184 1580
rect 188 1576 190 1580
rect 182 1574 190 1576
rect 206 1580 214 1582
rect 206 1576 208 1580
rect 212 1576 214 1580
rect 206 1574 214 1576
rect 230 1580 238 1582
rect 230 1576 232 1580
rect 236 1576 238 1580
rect 230 1574 238 1576
rect 254 1580 262 1582
rect 254 1576 256 1580
rect 260 1576 262 1580
rect 254 1574 262 1576
rect 278 1580 286 1582
rect 278 1576 280 1580
rect 284 1576 286 1580
rect 278 1574 286 1576
rect 302 1580 310 1582
rect 302 1576 304 1580
rect 308 1576 310 1580
rect 302 1574 310 1576
rect 326 1580 334 1582
rect 326 1576 328 1580
rect 332 1576 334 1580
rect 326 1574 334 1576
rect 350 1580 358 1582
rect 350 1576 352 1580
rect 356 1576 358 1580
rect 350 1574 358 1576
rect 374 1580 382 1582
rect 374 1576 376 1580
rect 380 1576 382 1580
rect 374 1574 382 1576
rect 398 1580 406 1582
rect 398 1576 400 1580
rect 404 1576 406 1580
rect 398 1574 406 1576
rect 422 1580 430 1582
rect 422 1576 424 1580
rect 428 1576 430 1580
rect 422 1574 430 1576
rect 446 1580 454 1582
rect 446 1576 448 1580
rect 452 1576 454 1580
rect 446 1574 454 1576
rect 470 1580 478 1582
rect 470 1576 472 1580
rect 476 1576 478 1580
rect 470 1574 478 1576
rect 494 1580 502 1582
rect 494 1576 496 1580
rect 500 1576 502 1580
rect 494 1574 502 1576
rect 98 1568 106 1570
rect 98 1564 100 1568
rect 104 1564 106 1568
rect 98 1562 106 1564
rect 122 1568 130 1570
rect 122 1564 124 1568
rect 128 1564 130 1568
rect 122 1562 130 1564
rect 146 1568 154 1570
rect 146 1564 148 1568
rect 152 1564 154 1568
rect 146 1562 154 1564
rect 170 1568 178 1570
rect 170 1564 172 1568
rect 176 1564 178 1568
rect 170 1562 178 1564
rect 194 1568 202 1570
rect 194 1564 196 1568
rect 200 1564 202 1568
rect 194 1562 202 1564
rect 218 1568 226 1570
rect 218 1564 220 1568
rect 224 1564 226 1568
rect 218 1562 226 1564
rect 242 1568 250 1570
rect 242 1564 244 1568
rect 248 1564 250 1568
rect 242 1562 250 1564
rect 266 1568 274 1570
rect 266 1564 268 1568
rect 272 1564 274 1568
rect 266 1562 274 1564
rect 290 1568 298 1570
rect 290 1564 292 1568
rect 296 1564 298 1568
rect 290 1562 298 1564
rect 314 1568 322 1570
rect 314 1564 316 1568
rect 320 1564 322 1568
rect 314 1562 322 1564
rect 338 1568 346 1570
rect 338 1564 340 1568
rect 344 1564 346 1568
rect 338 1562 346 1564
rect 362 1568 370 1570
rect 362 1564 364 1568
rect 368 1564 370 1568
rect 362 1562 370 1564
rect 386 1568 394 1570
rect 386 1564 388 1568
rect 392 1564 394 1568
rect 386 1562 394 1564
rect 410 1568 418 1570
rect 410 1564 412 1568
rect 416 1564 418 1568
rect 410 1562 418 1564
rect 434 1568 442 1570
rect 434 1564 436 1568
rect 440 1564 442 1568
rect 434 1562 442 1564
rect 458 1568 466 1570
rect 458 1564 460 1568
rect 464 1564 466 1568
rect 458 1562 466 1564
rect 482 1568 490 1570
rect 482 1564 484 1568
rect 488 1564 490 1568
rect 482 1562 490 1564
rect 110 1556 118 1558
rect 110 1552 112 1556
rect 116 1552 118 1556
rect 110 1550 118 1552
rect 134 1556 142 1558
rect 134 1552 136 1556
rect 140 1552 142 1556
rect 134 1550 142 1552
rect 158 1556 166 1558
rect 158 1552 160 1556
rect 164 1552 166 1556
rect 158 1550 166 1552
rect 182 1556 190 1558
rect 182 1552 184 1556
rect 188 1552 190 1556
rect 182 1550 190 1552
rect 206 1556 214 1558
rect 206 1552 208 1556
rect 212 1552 214 1556
rect 206 1550 214 1552
rect 230 1556 238 1558
rect 230 1552 232 1556
rect 236 1552 238 1556
rect 230 1550 238 1552
rect 254 1556 262 1558
rect 254 1552 256 1556
rect 260 1552 262 1556
rect 254 1550 262 1552
rect 278 1556 286 1558
rect 278 1552 280 1556
rect 284 1552 286 1556
rect 278 1550 286 1552
rect 302 1556 310 1558
rect 302 1552 304 1556
rect 308 1552 310 1556
rect 302 1550 310 1552
rect 326 1556 334 1558
rect 326 1552 328 1556
rect 332 1552 334 1556
rect 326 1550 334 1552
rect 350 1556 358 1558
rect 350 1552 352 1556
rect 356 1552 358 1556
rect 350 1550 358 1552
rect 374 1556 382 1558
rect 374 1552 376 1556
rect 380 1552 382 1556
rect 374 1550 382 1552
rect 398 1556 406 1558
rect 398 1552 400 1556
rect 404 1552 406 1556
rect 398 1550 406 1552
rect 422 1556 430 1558
rect 422 1552 424 1556
rect 428 1552 430 1556
rect 422 1550 430 1552
rect 446 1556 454 1558
rect 446 1552 448 1556
rect 452 1552 454 1556
rect 446 1550 454 1552
rect 470 1556 478 1558
rect 470 1552 472 1556
rect 476 1552 478 1556
rect 470 1550 478 1552
rect 494 1556 502 1558
rect 494 1552 496 1556
rect 500 1552 502 1556
rect 494 1550 502 1552
rect 98 1544 106 1546
rect 98 1540 100 1544
rect 104 1540 106 1544
rect 98 1538 106 1540
rect 122 1544 130 1546
rect 122 1540 124 1544
rect 128 1540 130 1544
rect 122 1538 130 1540
rect 146 1544 154 1546
rect 146 1540 148 1544
rect 152 1540 154 1544
rect 146 1538 154 1540
rect 170 1544 178 1546
rect 170 1540 172 1544
rect 176 1540 178 1544
rect 170 1538 178 1540
rect 194 1544 202 1546
rect 194 1540 196 1544
rect 200 1540 202 1544
rect 194 1538 202 1540
rect 218 1544 226 1546
rect 218 1540 220 1544
rect 224 1540 226 1544
rect 218 1538 226 1540
rect 242 1544 250 1546
rect 242 1540 244 1544
rect 248 1540 250 1544
rect 242 1538 250 1540
rect 266 1544 274 1546
rect 266 1540 268 1544
rect 272 1540 274 1544
rect 266 1538 274 1540
rect 290 1544 298 1546
rect 290 1540 292 1544
rect 296 1540 298 1544
rect 290 1538 298 1540
rect 314 1544 322 1546
rect 314 1540 316 1544
rect 320 1540 322 1544
rect 314 1538 322 1540
rect 338 1544 346 1546
rect 338 1540 340 1544
rect 344 1540 346 1544
rect 338 1538 346 1540
rect 362 1544 370 1546
rect 362 1540 364 1544
rect 368 1540 370 1544
rect 362 1538 370 1540
rect 386 1544 394 1546
rect 386 1540 388 1544
rect 392 1540 394 1544
rect 386 1538 394 1540
rect 410 1544 418 1546
rect 410 1540 412 1544
rect 416 1540 418 1544
rect 410 1538 418 1540
rect 434 1544 442 1546
rect 434 1540 436 1544
rect 440 1540 442 1544
rect 434 1538 442 1540
rect 458 1544 466 1546
rect 458 1540 460 1544
rect 464 1540 466 1544
rect 458 1538 466 1540
rect 482 1544 490 1546
rect 482 1540 484 1544
rect 488 1540 490 1544
rect 482 1538 490 1540
<< nwell >>
rect 30 1208 572 1304
rect 28 950 572 1208
rect 28 850 570 950
rect 284 848 570 850
rect -12 507 606 677
rect -6 498 606 507
rect -6 22 22 498
rect 572 22 606 498
rect -6 -6 606 22
<< ntransistor >>
rect 38 706 42 766
rect 54 706 58 766
rect 88 706 92 766
rect 104 706 108 766
rect 120 706 124 766
rect 136 706 140 766
rect 152 706 156 766
rect 168 706 172 766
rect 184 706 188 766
rect 200 706 204 766
rect 216 706 220 766
rect 232 706 236 766
rect 248 706 252 766
rect 264 706 268 766
rect 280 706 284 766
rect 296 706 300 766
rect 396 707 400 767
rect 412 707 416 767
rect 428 707 432 767
rect 444 707 448 767
rect 460 707 464 767
rect 476 707 480 767
rect 492 707 496 767
rect 508 707 512 767
rect 524 707 528 767
rect 540 707 544 767
rect 556 707 560 767
rect 572 707 576 767
rect 76 432 276 438
rect 76 342 276 348
rect 76 300 276 306
rect 76 212 276 218
rect 76 170 276 176
rect 76 82 276 88
rect 324 432 524 438
rect 324 342 524 348
rect 324 300 524 306
rect 324 212 524 218
rect 324 170 524 176
rect 324 82 524 88
<< ptransistor >>
rect 76 1248 276 1254
rect 76 1160 276 1166
rect 76 1118 276 1124
rect 76 1032 276 1038
rect 76 990 276 996
rect 76 902 276 908
rect 324 1248 524 1254
rect 324 1160 524 1166
rect 324 1118 524 1124
rect 324 1032 524 1038
rect 324 990 524 996
rect 324 902 524 908
rect 38 539 42 643
rect 54 539 58 643
rect 88 539 92 643
rect 104 539 108 643
rect 120 539 124 643
rect 136 539 140 643
rect 152 539 156 643
rect 168 539 172 643
rect 184 539 188 643
rect 200 539 204 643
rect 216 539 220 643
rect 232 539 236 643
rect 248 539 252 643
rect 264 539 268 643
rect 280 539 284 643
rect 296 539 300 643
rect 396 539 400 643
rect 412 539 416 643
rect 428 539 432 643
rect 444 539 448 643
rect 460 539 464 643
rect 476 539 480 643
rect 492 539 496 643
rect 508 539 512 643
rect 524 539 528 643
rect 540 539 544 643
rect 556 539 560 643
rect 572 539 576 643
<< ndiffusion >>
rect 26 760 38 766
rect 26 722 28 760
rect 36 722 38 760
rect 26 706 38 722
rect 42 760 54 766
rect 42 752 44 760
rect 52 752 54 760
rect 42 740 54 752
rect 42 732 44 740
rect 52 732 54 740
rect 42 720 54 732
rect 42 712 44 720
rect 52 712 54 720
rect 42 706 54 712
rect 58 758 70 766
rect 58 710 60 758
rect 68 710 70 758
rect 58 706 70 710
rect 76 759 88 766
rect 76 721 78 759
rect 86 721 88 759
rect 76 706 88 721
rect 92 756 104 766
rect 92 748 94 756
rect 102 748 104 756
rect 92 736 104 748
rect 92 728 94 736
rect 102 728 104 736
rect 92 716 104 728
rect 92 708 94 716
rect 102 708 104 716
rect 92 706 104 708
rect 108 759 120 766
rect 108 711 110 759
rect 118 711 120 759
rect 108 706 120 711
rect 124 756 136 766
rect 124 748 126 756
rect 134 748 136 756
rect 124 736 136 748
rect 124 728 126 736
rect 134 728 136 736
rect 124 716 136 728
rect 124 708 126 716
rect 134 708 136 716
rect 124 706 136 708
rect 140 759 152 766
rect 140 711 142 759
rect 150 711 152 759
rect 140 706 152 711
rect 156 756 168 766
rect 156 748 158 756
rect 166 748 168 756
rect 156 736 168 748
rect 156 728 158 736
rect 166 728 168 736
rect 156 716 168 728
rect 156 708 158 716
rect 166 708 168 716
rect 156 706 168 708
rect 172 759 184 766
rect 172 711 174 759
rect 182 711 184 759
rect 172 706 184 711
rect 188 756 200 766
rect 188 748 190 756
rect 198 748 200 756
rect 188 736 200 748
rect 188 728 190 736
rect 198 728 200 736
rect 188 716 200 728
rect 188 708 190 716
rect 198 708 200 716
rect 188 706 200 708
rect 204 760 216 766
rect 204 712 206 760
rect 214 712 216 760
rect 204 706 216 712
rect 220 756 232 766
rect 220 748 222 756
rect 230 748 232 756
rect 220 736 232 748
rect 220 728 222 736
rect 230 728 232 736
rect 220 716 232 728
rect 220 708 222 716
rect 230 708 232 716
rect 220 706 232 708
rect 236 758 248 766
rect 236 730 238 758
rect 246 730 248 758
rect 236 706 248 730
rect 252 756 264 766
rect 252 708 254 756
rect 262 708 264 756
rect 252 706 264 708
rect 268 758 280 766
rect 268 730 270 758
rect 278 730 280 758
rect 268 718 280 730
rect 268 710 270 718
rect 278 710 280 718
rect 268 706 280 710
rect 284 763 296 766
rect 284 755 286 763
rect 294 755 296 763
rect 284 752 296 755
rect 284 744 286 752
rect 294 744 296 752
rect 284 740 296 744
rect 284 732 286 740
rect 294 732 296 740
rect 284 728 296 732
rect 284 720 286 728
rect 294 720 296 728
rect 284 706 296 720
rect 300 764 312 766
rect 300 756 302 764
rect 310 756 312 764
rect 300 752 312 756
rect 300 744 302 752
rect 310 744 312 752
rect 300 741 312 744
rect 300 733 302 741
rect 310 733 312 741
rect 300 728 312 733
rect 300 720 302 728
rect 310 720 312 728
rect 300 716 312 720
rect 300 708 302 716
rect 310 708 312 716
rect 300 706 312 708
rect 384 760 396 767
rect 384 752 386 760
rect 394 752 396 760
rect 384 740 396 752
rect 384 732 386 740
rect 394 732 396 740
rect 384 720 396 732
rect 384 712 386 720
rect 394 712 396 720
rect 384 707 396 712
rect 400 760 412 767
rect 400 712 402 760
rect 410 712 412 760
rect 400 707 412 712
rect 416 748 428 767
rect 416 730 418 748
rect 426 730 428 748
rect 416 717 428 730
rect 416 709 418 717
rect 426 709 428 717
rect 416 707 428 709
rect 432 760 444 767
rect 432 712 434 760
rect 442 712 444 760
rect 432 707 444 712
rect 448 761 460 767
rect 448 753 450 761
rect 458 753 460 761
rect 448 741 460 753
rect 448 733 450 741
rect 458 733 460 741
rect 448 721 460 733
rect 448 713 450 721
rect 458 713 460 721
rect 448 707 460 713
rect 464 761 476 767
rect 464 713 466 761
rect 474 713 476 761
rect 464 707 476 713
rect 480 761 492 767
rect 480 753 482 761
rect 490 753 492 761
rect 480 741 492 753
rect 480 733 482 741
rect 490 733 492 741
rect 480 721 492 733
rect 480 713 482 721
rect 490 713 492 721
rect 480 707 492 713
rect 496 761 508 767
rect 496 713 498 761
rect 506 713 508 761
rect 496 707 508 713
rect 512 761 524 767
rect 512 753 514 761
rect 522 753 524 761
rect 512 741 524 753
rect 512 733 514 741
rect 522 733 524 741
rect 512 721 524 733
rect 512 713 514 721
rect 522 713 524 721
rect 512 707 524 713
rect 528 761 540 767
rect 528 713 530 761
rect 538 713 540 761
rect 528 707 540 713
rect 544 761 556 767
rect 544 753 546 761
rect 554 753 556 761
rect 544 741 556 753
rect 544 733 546 741
rect 554 733 556 741
rect 544 721 556 733
rect 544 713 546 721
rect 554 713 556 721
rect 544 707 556 713
rect 560 761 572 767
rect 560 713 562 761
rect 570 713 572 761
rect 560 707 572 713
rect 576 761 582 767
rect 576 753 578 761
rect 576 741 586 753
rect 576 733 578 741
rect 576 721 586 733
rect 576 713 578 721
rect 576 707 586 713
rect 94 701 100 706
rect 126 701 134 706
rect 158 701 166 706
rect 222 701 230 706
rect 384 701 394 707
rect 418 701 426 707
rect 450 701 456 707
rect 482 701 490 707
rect 514 701 522 707
rect 546 701 552 707
rect 578 701 586 707
rect 76 454 276 456
rect 76 446 108 454
rect 126 446 138 454
rect 156 446 168 454
rect 186 446 198 454
rect 216 446 228 454
rect 236 446 276 454
rect 76 438 276 446
rect 76 400 276 432
rect 76 392 112 400
rect 240 392 276 400
rect 76 388 276 392
rect 76 380 112 388
rect 240 380 276 388
rect 76 348 276 380
rect 76 334 276 342
rect 76 326 110 334
rect 128 326 140 334
rect 158 326 170 334
rect 188 326 200 334
rect 218 326 230 334
rect 238 326 276 334
rect 76 322 276 326
rect 76 314 110 322
rect 128 314 140 322
rect 158 314 170 322
rect 188 314 200 322
rect 218 314 230 322
rect 238 314 276 322
rect 76 306 276 314
rect 76 268 276 300
rect 76 250 112 268
rect 240 250 276 268
rect 76 218 276 250
rect 76 204 276 212
rect 76 196 109 204
rect 127 196 139 204
rect 157 196 169 204
rect 187 196 199 204
rect 217 196 229 204
rect 237 196 276 204
rect 76 192 276 196
rect 76 184 109 192
rect 127 184 139 192
rect 157 184 169 192
rect 187 184 199 192
rect 217 184 229 192
rect 237 184 276 192
rect 76 176 276 184
rect 76 138 276 170
rect 76 120 112 138
rect 240 120 276 138
rect 76 88 276 120
rect 324 454 524 456
rect 324 446 364 454
rect 382 446 394 454
rect 412 446 424 454
rect 442 446 454 454
rect 472 446 484 454
rect 492 446 524 454
rect 324 438 524 446
rect 76 75 276 82
rect 76 67 78 75
rect 86 74 276 75
rect 86 67 107 74
rect 76 66 107 67
rect 115 66 118 74
rect 236 66 276 74
rect 76 64 276 66
rect 324 400 524 432
rect 324 392 360 400
rect 488 392 524 400
rect 324 388 524 392
rect 324 380 360 388
rect 488 380 524 388
rect 324 348 524 380
rect 324 335 524 342
rect 324 327 363 335
rect 381 327 393 335
rect 411 327 423 335
rect 441 327 453 335
rect 471 327 483 335
rect 491 327 524 335
rect 324 323 524 327
rect 324 315 363 323
rect 381 315 393 323
rect 411 315 423 323
rect 441 315 453 323
rect 471 315 483 323
rect 491 315 524 323
rect 324 306 524 315
rect 324 268 524 300
rect 324 250 360 268
rect 488 250 524 268
rect 324 218 524 250
rect 324 204 524 212
rect 324 196 364 204
rect 382 196 394 204
rect 412 196 424 204
rect 442 196 454 204
rect 472 196 484 204
rect 492 196 524 204
rect 324 192 524 196
rect 324 184 364 192
rect 382 184 394 192
rect 412 184 424 192
rect 442 184 454 192
rect 472 184 484 192
rect 492 184 524 192
rect 324 176 524 184
rect 324 138 524 170
rect 324 120 360 138
rect 488 120 524 138
rect 324 88 524 120
rect 324 74 524 82
rect 324 66 364 74
rect 492 66 524 74
rect 324 64 524 66
<< pdiffusion >>
rect 72 1270 280 1272
rect 72 1262 90 1270
rect 108 1262 112 1270
rect 120 1262 132 1270
rect 150 1262 162 1270
rect 180 1262 192 1270
rect 210 1262 222 1270
rect 230 1262 280 1270
rect 72 1260 280 1262
rect 76 1258 280 1260
rect 76 1254 276 1258
rect 76 1216 276 1248
rect 76 1198 112 1216
rect 240 1198 276 1216
rect 76 1166 276 1198
rect 76 1152 276 1160
rect 76 1144 123 1152
rect 141 1144 153 1152
rect 171 1144 183 1152
rect 201 1144 213 1152
rect 231 1144 276 1152
rect 76 1140 276 1144
rect 76 1132 123 1140
rect 141 1132 153 1140
rect 171 1132 183 1140
rect 201 1132 213 1140
rect 231 1132 276 1140
rect 76 1124 276 1132
rect 76 1087 276 1118
rect 76 1069 112 1087
rect 240 1069 276 1087
rect 76 1038 276 1069
rect 76 1024 276 1032
rect 76 1016 122 1024
rect 140 1016 152 1024
rect 170 1016 182 1024
rect 200 1016 212 1024
rect 230 1016 276 1024
rect 76 1012 276 1016
rect 76 1004 122 1012
rect 140 1004 152 1012
rect 170 1004 182 1012
rect 200 1004 212 1012
rect 230 1004 276 1012
rect 76 996 276 1004
rect 76 958 276 990
rect 76 940 112 958
rect 240 940 276 958
rect 76 908 276 940
rect 320 1270 528 1272
rect 320 1262 366 1270
rect 374 1262 386 1270
rect 404 1262 416 1270
rect 434 1262 446 1270
rect 464 1262 476 1270
rect 484 1262 488 1270
rect 506 1262 528 1270
rect 320 1260 528 1262
rect 320 1258 524 1260
rect 324 1254 524 1258
rect 76 894 276 902
rect 76 886 123 894
rect 141 886 153 894
rect 171 886 183 894
rect 201 886 213 894
rect 231 886 276 894
rect 76 884 276 886
rect 324 1216 524 1248
rect 324 1198 360 1216
rect 488 1198 524 1216
rect 324 1166 524 1198
rect 324 1152 524 1160
rect 324 1144 368 1152
rect 386 1144 398 1152
rect 416 1144 428 1152
rect 446 1144 458 1152
rect 476 1144 524 1152
rect 324 1140 524 1144
rect 324 1132 368 1140
rect 386 1132 398 1140
rect 416 1132 428 1140
rect 446 1132 458 1140
rect 476 1132 524 1140
rect 324 1124 524 1132
rect 324 1087 524 1118
rect 324 1069 360 1087
rect 488 1069 524 1087
rect 324 1038 524 1069
rect 324 1024 524 1032
rect 324 1016 367 1024
rect 385 1016 397 1024
rect 415 1016 427 1024
rect 445 1016 457 1024
rect 475 1016 524 1024
rect 324 1012 524 1016
rect 324 1004 367 1012
rect 385 1004 397 1012
rect 415 1004 427 1012
rect 445 1004 457 1012
rect 475 1004 524 1012
rect 324 996 524 1004
rect 324 958 524 990
rect 324 940 360 958
rect 488 940 524 958
rect 324 908 524 940
rect 324 894 524 902
rect 324 886 369 894
rect 387 886 399 894
rect 417 886 429 894
rect 447 886 459 894
rect 477 886 524 894
rect 324 884 524 886
rect 126 643 134 649
rect 158 643 166 649
rect 222 643 230 649
rect 384 643 394 649
rect 418 643 426 649
rect 450 643 456 649
rect 482 643 490 649
rect 514 643 522 649
rect 546 643 552 649
rect 578 643 586 649
rect 26 629 38 643
rect 26 541 28 629
rect 36 541 38 629
rect 26 539 38 541
rect 42 641 54 643
rect 42 633 44 641
rect 52 633 54 641
rect 42 621 54 633
rect 42 613 44 621
rect 52 613 54 621
rect 42 601 54 613
rect 42 593 44 601
rect 52 593 54 601
rect 42 581 54 593
rect 42 573 44 581
rect 52 573 54 581
rect 42 561 54 573
rect 42 553 44 561
rect 52 553 54 561
rect 42 539 54 553
rect 58 639 70 643
rect 58 541 60 639
rect 68 541 70 639
rect 58 539 70 541
rect 76 629 88 643
rect 76 541 78 629
rect 86 541 88 629
rect 76 539 88 541
rect 92 641 104 643
rect 92 633 94 641
rect 102 633 104 641
rect 92 621 104 633
rect 92 613 94 621
rect 102 613 104 621
rect 92 601 104 613
rect 92 593 94 601
rect 102 593 104 601
rect 92 581 104 593
rect 92 573 94 581
rect 102 573 104 581
rect 92 561 104 573
rect 92 553 94 561
rect 102 553 104 561
rect 92 539 104 553
rect 108 639 120 643
rect 108 541 110 639
rect 118 541 120 639
rect 108 539 120 541
rect 124 633 136 643
rect 124 625 126 633
rect 134 625 136 633
rect 124 613 136 625
rect 124 605 126 613
rect 134 605 136 613
rect 124 593 136 605
rect 124 585 126 593
rect 134 585 136 593
rect 124 573 136 585
rect 124 565 126 573
rect 134 565 136 573
rect 124 539 136 565
rect 140 639 152 643
rect 140 541 142 639
rect 150 541 152 639
rect 140 539 152 541
rect 156 633 168 643
rect 156 625 158 633
rect 166 625 168 633
rect 156 613 168 625
rect 156 605 158 613
rect 166 605 168 613
rect 156 583 168 605
rect 156 565 158 583
rect 166 565 168 583
rect 156 553 168 565
rect 156 545 158 553
rect 166 545 168 553
rect 156 539 168 545
rect 172 640 184 643
rect 172 542 174 640
rect 182 542 184 640
rect 172 539 184 542
rect 188 633 200 643
rect 188 625 190 633
rect 198 625 200 633
rect 188 613 200 625
rect 188 605 190 613
rect 198 605 200 613
rect 188 593 200 605
rect 188 585 190 593
rect 198 585 200 593
rect 188 573 200 585
rect 188 565 190 573
rect 198 565 200 573
rect 188 553 200 565
rect 188 545 190 553
rect 198 545 200 553
rect 188 539 200 545
rect 204 639 216 643
rect 204 541 206 639
rect 214 541 216 639
rect 204 539 216 541
rect 220 641 232 643
rect 220 633 222 641
rect 230 633 232 641
rect 220 621 232 633
rect 220 613 222 621
rect 230 613 232 621
rect 220 601 232 613
rect 220 593 222 601
rect 230 593 232 601
rect 220 581 232 593
rect 220 573 222 581
rect 230 573 232 581
rect 220 561 232 573
rect 220 553 222 561
rect 230 553 232 561
rect 220 539 232 553
rect 236 640 248 643
rect 236 542 238 640
rect 246 542 248 640
rect 236 539 248 542
rect 252 623 264 643
rect 252 545 254 623
rect 262 545 264 623
rect 252 539 264 545
rect 268 640 280 643
rect 268 632 270 640
rect 278 632 280 640
rect 268 614 280 632
rect 268 556 270 614
rect 278 556 280 614
rect 268 539 280 556
rect 284 641 296 643
rect 284 543 286 641
rect 294 543 296 641
rect 284 539 296 543
rect 300 619 312 643
rect 300 541 302 619
rect 310 541 312 619
rect 300 539 312 541
rect 384 633 396 643
rect 384 625 386 633
rect 394 625 396 633
rect 384 613 396 625
rect 384 605 386 613
rect 394 605 396 613
rect 384 583 396 605
rect 384 565 386 583
rect 394 565 396 583
rect 384 553 396 565
rect 384 545 386 553
rect 394 545 396 553
rect 384 539 396 545
rect 400 633 412 643
rect 400 545 402 633
rect 410 545 412 633
rect 400 539 412 545
rect 416 633 428 643
rect 416 625 418 633
rect 426 625 428 633
rect 416 613 428 625
rect 416 605 418 613
rect 426 605 428 613
rect 416 583 428 605
rect 416 565 418 583
rect 426 565 428 583
rect 416 553 428 565
rect 416 545 418 553
rect 426 545 428 553
rect 416 539 428 545
rect 432 633 444 643
rect 432 545 434 633
rect 442 545 444 633
rect 432 539 444 545
rect 448 633 460 643
rect 448 625 450 633
rect 458 625 460 633
rect 448 613 460 625
rect 448 605 450 613
rect 458 605 460 613
rect 448 583 460 605
rect 448 565 450 583
rect 458 565 460 583
rect 448 553 460 565
rect 448 545 450 553
rect 458 545 460 553
rect 448 539 460 545
rect 464 633 476 643
rect 464 545 466 633
rect 474 545 476 633
rect 464 539 476 545
rect 480 633 492 643
rect 480 625 482 633
rect 490 625 492 633
rect 480 613 492 625
rect 480 605 482 613
rect 490 605 492 613
rect 480 583 492 605
rect 480 565 482 583
rect 490 565 492 583
rect 480 553 492 565
rect 480 545 482 553
rect 490 545 492 553
rect 480 539 492 545
rect 496 633 508 643
rect 496 545 498 633
rect 506 545 508 633
rect 496 539 508 545
rect 512 633 524 643
rect 512 625 514 633
rect 522 625 524 633
rect 512 613 524 625
rect 512 605 514 613
rect 522 605 524 613
rect 512 583 524 605
rect 512 565 514 583
rect 522 565 524 583
rect 512 553 524 565
rect 512 545 514 553
rect 522 545 524 553
rect 512 539 524 545
rect 528 633 540 643
rect 528 545 530 633
rect 538 545 540 633
rect 528 539 540 545
rect 544 633 556 643
rect 544 625 546 633
rect 554 625 556 633
rect 544 613 556 625
rect 544 605 546 613
rect 554 605 556 613
rect 544 583 556 605
rect 544 565 546 583
rect 554 565 556 583
rect 544 553 556 565
rect 544 545 546 553
rect 554 545 556 553
rect 544 539 556 545
rect 560 633 572 643
rect 560 545 562 633
rect 570 545 572 633
rect 560 539 572 545
rect 576 633 586 643
rect 576 625 578 633
rect 576 613 586 625
rect 576 605 578 613
rect 576 593 586 605
rect 576 585 578 593
rect 576 573 586 585
rect 576 565 578 573
rect 576 553 586 565
rect 576 545 578 553
rect 576 539 586 545
rect 158 535 166 539
rect 384 535 394 539
rect 482 535 490 539
rect 578 535 586 539
<< ndcontact >>
rect 28 722 36 760
rect 44 752 52 760
rect 44 732 52 740
rect 44 712 52 720
rect 60 710 68 758
rect 78 721 86 759
rect 94 748 102 756
rect 94 728 102 736
rect 94 708 102 716
rect 110 711 118 759
rect 126 748 134 756
rect 126 728 134 736
rect 126 708 134 716
rect 142 711 150 759
rect 158 748 166 756
rect 158 728 166 736
rect 158 708 166 716
rect 174 711 182 759
rect 190 748 198 756
rect 190 728 198 736
rect 190 708 198 716
rect 206 712 214 760
rect 222 748 230 756
rect 222 728 230 736
rect 222 708 230 716
rect 238 730 246 758
rect 254 708 262 756
rect 270 730 278 758
rect 270 710 278 718
rect 286 755 294 763
rect 286 744 294 752
rect 286 732 294 740
rect 286 720 294 728
rect 302 756 310 764
rect 302 744 310 752
rect 302 733 310 741
rect 302 720 310 728
rect 302 708 310 716
rect 386 752 394 760
rect 386 732 394 740
rect 386 712 394 720
rect 402 712 410 760
rect 418 730 426 748
rect 418 709 426 717
rect 434 712 442 760
rect 450 753 458 761
rect 450 733 458 741
rect 450 713 458 721
rect 466 713 474 761
rect 482 753 490 761
rect 482 733 490 741
rect 482 713 490 721
rect 498 713 506 761
rect 514 753 522 761
rect 514 733 522 741
rect 514 713 522 721
rect 530 713 538 761
rect 546 753 554 761
rect 546 733 554 741
rect 546 713 554 721
rect 562 713 570 761
rect 578 753 586 761
rect 578 733 586 741
rect 578 713 586 721
rect 108 446 126 454
rect 138 446 156 454
rect 168 446 186 454
rect 198 446 216 454
rect 228 446 236 454
rect 112 392 240 400
rect 112 380 240 388
rect 110 326 128 334
rect 140 326 158 334
rect 170 326 188 334
rect 200 326 218 334
rect 230 326 238 334
rect 110 314 128 322
rect 140 314 158 322
rect 170 314 188 322
rect 200 314 218 322
rect 230 314 238 322
rect 112 250 240 268
rect 109 196 127 204
rect 139 196 157 204
rect 169 196 187 204
rect 199 196 217 204
rect 229 196 237 204
rect 109 184 127 192
rect 139 184 157 192
rect 169 184 187 192
rect 199 184 217 192
rect 229 184 237 192
rect 112 120 240 138
rect 364 446 382 454
rect 394 446 412 454
rect 424 446 442 454
rect 454 446 472 454
rect 484 446 492 454
rect 78 67 86 75
rect 107 66 115 74
rect 118 66 236 74
rect 360 392 488 400
rect 360 380 488 388
rect 363 327 381 335
rect 393 327 411 335
rect 423 327 441 335
rect 453 327 471 335
rect 483 327 491 335
rect 363 315 381 323
rect 393 315 411 323
rect 423 315 441 323
rect 453 315 471 323
rect 483 315 491 323
rect 360 250 488 268
rect 364 196 382 204
rect 394 196 412 204
rect 424 196 442 204
rect 454 196 472 204
rect 484 196 492 204
rect 364 184 382 192
rect 394 184 412 192
rect 424 184 442 192
rect 454 184 472 192
rect 484 184 492 192
rect 360 120 488 138
rect 364 66 492 74
<< pdcontact >>
rect 90 1262 108 1270
rect 112 1262 120 1270
rect 132 1262 150 1270
rect 162 1262 180 1270
rect 192 1262 210 1270
rect 222 1262 230 1270
rect 112 1198 240 1216
rect 123 1144 141 1152
rect 153 1144 171 1152
rect 183 1144 201 1152
rect 213 1144 231 1152
rect 123 1132 141 1140
rect 153 1132 171 1140
rect 183 1132 201 1140
rect 213 1132 231 1140
rect 112 1069 240 1087
rect 122 1016 140 1024
rect 152 1016 170 1024
rect 182 1016 200 1024
rect 212 1016 230 1024
rect 122 1004 140 1012
rect 152 1004 170 1012
rect 182 1004 200 1012
rect 212 1004 230 1012
rect 112 940 240 958
rect 366 1262 374 1270
rect 386 1262 404 1270
rect 416 1262 434 1270
rect 446 1262 464 1270
rect 476 1262 484 1270
rect 488 1262 506 1270
rect 123 886 141 894
rect 153 886 171 894
rect 183 886 201 894
rect 213 886 231 894
rect 360 1198 488 1216
rect 368 1144 386 1152
rect 398 1144 416 1152
rect 428 1144 446 1152
rect 458 1144 476 1152
rect 368 1132 386 1140
rect 398 1132 416 1140
rect 428 1132 446 1140
rect 458 1132 476 1140
rect 360 1069 488 1087
rect 367 1016 385 1024
rect 397 1016 415 1024
rect 427 1016 445 1024
rect 457 1016 475 1024
rect 367 1004 385 1012
rect 397 1004 415 1012
rect 427 1004 445 1012
rect 457 1004 475 1012
rect 360 940 488 958
rect 369 886 387 894
rect 399 886 417 894
rect 429 886 447 894
rect 459 886 477 894
rect 28 541 36 629
rect 44 633 52 641
rect 44 613 52 621
rect 44 593 52 601
rect 44 573 52 581
rect 44 553 52 561
rect 60 541 68 639
rect 78 541 86 629
rect 94 633 102 641
rect 94 613 102 621
rect 94 593 102 601
rect 94 573 102 581
rect 94 553 102 561
rect 110 541 118 639
rect 126 625 134 633
rect 126 605 134 613
rect 126 585 134 593
rect 126 565 134 573
rect 142 541 150 639
rect 158 625 166 633
rect 158 605 166 613
rect 158 565 166 583
rect 158 545 166 553
rect 174 542 182 640
rect 190 625 198 633
rect 190 605 198 613
rect 190 585 198 593
rect 190 565 198 573
rect 190 545 198 553
rect 206 541 214 639
rect 222 633 230 641
rect 222 613 230 621
rect 222 593 230 601
rect 222 573 230 581
rect 222 553 230 561
rect 238 542 246 640
rect 254 545 262 623
rect 270 632 278 640
rect 270 556 278 614
rect 286 543 294 641
rect 302 541 310 619
rect 386 625 394 633
rect 386 605 394 613
rect 386 565 394 583
rect 386 545 394 553
rect 402 545 410 633
rect 418 625 426 633
rect 418 605 426 613
rect 418 565 426 583
rect 418 545 426 553
rect 434 545 442 633
rect 450 625 458 633
rect 450 605 458 613
rect 450 565 458 583
rect 450 545 458 553
rect 466 545 474 633
rect 482 625 490 633
rect 482 605 490 613
rect 482 565 490 583
rect 482 545 490 553
rect 498 545 506 633
rect 514 625 522 633
rect 514 605 522 613
rect 514 565 522 583
rect 514 545 522 553
rect 530 545 538 633
rect 546 625 554 633
rect 546 605 554 613
rect 546 565 554 583
rect 546 545 554 553
rect 562 545 570 633
rect 578 625 586 633
rect 578 605 586 613
rect 578 585 586 593
rect 578 565 586 573
rect 578 545 586 553
<< psubstratepdiff >>
rect 0 1334 600 1340
rect 0 826 2 1334
rect 10 1314 14 1334
rect 232 1316 368 1334
rect 576 1332 600 1334
rect 576 1316 580 1332
rect 20 1314 580 1316
rect 20 840 22 1314
rect 234 840 294 842
rect 306 840 366 842
rect 578 840 580 1314
rect 20 839 580 840
rect 20 826 30 839
rect 0 821 30 826
rect 58 821 78 839
rect 226 821 296 839
rect 304 821 368 839
rect 576 824 580 839
rect 598 824 600 1332
rect 576 821 600 824
rect 0 820 600 821
rect 0 814 12 820
rect 0 686 2 814
rect 10 697 12 814
rect 586 813 600 820
rect 586 805 590 813
rect 598 805 600 813
rect 586 793 600 805
rect 586 785 590 793
rect 598 785 600 793
rect 586 773 600 785
rect 586 767 590 773
rect 582 765 590 767
rect 598 765 600 773
rect 582 761 600 765
rect 586 753 600 761
rect 586 745 590 753
rect 598 745 600 753
rect 586 733 600 745
rect 586 725 590 733
rect 598 725 600 733
rect 586 713 600 725
rect 10 690 14 697
rect 30 694 46 697
rect 30 690 34 694
rect 10 686 34 690
rect 42 690 46 694
rect 94 695 100 701
rect 62 693 100 695
rect 62 690 76 693
rect 42 686 76 690
rect 0 685 76 686
rect 84 685 90 693
rect 98 689 100 693
rect 126 695 134 701
rect 158 695 166 701
rect 126 693 168 695
rect 126 689 128 693
rect 98 685 128 689
rect 166 690 168 693
rect 222 697 230 701
rect 194 695 270 697
rect 194 690 198 695
rect 166 687 198 690
rect 206 687 216 695
rect 224 687 248 695
rect 256 690 270 695
rect 384 697 394 701
rect 418 697 426 701
rect 450 697 456 701
rect 296 694 456 697
rect 296 693 446 694
rect 296 690 388 693
rect 256 687 388 690
rect 166 685 388 687
rect 426 686 446 693
rect 454 691 456 694
rect 482 697 490 701
rect 514 697 522 701
rect 546 697 552 701
rect 482 693 552 697
rect 586 705 590 713
rect 598 705 600 713
rect 586 701 600 705
rect 578 693 600 701
rect 482 691 484 693
rect 454 686 484 691
rect 426 685 484 686
rect 502 685 514 693
rect 522 692 552 693
rect 522 685 542 692
rect 0 684 542 685
rect 550 691 552 692
rect 578 691 580 693
rect 550 685 580 691
rect 598 685 600 693
rect 550 684 600 685
rect 0 683 600 684
rect 28 486 562 492
rect 28 484 106 486
rect 28 456 34 484
rect 72 468 106 484
rect 234 478 364 486
rect 72 466 108 468
rect 52 460 108 466
rect 52 456 60 460
rect 28 444 60 456
rect 28 416 34 444
rect 52 416 60 444
rect 76 458 108 460
rect 126 458 138 468
rect 156 458 168 468
rect 186 458 198 468
rect 216 458 228 468
rect 234 466 296 478
rect 236 460 296 466
rect 304 460 364 478
rect 492 484 562 486
rect 236 458 276 460
rect 76 456 276 458
rect 286 448 314 460
rect 28 404 60 416
rect 28 376 34 404
rect 52 376 60 404
rect 28 364 60 376
rect 28 336 34 364
rect 52 336 60 364
rect 28 324 60 336
rect 28 296 34 324
rect 52 296 60 324
rect 28 284 60 296
rect 28 256 34 284
rect 52 256 60 284
rect 28 244 60 256
rect 28 216 34 244
rect 52 216 60 244
rect 28 204 60 216
rect 28 176 34 204
rect 52 176 60 204
rect 28 164 60 176
rect 28 136 34 164
rect 52 136 60 164
rect 28 124 60 136
rect 28 96 34 124
rect 52 96 60 124
rect 28 84 60 96
rect 28 66 34 84
rect 52 66 60 84
rect 286 430 296 448
rect 304 430 314 448
rect 324 458 364 460
rect 382 458 394 468
rect 412 458 424 468
rect 442 458 454 468
rect 472 458 484 468
rect 492 466 542 484
rect 560 466 562 484
rect 492 461 562 466
rect 492 460 542 461
rect 492 458 524 460
rect 324 456 524 458
rect 540 453 542 460
rect 560 453 562 461
rect 540 441 562 453
rect 286 418 314 430
rect 286 400 296 418
rect 304 400 314 418
rect 286 388 314 400
rect 286 370 296 388
rect 304 370 314 388
rect 286 358 314 370
rect 286 340 296 358
rect 304 340 314 358
rect 286 328 314 340
rect 286 310 296 328
rect 304 310 314 328
rect 286 288 314 310
rect 286 280 296 288
rect 304 280 314 288
rect 286 268 314 280
rect 286 250 296 268
rect 304 250 314 268
rect 286 238 314 250
rect 286 220 296 238
rect 304 220 314 238
rect 286 208 314 220
rect 286 190 296 208
rect 304 190 314 208
rect 286 178 314 190
rect 286 170 296 178
rect 304 170 314 178
rect 286 148 314 170
rect 286 130 296 148
rect 304 130 314 148
rect 286 118 314 130
rect 286 110 296 118
rect 304 110 314 118
rect 28 60 60 66
rect 76 60 78 64
rect 28 58 78 60
rect 28 50 34 58
rect 42 50 48 58
rect 86 56 107 64
rect 76 50 107 56
rect 28 44 107 50
rect 28 38 78 44
rect 28 30 48 38
rect 86 36 107 44
rect 115 62 276 64
rect 115 36 128 62
rect 76 34 128 36
rect 136 34 148 62
rect 156 34 168 62
rect 176 34 188 62
rect 196 34 208 62
rect 216 34 228 62
rect 236 60 276 62
rect 286 60 314 110
rect 540 413 542 441
rect 560 413 562 441
rect 540 401 562 413
rect 540 373 542 401
rect 560 373 562 401
rect 540 361 562 373
rect 540 333 542 361
rect 560 333 562 361
rect 540 321 562 333
rect 540 293 542 321
rect 560 293 562 321
rect 540 281 562 293
rect 540 253 542 281
rect 560 253 562 281
rect 540 241 562 253
rect 540 213 542 241
rect 560 213 562 241
rect 540 201 562 213
rect 540 173 542 201
rect 560 173 562 201
rect 540 161 562 173
rect 540 133 542 161
rect 560 133 562 161
rect 540 121 562 133
rect 540 93 542 121
rect 560 93 562 121
rect 324 62 484 64
rect 324 60 364 62
rect 236 34 364 60
rect 372 34 384 62
rect 392 34 404 62
rect 412 34 424 62
rect 432 34 444 62
rect 452 34 464 62
rect 472 36 484 62
rect 492 60 524 64
rect 540 81 562 93
rect 540 63 542 81
rect 560 63 562 81
rect 540 60 562 63
rect 492 58 562 60
rect 492 50 526 58
rect 544 50 552 58
rect 560 50 562 58
rect 492 40 562 50
rect 492 36 526 40
rect 472 34 526 36
rect 76 32 526 34
rect 534 38 562 40
rect 534 32 552 38
rect 76 30 552 32
rect 560 30 562 38
rect 28 28 562 30
<< nsubstratendiff >>
rect 38 1294 562 1296
rect 38 1290 296 1294
rect 38 1280 90 1290
rect 38 1252 40 1280
rect 58 1272 90 1280
rect 108 1272 112 1290
rect 120 1272 132 1290
rect 150 1272 162 1290
rect 180 1272 192 1290
rect 210 1272 222 1290
rect 230 1286 296 1290
rect 304 1290 562 1294
rect 304 1286 366 1290
rect 230 1274 366 1286
rect 230 1272 296 1274
rect 58 1260 72 1272
rect 58 1252 60 1260
rect 280 1258 296 1272
rect 38 1240 60 1252
rect 38 1212 40 1240
rect 58 1212 60 1240
rect 38 1200 60 1212
rect 38 1172 40 1200
rect 58 1172 60 1200
rect 38 1160 60 1172
rect 38 1132 40 1160
rect 58 1132 60 1160
rect 38 1120 60 1132
rect 38 1092 40 1120
rect 58 1092 60 1120
rect 38 1080 60 1092
rect 38 1052 40 1080
rect 58 1052 60 1080
rect 38 1040 60 1052
rect 38 1012 40 1040
rect 58 1012 60 1040
rect 38 1000 60 1012
rect 38 972 40 1000
rect 58 972 60 1000
rect 38 960 60 972
rect 38 932 40 960
rect 58 932 60 960
rect 38 920 60 932
rect 38 892 40 920
rect 58 892 60 920
rect 284 1246 296 1258
rect 304 1272 366 1274
rect 374 1272 386 1290
rect 404 1272 416 1290
rect 434 1272 446 1290
rect 464 1272 476 1290
rect 484 1272 488 1290
rect 506 1280 562 1290
rect 506 1272 542 1280
rect 304 1258 320 1272
rect 528 1260 542 1272
rect 304 1246 316 1258
rect 284 1234 316 1246
rect 284 1206 296 1234
rect 304 1206 316 1234
rect 284 1194 316 1206
rect 284 1166 296 1194
rect 304 1166 316 1194
rect 284 1154 316 1166
rect 284 1126 296 1154
rect 304 1126 316 1154
rect 284 1114 316 1126
rect 284 1086 296 1114
rect 304 1086 316 1114
rect 284 1074 316 1086
rect 284 1046 296 1074
rect 304 1046 316 1074
rect 284 1034 316 1046
rect 284 1006 296 1034
rect 304 1006 316 1034
rect 284 994 316 1006
rect 284 966 296 994
rect 304 966 316 994
rect 284 954 316 966
rect 284 926 296 954
rect 304 926 316 954
rect 284 914 316 926
rect 38 880 60 892
rect 76 882 276 884
rect 76 880 103 882
rect 38 862 40 880
rect 58 874 103 880
rect 111 874 123 882
rect 141 874 153 882
rect 171 874 183 882
rect 201 874 213 882
rect 231 880 276 882
rect 284 886 296 914
rect 304 886 316 914
rect 540 1252 542 1260
rect 560 1252 562 1280
rect 540 1240 562 1252
rect 540 1212 542 1240
rect 560 1212 562 1240
rect 540 1200 562 1212
rect 540 1172 542 1200
rect 560 1172 562 1200
rect 540 1160 562 1172
rect 540 1132 542 1160
rect 560 1132 562 1160
rect 540 1120 562 1132
rect 540 1092 542 1120
rect 560 1092 562 1120
rect 540 1080 562 1092
rect 540 1052 542 1080
rect 560 1052 562 1080
rect 540 1040 562 1052
rect 540 1012 542 1040
rect 560 1012 562 1040
rect 540 1000 562 1012
rect 540 972 542 1000
rect 560 972 562 1000
rect 540 960 562 972
rect 540 932 542 960
rect 560 932 562 960
rect 540 920 562 932
rect 284 880 316 886
rect 324 882 524 884
rect 324 880 369 882
rect 231 874 369 880
rect 387 874 399 882
rect 417 874 429 882
rect 447 874 459 882
rect 477 874 489 882
rect 497 880 524 882
rect 540 892 542 920
rect 560 892 562 920
rect 540 880 562 892
rect 497 874 542 880
rect 58 870 296 874
rect 58 862 93 870
rect 231 866 296 870
rect 304 870 542 874
rect 304 866 369 870
rect 231 862 369 866
rect 507 862 542 870
rect 560 862 562 880
rect 38 860 562 862
rect 0 664 600 665
rect 0 663 580 664
rect 0 662 34 663
rect 0 644 2 662
rect 10 659 34 662
rect 10 653 14 659
rect 10 644 12 653
rect 30 655 34 659
rect 42 659 76 663
rect 42 655 46 659
rect 30 653 46 655
rect 62 655 76 659
rect 84 655 90 663
rect 98 659 128 663
rect 98 655 100 659
rect 62 653 100 655
rect 0 632 12 644
rect 126 655 128 659
rect 136 655 148 663
rect 166 659 196 663
rect 166 655 168 659
rect 126 653 168 655
rect 126 649 134 653
rect 158 649 166 653
rect 194 655 196 659
rect 204 655 218 663
rect 226 659 274 663
rect 226 655 244 659
rect 194 653 244 655
rect 222 649 230 653
rect 270 655 274 659
rect 282 655 388 663
rect 406 655 418 663
rect 426 655 446 663
rect 454 659 484 663
rect 454 655 456 659
rect 270 653 456 655
rect 384 649 394 653
rect 418 649 426 653
rect 450 649 456 653
rect 482 655 484 659
rect 502 655 514 663
rect 522 655 542 663
rect 550 659 580 663
rect 550 655 552 659
rect 482 653 552 655
rect 482 649 490 653
rect 514 649 522 653
rect 546 649 552 653
rect 578 656 580 659
rect 578 649 590 656
rect 586 646 590 649
rect 598 646 600 664
rect 0 624 2 632
rect 10 624 12 632
rect 0 612 12 624
rect 0 604 2 612
rect 10 604 12 612
rect 0 592 12 604
rect 0 584 2 592
rect 10 584 12 592
rect 0 572 12 584
rect 0 564 2 572
rect 10 564 12 572
rect 0 552 12 564
rect 0 544 2 552
rect 10 544 12 552
rect 0 532 12 544
rect 586 634 600 646
rect 586 626 590 634
rect 598 626 600 634
rect 586 614 600 626
rect 586 606 590 614
rect 598 606 600 614
rect 586 594 600 606
rect 586 586 590 594
rect 598 586 600 594
rect 586 574 600 586
rect 586 566 590 574
rect 598 566 600 574
rect 586 554 600 566
rect 586 546 590 554
rect 598 546 600 554
rect 0 524 2 532
rect 10 524 12 532
rect 0 523 12 524
rect 72 523 86 531
rect 158 531 166 535
rect 384 531 394 535
rect 482 531 490 535
rect 586 535 600 546
rect 578 534 600 535
rect 578 531 590 534
rect 112 529 580 531
rect 112 526 386 529
rect 112 523 118 526
rect 0 518 118 523
rect 226 521 386 526
rect 394 521 482 529
rect 226 519 482 521
rect 490 521 580 529
rect 598 526 600 534
rect 490 519 527 521
rect 0 516 218 518
rect 0 512 34 516
rect 0 4 4 512
rect 12 508 34 512
rect 72 514 218 516
rect 226 516 480 519
rect 72 508 108 514
rect 226 508 389 516
rect 457 511 480 516
rect 508 513 527 519
rect 535 513 540 521
rect 588 513 600 526
rect 508 512 600 513
rect 508 511 590 512
rect 457 508 590 511
rect 12 506 108 508
rect 216 506 590 508
rect 12 504 590 506
rect 12 16 16 504
rect 578 502 590 504
rect 578 16 580 502
rect 12 12 580 16
rect 12 10 56 12
rect 74 10 116 12
rect 0 2 14 4
rect 42 2 46 10
rect 334 4 338 12
rect 476 10 538 12
rect 586 4 590 14
rect 598 4 600 512
rect 54 2 76 4
rect 114 2 478 4
rect 536 2 600 4
rect 0 0 600 2
<< psubstratepcontact >>
rect 2 1314 10 1334
rect 14 1316 232 1334
rect 368 1316 576 1334
rect 14 1314 20 1316
rect 2 826 20 1314
rect 30 821 58 839
rect 78 821 226 839
rect 296 821 304 839
rect 368 821 576 839
rect 580 824 598 1332
rect 2 686 10 814
rect 590 805 598 813
rect 590 785 598 793
rect 590 765 598 773
rect 590 745 598 753
rect 590 725 598 733
rect 34 686 42 694
rect 76 685 84 693
rect 90 685 98 693
rect 128 685 166 693
rect 198 687 206 695
rect 216 687 224 695
rect 248 687 256 695
rect 388 685 426 693
rect 446 686 454 694
rect 590 705 598 713
rect 484 685 502 693
rect 514 685 522 693
rect 542 684 550 692
rect 580 685 598 693
rect 34 466 72 484
rect 106 468 234 486
rect 34 456 52 466
rect 34 416 52 444
rect 108 458 126 468
rect 138 458 156 468
rect 168 458 186 468
rect 198 458 216 468
rect 228 466 234 468
rect 228 458 236 466
rect 296 460 304 478
rect 364 468 492 486
rect 34 376 52 404
rect 34 336 52 364
rect 34 296 52 324
rect 34 256 52 284
rect 34 216 52 244
rect 34 176 52 204
rect 34 136 52 164
rect 34 96 52 124
rect 34 66 52 84
rect 296 430 304 448
rect 364 458 382 468
rect 394 458 412 468
rect 424 458 442 468
rect 454 458 472 468
rect 484 458 492 468
rect 542 466 560 484
rect 542 453 560 461
rect 296 400 304 418
rect 296 370 304 388
rect 296 340 304 358
rect 296 310 304 328
rect 296 280 304 288
rect 296 250 304 268
rect 296 220 304 238
rect 296 190 304 208
rect 296 170 304 178
rect 296 130 304 148
rect 296 110 304 118
rect 78 58 86 64
rect 34 50 42 58
rect 48 56 86 58
rect 48 50 76 56
rect 78 38 86 44
rect 48 36 86 38
rect 107 36 115 64
rect 48 30 76 36
rect 128 34 136 62
rect 148 34 156 62
rect 168 34 176 62
rect 188 34 196 62
rect 208 34 216 62
rect 228 34 236 62
rect 542 413 560 441
rect 542 373 560 401
rect 542 333 560 361
rect 542 293 560 321
rect 542 253 560 281
rect 542 213 560 241
rect 542 173 560 201
rect 542 133 560 161
rect 542 93 560 121
rect 364 34 372 62
rect 384 34 392 62
rect 404 34 412 62
rect 424 34 432 62
rect 444 34 452 62
rect 464 34 472 62
rect 484 36 492 64
rect 542 63 560 81
rect 526 50 544 58
rect 552 50 560 58
rect 526 32 534 40
rect 552 30 560 38
<< nsubstratencontact >>
rect 40 1252 58 1280
rect 90 1272 108 1290
rect 112 1272 120 1290
rect 132 1272 150 1290
rect 162 1272 180 1290
rect 192 1272 210 1290
rect 222 1272 230 1290
rect 296 1286 304 1294
rect 40 1212 58 1240
rect 40 1172 58 1200
rect 40 1132 58 1160
rect 40 1092 58 1120
rect 40 1052 58 1080
rect 40 1012 58 1040
rect 40 972 58 1000
rect 40 932 58 960
rect 40 892 58 920
rect 296 1246 304 1274
rect 366 1272 374 1290
rect 386 1272 404 1290
rect 416 1272 434 1290
rect 446 1272 464 1290
rect 476 1272 484 1290
rect 488 1272 506 1290
rect 296 1206 304 1234
rect 296 1166 304 1194
rect 296 1126 304 1154
rect 296 1086 304 1114
rect 296 1046 304 1074
rect 296 1006 304 1034
rect 296 966 304 994
rect 296 926 304 954
rect 40 862 58 880
rect 103 874 111 882
rect 123 874 141 882
rect 153 874 171 882
rect 183 874 201 882
rect 213 874 231 882
rect 296 886 304 914
rect 542 1252 560 1280
rect 542 1212 560 1240
rect 542 1172 560 1200
rect 542 1132 560 1160
rect 542 1092 560 1120
rect 542 1052 560 1080
rect 542 1012 560 1040
rect 542 972 560 1000
rect 542 932 560 960
rect 369 874 387 882
rect 399 874 417 882
rect 429 874 447 882
rect 459 874 477 882
rect 489 874 497 882
rect 542 892 560 920
rect 93 862 231 870
rect 296 866 304 874
rect 369 862 507 870
rect 542 862 560 880
rect 2 644 10 662
rect 34 655 42 663
rect 76 655 84 663
rect 90 655 98 663
rect 128 655 136 663
rect 148 655 166 663
rect 196 655 204 663
rect 218 655 226 663
rect 274 655 282 663
rect 388 655 406 663
rect 418 655 426 663
rect 446 655 454 663
rect 484 655 502 663
rect 514 655 522 663
rect 542 655 550 663
rect 580 656 598 664
rect 590 646 598 656
rect 2 624 10 632
rect 2 604 10 612
rect 2 584 10 592
rect 2 564 10 572
rect 2 544 10 552
rect 590 626 598 634
rect 590 606 598 614
rect 590 586 598 594
rect 590 566 598 574
rect 590 546 598 554
rect 2 524 10 532
rect 590 531 598 534
rect 118 518 226 526
rect 386 521 394 529
rect 482 519 490 529
rect 580 526 598 531
rect 580 521 588 526
rect 4 10 12 512
rect 34 508 72 516
rect 218 514 226 518
rect 108 508 226 514
rect 389 508 457 516
rect 480 511 508 519
rect 527 513 535 521
rect 540 513 588 521
rect 108 506 216 508
rect 590 502 598 512
rect 580 14 598 502
rect 580 12 586 14
rect 56 10 74 12
rect 116 10 334 12
rect 4 4 42 10
rect 14 2 42 4
rect 46 4 334 10
rect 338 10 476 12
rect 538 10 586 12
rect 338 4 586 10
rect 590 4 598 14
rect 46 2 54 4
rect 76 2 114 4
rect 478 2 536 4
<< polysilicon >>
rect 62 1248 76 1254
rect 276 1248 282 1254
rect 62 1228 74 1248
rect 62 1190 64 1228
rect 72 1190 74 1228
rect 62 1166 74 1190
rect 278 1166 282 1248
rect 62 1160 76 1166
rect 276 1160 282 1166
rect 62 1124 74 1160
rect 278 1124 282 1160
rect 62 1118 76 1124
rect 276 1118 282 1124
rect 62 1098 74 1118
rect 62 1060 64 1098
rect 72 1060 74 1098
rect 62 1038 74 1060
rect 278 1038 282 1118
rect 62 1032 76 1038
rect 276 1032 282 1038
rect 62 996 74 1032
rect 278 996 282 1032
rect 62 990 76 996
rect 276 990 282 996
rect 62 962 74 990
rect 62 904 64 962
rect 72 908 74 962
rect 278 908 282 990
rect 72 904 76 908
rect 62 902 76 904
rect 276 902 282 908
rect 318 1248 324 1254
rect 524 1248 538 1254
rect 318 1166 322 1248
rect 526 1225 538 1248
rect 526 1187 528 1225
rect 536 1187 538 1225
rect 526 1166 538 1187
rect 318 1160 324 1166
rect 524 1160 538 1166
rect 318 1124 322 1160
rect 526 1124 538 1160
rect 318 1118 324 1124
rect 524 1118 538 1124
rect 318 1038 322 1118
rect 526 1098 538 1118
rect 526 1060 528 1098
rect 536 1060 538 1098
rect 526 1038 538 1060
rect 318 1032 324 1038
rect 524 1032 538 1038
rect 318 996 322 1032
rect 526 996 538 1032
rect 318 990 324 996
rect 524 990 538 996
rect 318 908 322 990
rect 526 968 538 990
rect 526 910 528 968
rect 536 910 538 968
rect 526 908 538 910
rect 318 902 324 908
rect 524 902 538 908
rect 222 809 580 810
rect 222 791 223 809
rect 251 799 551 809
rect 251 791 387 799
rect 222 790 387 791
rect 386 781 387 790
rect 415 791 551 799
rect 579 791 580 809
rect 415 790 580 791
rect 415 781 416 790
rect 386 780 416 781
rect 48 778 70 780
rect 48 770 50 778
rect 68 770 70 778
rect 38 766 42 770
rect 48 768 70 770
rect 88 768 156 772
rect 54 766 58 768
rect 88 766 92 768
rect 104 766 108 768
rect 120 766 124 768
rect 136 766 140 768
rect 152 766 156 768
rect 168 768 236 772
rect 168 766 172 768
rect 184 766 188 768
rect 200 766 204 768
rect 216 766 220 768
rect 232 766 236 768
rect 248 766 252 770
rect 264 766 268 770
rect 280 766 284 770
rect 296 766 300 770
rect 396 767 400 780
rect 412 770 432 774
rect 412 767 416 770
rect 428 767 432 770
rect 444 769 464 773
rect 444 767 448 769
rect 460 767 464 769
rect 476 767 480 771
rect 492 767 496 771
rect 508 769 528 773
rect 508 767 512 769
rect 524 767 528 769
rect 540 769 560 773
rect 540 767 544 769
rect 556 767 560 769
rect 572 767 576 772
rect 38 704 42 706
rect 54 704 58 706
rect 16 702 42 704
rect 16 694 18 702
rect 26 700 42 702
rect 48 702 60 704
rect 26 694 28 700
rect 16 692 28 694
rect 48 694 50 702
rect 58 694 60 702
rect 88 700 92 706
rect 104 703 108 706
rect 120 703 124 706
rect 48 692 60 694
rect 102 701 124 703
rect 102 693 104 701
rect 122 693 124 701
rect 102 691 124 693
rect 136 701 140 706
rect 152 701 156 706
rect 168 704 172 706
rect 184 704 188 706
rect 168 702 192 704
rect 168 699 172 702
rect 170 694 172 699
rect 190 694 192 702
rect 200 701 204 706
rect 216 701 220 706
rect 232 701 236 706
rect 248 704 252 706
rect 264 704 268 706
rect 280 704 284 706
rect 296 704 300 706
rect 248 702 300 704
rect 248 700 274 702
rect 170 692 192 694
rect 272 694 274 700
rect 292 700 300 702
rect 396 705 400 707
rect 412 705 416 707
rect 396 701 416 705
rect 428 705 432 707
rect 444 705 448 707
rect 428 701 448 705
rect 460 705 464 707
rect 476 705 480 707
rect 292 694 294 700
rect 272 692 294 694
rect 458 703 480 705
rect 458 695 460 703
rect 478 695 480 703
rect 458 693 480 695
rect 492 705 496 707
rect 508 705 512 707
rect 492 701 512 705
rect 524 705 528 707
rect 540 705 544 707
rect 524 701 544 705
rect 556 705 560 707
rect 572 705 576 707
rect 554 703 576 705
rect 554 695 556 703
rect 574 695 576 703
rect 554 693 576 695
rect 62 678 294 680
rect 62 670 64 678
rect 82 670 160 678
rect 178 670 274 678
rect 292 670 294 678
rect 62 668 294 670
rect 16 655 28 657
rect 16 647 18 655
rect 26 649 28 655
rect 48 655 60 657
rect 26 647 42 649
rect 16 645 42 647
rect 48 647 50 655
rect 58 647 60 655
rect 102 655 124 657
rect 102 647 104 655
rect 122 647 124 655
rect 48 645 60 647
rect 38 643 42 645
rect 54 643 58 645
rect 88 643 92 647
rect 102 645 124 647
rect 104 643 108 645
rect 120 643 124 645
rect 170 655 192 657
rect 170 649 172 655
rect 136 643 140 647
rect 152 643 156 647
rect 168 647 172 649
rect 190 647 192 655
rect 246 655 268 657
rect 168 645 192 647
rect 168 643 172 645
rect 184 643 188 645
rect 200 643 204 647
rect 216 643 220 647
rect 246 647 248 655
rect 266 649 268 655
rect 266 647 300 649
rect 232 643 236 647
rect 246 645 300 647
rect 248 643 252 645
rect 264 643 268 645
rect 280 643 284 645
rect 296 643 300 645
rect 396 647 416 651
rect 396 643 400 647
rect 412 643 416 647
rect 428 647 448 651
rect 428 643 432 647
rect 444 643 448 647
rect 458 655 480 657
rect 458 647 460 655
rect 478 647 480 655
rect 458 645 480 647
rect 460 643 464 645
rect 476 643 480 645
rect 492 645 512 649
rect 492 643 496 645
rect 508 643 512 645
rect 524 645 544 649
rect 524 643 528 645
rect 540 643 544 645
rect 554 655 576 657
rect 554 647 556 655
rect 574 647 576 655
rect 554 645 576 647
rect 556 643 560 645
rect 572 643 576 645
rect 38 537 42 539
rect 54 537 58 539
rect 88 537 92 539
rect 104 537 108 539
rect 120 537 124 539
rect 136 537 140 539
rect 152 537 156 539
rect 20 535 42 537
rect 20 527 22 535
rect 40 527 42 535
rect 20 525 42 527
rect 48 535 70 537
rect 48 527 50 535
rect 68 527 70 535
rect 88 535 156 537
rect 48 525 70 527
rect 88 527 90 535
rect 108 533 156 535
rect 108 527 110 533
rect 168 537 172 539
rect 184 537 188 539
rect 200 537 204 539
rect 216 537 220 539
rect 232 537 236 539
rect 168 533 236 537
rect 248 535 252 539
rect 264 535 268 539
rect 280 535 284 539
rect 296 535 300 539
rect 396 535 400 539
rect 412 537 416 539
rect 428 537 432 539
rect 412 533 432 537
rect 444 537 448 539
rect 460 537 464 539
rect 444 533 464 537
rect 476 535 480 539
rect 492 535 496 539
rect 508 537 512 539
rect 524 537 528 539
rect 508 533 528 537
rect 540 537 544 539
rect 556 537 560 539
rect 540 533 560 537
rect 572 535 576 539
rect 88 525 110 527
rect 62 434 76 438
rect 62 86 64 434
rect 72 432 76 434
rect 276 432 284 438
rect 72 348 74 432
rect 278 348 284 432
rect 72 342 76 348
rect 276 342 284 348
rect 72 306 74 342
rect 278 306 284 342
rect 72 300 76 306
rect 276 300 284 306
rect 72 218 74 300
rect 278 218 284 300
rect 72 212 76 218
rect 276 212 284 218
rect 72 176 74 212
rect 278 176 284 212
rect 72 170 76 176
rect 276 170 284 176
rect 72 88 74 170
rect 278 88 284 170
rect 72 86 76 88
rect 62 82 76 86
rect 276 82 284 88
rect 316 432 324 438
rect 524 434 538 438
rect 524 432 528 434
rect 316 348 322 432
rect 526 348 528 432
rect 316 342 324 348
rect 524 342 528 348
rect 316 306 322 342
rect 526 306 528 342
rect 316 300 324 306
rect 524 300 528 306
rect 316 218 322 300
rect 526 218 528 300
rect 316 212 324 218
rect 524 212 528 218
rect 316 176 322 212
rect 526 176 528 212
rect 316 170 324 176
rect 524 170 528 176
rect 316 88 322 170
rect 526 88 528 170
rect 316 82 324 88
rect 524 86 528 88
rect 536 86 538 434
rect 524 82 538 86
<< polycontact >>
rect 64 1190 72 1228
rect 64 1060 72 1098
rect 64 904 72 962
rect 528 1187 536 1225
rect 528 1060 536 1098
rect 528 910 536 968
rect 223 791 251 809
rect 387 781 415 799
rect 551 791 579 809
rect 50 770 68 778
rect 18 694 26 702
rect 50 694 58 702
rect 104 693 122 701
rect 172 694 190 702
rect 274 694 292 702
rect 460 695 478 703
rect 556 695 574 703
rect 64 670 82 678
rect 160 670 178 678
rect 274 670 292 678
rect 18 647 26 655
rect 50 647 58 655
rect 104 647 122 655
rect 172 647 190 655
rect 248 647 266 655
rect 460 647 478 655
rect 556 647 574 655
rect 22 527 40 535
rect 50 527 68 535
rect 90 527 108 535
rect 64 86 72 434
rect 528 86 536 434
<< metal1 >>
rect 124 1400 476 1480
rect 204 1380 396 1400
rect 224 1360 376 1380
rect 0 1334 232 1338
rect 0 826 2 1334
rect 10 1314 14 1334
rect 28 1308 234 1310
rect 226 1300 234 1308
rect 36 1290 234 1300
rect 36 1282 40 1290
rect 36 1280 60 1282
rect 36 1252 40 1280
rect 58 1262 60 1280
rect 88 1272 90 1290
rect 108 1272 112 1290
rect 120 1272 122 1290
rect 88 1270 122 1272
rect 88 1262 90 1270
rect 108 1262 112 1270
rect 120 1262 122 1270
rect 130 1272 132 1290
rect 150 1272 152 1290
rect 130 1270 152 1272
rect 130 1262 132 1270
rect 150 1262 152 1270
rect 160 1272 162 1290
rect 180 1272 182 1290
rect 160 1270 182 1272
rect 160 1262 162 1270
rect 180 1262 182 1270
rect 190 1272 192 1290
rect 210 1272 212 1290
rect 190 1270 212 1272
rect 190 1262 192 1270
rect 210 1262 212 1270
rect 220 1272 222 1290
rect 230 1272 234 1290
rect 220 1270 234 1272
rect 220 1262 222 1270
rect 230 1262 234 1270
rect 58 1252 234 1262
rect 36 1251 234 1252
rect 36 1250 64 1251
rect 36 1242 40 1250
rect 58 1243 64 1250
rect 72 1244 234 1251
rect 72 1243 84 1244
rect 58 1242 84 1243
rect 36 1240 84 1242
rect 36 1212 40 1240
rect 58 1236 84 1240
rect 232 1236 234 1244
rect 58 1234 234 1236
rect 240 1308 360 1360
rect 368 1334 600 1338
rect 576 1332 600 1334
rect 576 1316 580 1332
rect 78 1233 104 1234
rect 36 1210 58 1212
rect 36 1202 40 1210
rect 36 1200 58 1202
rect 36 1172 40 1200
rect 78 1185 82 1233
rect 100 1185 104 1233
rect 240 1224 286 1308
rect 112 1216 286 1224
rect 240 1198 286 1216
rect 112 1191 286 1198
rect 78 1184 104 1185
rect 58 1180 234 1184
rect 58 1179 84 1180
rect 58 1172 64 1179
rect 36 1170 64 1172
rect 36 1162 40 1170
rect 58 1162 64 1170
rect 36 1160 64 1162
rect 36 1132 40 1160
rect 58 1132 64 1160
rect 36 1130 64 1132
rect 36 1122 40 1130
rect 58 1122 64 1130
rect 36 1120 64 1122
rect 36 1092 40 1120
rect 58 1111 64 1120
rect 72 1172 84 1179
rect 232 1172 234 1180
rect 72 1152 234 1172
rect 72 1144 83 1152
rect 121 1144 123 1152
rect 141 1144 143 1152
rect 151 1144 153 1152
rect 171 1144 173 1152
rect 181 1144 183 1152
rect 201 1144 203 1152
rect 211 1144 213 1152
rect 231 1144 234 1152
rect 72 1140 234 1144
rect 72 1132 83 1140
rect 121 1132 123 1140
rect 141 1132 143 1140
rect 151 1132 153 1140
rect 171 1132 173 1140
rect 181 1132 183 1140
rect 201 1132 203 1140
rect 211 1132 213 1140
rect 231 1132 234 1140
rect 72 1113 234 1132
rect 72 1111 84 1113
rect 58 1104 84 1111
rect 232 1105 234 1113
rect 36 1090 58 1092
rect 36 1082 40 1090
rect 36 1080 58 1082
rect 36 1052 40 1080
rect 78 1055 84 1104
rect 102 1104 234 1105
rect 102 1055 104 1104
rect 240 1096 286 1191
rect 111 1087 286 1096
rect 111 1069 112 1087
rect 240 1069 286 1087
rect 111 1061 286 1069
rect 78 1054 104 1055
rect 58 1052 234 1054
rect 36 1050 84 1052
rect 36 1042 40 1050
rect 58 1049 84 1050
rect 58 1042 64 1049
rect 36 1040 64 1042
rect 36 1012 40 1040
rect 58 1012 64 1040
rect 36 1010 64 1012
rect 36 1002 40 1010
rect 58 1002 64 1010
rect 36 1000 64 1002
rect 36 972 40 1000
rect 58 981 64 1000
rect 72 1044 84 1049
rect 232 1044 234 1052
rect 72 1024 234 1044
rect 72 1016 82 1024
rect 120 1016 122 1024
rect 140 1016 142 1024
rect 150 1016 152 1024
rect 170 1016 172 1024
rect 180 1016 182 1024
rect 200 1016 202 1024
rect 210 1016 212 1024
rect 230 1016 234 1024
rect 72 1012 234 1016
rect 72 1004 82 1012
rect 120 1004 122 1012
rect 140 1004 142 1012
rect 150 1004 152 1012
rect 170 1004 172 1012
rect 180 1004 182 1012
rect 200 1004 202 1012
rect 210 1004 212 1012
rect 230 1004 234 1012
rect 72 986 234 1004
rect 72 981 84 986
rect 58 978 84 981
rect 232 978 234 986
rect 58 976 234 978
rect 36 970 58 972
rect 36 962 40 970
rect 78 975 104 976
rect 36 960 58 962
rect 36 932 40 960
rect 36 930 58 932
rect 36 922 40 930
rect 36 920 58 922
rect 36 892 40 920
rect 36 890 58 892
rect 36 882 40 890
rect 36 880 58 882
rect 28 862 40 880
rect 28 860 58 862
rect 64 962 72 963
rect 64 872 72 904
rect 78 927 84 975
rect 102 927 104 975
rect 240 966 286 1061
rect 111 958 286 966
rect 111 940 112 958
rect 240 940 286 958
rect 111 933 286 940
rect 78 924 104 927
rect 78 922 232 924
rect 78 914 82 922
rect 230 914 232 922
rect 78 894 232 914
rect 78 886 80 894
rect 88 886 91 894
rect 99 886 102 894
rect 110 886 113 894
rect 121 886 123 894
rect 141 886 143 894
rect 151 886 153 894
rect 171 886 173 894
rect 181 886 183 894
rect 201 886 203 894
rect 211 886 213 894
rect 231 886 232 894
rect 78 882 232 886
rect 78 878 93 882
rect 88 874 93 878
rect 101 874 103 882
rect 111 874 113 882
rect 121 874 123 882
rect 141 874 143 882
rect 151 874 153 882
rect 171 874 173 882
rect 181 874 183 882
rect 201 874 203 882
rect 211 874 213 882
rect 231 874 232 882
rect 64 870 82 872
rect 64 860 82 862
rect 88 870 232 874
rect 88 862 93 870
rect 231 862 232 870
rect 88 860 232 862
rect 20 842 30 850
rect 20 839 58 842
rect 20 826 30 839
rect 0 821 30 826
rect 0 818 58 821
rect 0 814 14 818
rect 0 686 2 814
rect 10 790 14 814
rect 22 810 26 818
rect 54 810 58 818
rect 22 808 58 810
rect 10 786 22 790
rect 64 796 72 860
rect 226 842 231 850
rect 78 839 231 842
rect 226 821 231 839
rect 78 820 231 821
rect 78 818 216 820
rect 240 814 286 933
rect 294 1294 306 1296
rect 294 1286 296 1294
rect 304 1286 306 1294
rect 294 1284 306 1286
rect 294 1276 296 1284
rect 304 1276 306 1284
rect 294 1274 306 1276
rect 294 1246 296 1274
rect 304 1246 306 1274
rect 294 1244 306 1246
rect 294 1236 296 1244
rect 304 1236 306 1244
rect 294 1234 306 1236
rect 294 1206 296 1234
rect 304 1206 306 1234
rect 294 1204 306 1206
rect 294 1196 296 1204
rect 304 1196 306 1204
rect 294 1194 306 1196
rect 294 1166 296 1194
rect 304 1166 306 1194
rect 294 1164 306 1166
rect 294 1156 296 1164
rect 304 1156 306 1164
rect 294 1154 306 1156
rect 294 1126 296 1154
rect 304 1126 306 1154
rect 294 1124 306 1126
rect 294 1116 296 1124
rect 304 1116 306 1124
rect 294 1114 306 1116
rect 294 1086 296 1114
rect 304 1086 306 1114
rect 294 1084 306 1086
rect 294 1076 296 1084
rect 304 1076 306 1084
rect 294 1074 306 1076
rect 294 1046 296 1074
rect 304 1046 306 1074
rect 294 1044 306 1046
rect 294 1036 296 1044
rect 304 1036 306 1044
rect 294 1034 306 1036
rect 294 1006 296 1034
rect 304 1006 306 1034
rect 294 1004 306 1006
rect 294 996 296 1004
rect 304 996 306 1004
rect 294 994 306 996
rect 294 966 296 994
rect 304 966 306 994
rect 294 964 306 966
rect 294 956 296 964
rect 304 956 306 964
rect 294 954 306 956
rect 294 926 296 954
rect 304 926 306 954
rect 294 924 306 926
rect 294 916 296 924
rect 304 916 306 924
rect 294 914 306 916
rect 294 886 296 914
rect 304 886 306 914
rect 294 884 306 886
rect 294 876 296 884
rect 304 876 306 884
rect 294 874 306 876
rect 294 866 296 874
rect 304 866 306 874
rect 294 860 306 866
rect 314 1224 360 1308
rect 366 1302 374 1310
rect 366 1290 564 1302
rect 374 1272 376 1290
rect 366 1270 376 1272
rect 374 1262 376 1270
rect 384 1272 386 1290
rect 404 1272 406 1290
rect 384 1270 406 1272
rect 384 1262 386 1270
rect 404 1262 406 1270
rect 414 1272 416 1290
rect 434 1272 436 1290
rect 414 1270 436 1272
rect 414 1262 416 1270
rect 434 1262 436 1270
rect 444 1272 446 1290
rect 464 1272 466 1290
rect 444 1270 466 1272
rect 444 1262 446 1270
rect 464 1262 466 1270
rect 474 1272 476 1290
rect 484 1272 488 1290
rect 506 1272 508 1290
rect 474 1270 508 1272
rect 474 1262 476 1270
rect 484 1262 488 1270
rect 506 1262 508 1270
rect 536 1282 542 1290
rect 560 1282 564 1290
rect 536 1280 564 1282
rect 536 1262 542 1280
rect 366 1252 542 1262
rect 560 1252 564 1280
rect 366 1250 564 1252
rect 366 1244 528 1250
rect 366 1236 368 1244
rect 516 1242 528 1244
rect 536 1242 542 1250
rect 560 1242 564 1250
rect 516 1240 564 1242
rect 516 1236 542 1240
rect 366 1232 542 1236
rect 497 1229 522 1232
rect 314 1216 489 1224
rect 314 1198 360 1216
rect 488 1198 489 1216
rect 314 1191 489 1198
rect 314 1096 360 1191
rect 497 1181 498 1229
rect 516 1181 522 1229
rect 560 1212 564 1240
rect 542 1210 564 1212
rect 560 1202 564 1210
rect 542 1200 564 1202
rect 366 1178 542 1181
rect 366 1170 368 1178
rect 516 1176 542 1178
rect 516 1170 528 1176
rect 366 1152 528 1170
rect 366 1144 368 1152
rect 386 1144 388 1152
rect 396 1144 398 1152
rect 416 1144 418 1152
rect 426 1144 428 1152
rect 446 1144 448 1152
rect 456 1144 458 1152
rect 476 1144 478 1152
rect 516 1144 528 1152
rect 366 1140 528 1144
rect 366 1132 368 1140
rect 386 1132 388 1140
rect 396 1132 398 1140
rect 416 1132 418 1140
rect 426 1132 428 1140
rect 446 1132 448 1140
rect 456 1132 458 1140
rect 476 1132 478 1140
rect 516 1132 528 1140
rect 366 1114 528 1132
rect 366 1106 368 1114
rect 516 1108 528 1114
rect 536 1172 542 1176
rect 560 1172 564 1200
rect 536 1170 564 1172
rect 536 1162 542 1170
rect 560 1162 564 1170
rect 536 1160 564 1162
rect 536 1132 542 1160
rect 560 1132 564 1160
rect 536 1130 564 1132
rect 536 1122 542 1130
rect 560 1122 564 1130
rect 536 1120 564 1122
rect 536 1108 542 1120
rect 516 1106 542 1108
rect 366 1104 542 1106
rect 497 1103 522 1104
rect 314 1087 489 1096
rect 314 1069 360 1087
rect 488 1069 489 1087
rect 314 1061 489 1069
rect 314 966 360 1061
rect 497 1055 498 1103
rect 516 1055 522 1103
rect 560 1092 564 1120
rect 542 1090 564 1092
rect 560 1082 564 1090
rect 542 1080 564 1082
rect 497 1054 522 1055
rect 366 1052 542 1054
rect 560 1052 564 1080
rect 366 1044 368 1052
rect 516 1050 564 1052
rect 516 1049 542 1050
rect 516 1044 528 1049
rect 366 1024 528 1044
rect 366 1016 367 1024
rect 385 1016 387 1024
rect 395 1016 397 1024
rect 415 1016 417 1024
rect 425 1016 427 1024
rect 445 1016 447 1024
rect 455 1016 457 1024
rect 475 1016 477 1024
rect 515 1016 528 1024
rect 366 1012 528 1016
rect 366 1004 367 1012
rect 385 1004 387 1012
rect 395 1004 397 1012
rect 415 1004 417 1012
rect 425 1004 427 1012
rect 445 1004 447 1012
rect 455 1004 457 1012
rect 475 1004 477 1012
rect 515 1004 528 1012
rect 366 986 528 1004
rect 366 978 368 986
rect 516 981 528 986
rect 536 1042 542 1049
rect 560 1042 564 1050
rect 536 1040 564 1042
rect 536 1012 542 1040
rect 560 1012 564 1040
rect 536 1010 564 1012
rect 536 1002 542 1010
rect 560 1002 564 1010
rect 536 1000 564 1002
rect 536 981 542 1000
rect 516 978 542 981
rect 366 976 542 978
rect 497 974 522 976
rect 314 958 489 966
rect 314 940 360 958
rect 488 940 489 958
rect 314 933 489 940
rect 296 839 304 842
rect 296 820 304 821
rect 314 814 360 933
rect 497 926 500 974
rect 518 926 522 974
rect 560 972 564 1000
rect 542 970 564 972
rect 497 924 522 926
rect 368 922 522 924
rect 368 914 370 922
rect 518 914 522 922
rect 368 894 522 914
rect 368 886 369 894
rect 387 886 389 894
rect 397 886 399 894
rect 417 886 419 894
rect 427 886 429 894
rect 447 886 449 894
rect 457 886 459 894
rect 477 886 479 894
rect 487 886 490 894
rect 498 886 501 894
rect 509 886 512 894
rect 520 886 522 894
rect 368 882 522 886
rect 368 874 369 882
rect 387 874 389 882
rect 397 874 399 882
rect 417 874 419 882
rect 427 874 429 882
rect 447 874 449 882
rect 457 874 459 882
rect 477 874 479 882
rect 487 874 489 882
rect 497 874 499 882
rect 507 878 522 882
rect 507 874 512 878
rect 368 870 512 874
rect 528 872 536 910
rect 368 862 369 870
rect 507 862 512 870
rect 368 860 512 862
rect 518 870 536 872
rect 518 860 536 862
rect 560 962 564 970
rect 542 960 564 962
rect 560 932 564 960
rect 542 930 564 932
rect 560 922 564 930
rect 542 920 564 922
rect 560 892 564 920
rect 542 890 564 892
rect 560 882 564 890
rect 542 880 572 882
rect 560 862 572 880
rect 542 860 572 862
rect 576 842 580 850
rect 368 839 580 842
rect 576 824 580 839
rect 598 824 600 1332
rect 576 823 600 824
rect 576 821 590 823
rect 368 820 590 821
rect 586 815 590 820
rect 598 815 600 823
rect 78 808 216 810
rect 222 809 580 814
rect 64 787 83 796
rect 10 708 14 786
rect 74 780 83 787
rect 222 791 223 809
rect 251 806 551 809
rect 251 791 380 806
rect 222 786 380 791
rect 28 770 50 778
rect 74 774 262 780
rect 268 776 380 786
rect 386 799 416 800
rect 386 781 387 799
rect 415 781 416 799
rect 386 780 416 781
rect 422 791 551 806
rect 579 791 580 809
rect 422 790 580 791
rect 586 813 600 815
rect 586 805 590 813
rect 598 805 600 813
rect 586 803 600 805
rect 586 795 590 803
rect 598 795 600 803
rect 586 793 600 795
rect 422 780 457 790
rect 586 785 590 793
rect 598 785 600 793
rect 586 784 600 785
rect 254 770 262 774
rect 300 774 380 776
rect 422 774 430 780
rect 584 783 600 784
rect 584 776 590 783
rect 300 770 430 774
rect 578 775 590 776
rect 598 775 600 783
rect 578 773 600 775
rect 28 760 36 770
rect 28 720 36 722
rect 44 760 52 764
rect 44 750 52 752
rect 44 740 52 742
rect 44 730 52 732
rect 44 720 52 722
rect 38 712 44 714
rect 38 708 52 712
rect 60 758 68 764
rect 78 762 246 768
rect 78 759 86 762
rect 110 759 118 762
rect 94 746 102 748
rect 94 736 102 738
rect 94 726 102 728
rect 94 716 102 718
rect 68 710 70 716
rect 60 708 70 710
rect 10 686 12 708
rect 0 683 12 686
rect 38 696 44 708
rect 32 694 44 696
rect 0 662 12 665
rect 0 644 2 662
rect 10 644 12 662
rect 18 655 24 694
rect 32 686 34 694
rect 42 686 44 694
rect 32 684 44 686
rect 50 678 56 694
rect 64 678 70 708
rect 76 708 94 714
rect 142 759 150 762
rect 126 746 134 748
rect 126 736 134 738
rect 126 726 134 728
rect 126 716 134 718
rect 174 759 182 762
rect 158 746 166 748
rect 158 736 166 738
rect 158 726 166 728
rect 158 716 166 718
rect 76 693 98 708
rect 128 704 134 708
rect 206 760 214 762
rect 190 746 198 748
rect 190 736 198 738
rect 190 726 198 728
rect 190 716 198 718
rect 238 758 246 762
rect 206 708 214 712
rect 222 746 230 748
rect 222 736 230 738
rect 222 726 230 728
rect 238 728 246 730
rect 254 764 294 770
rect 316 766 430 770
rect 436 767 474 773
rect 254 756 262 764
rect 286 763 294 764
rect 222 716 230 718
rect 158 704 166 708
rect 128 693 166 704
rect 222 697 230 708
rect 84 685 90 693
rect 32 663 44 664
rect 32 655 34 663
rect 42 655 44 663
rect 32 653 44 655
rect 0 642 12 644
rect 0 634 2 642
rect 10 640 12 642
rect 10 636 22 640
rect 10 634 14 636
rect 0 632 14 634
rect 0 624 2 632
rect 10 624 14 632
rect 0 622 14 624
rect 0 614 2 622
rect 10 614 14 622
rect 0 612 14 614
rect 0 604 2 612
rect 10 604 14 612
rect 0 602 14 604
rect 0 594 2 602
rect 10 594 14 602
rect 0 592 14 594
rect 0 584 2 592
rect 10 584 14 592
rect 0 582 14 584
rect 0 574 2 582
rect 10 574 14 582
rect 0 572 14 574
rect 0 564 2 572
rect 10 564 14 572
rect 0 562 14 564
rect 0 554 2 562
rect 10 554 14 562
rect 0 552 14 554
rect 0 544 2 552
rect 10 548 14 552
rect 38 635 44 653
rect 50 655 56 670
rect 64 641 70 670
rect 44 631 52 633
rect 10 544 22 548
rect 0 542 16 544
rect 0 534 2 542
rect 10 534 16 542
rect 44 621 52 623
rect 44 611 52 613
rect 44 601 52 603
rect 44 591 52 593
rect 44 581 52 583
rect 44 571 52 573
rect 44 561 52 563
rect 60 639 70 641
rect 36 541 54 547
rect 68 632 70 639
rect 84 655 90 663
rect 106 655 112 693
rect 184 678 190 694
rect 196 695 230 697
rect 196 687 198 695
rect 214 687 216 695
rect 224 687 230 695
rect 196 684 230 687
rect 236 708 254 714
rect 270 728 278 730
rect 286 752 294 755
rect 286 740 294 744
rect 286 728 294 732
rect 302 752 310 756
rect 302 741 310 744
rect 302 728 310 733
rect 270 718 278 720
rect 302 716 310 720
rect 278 710 302 714
rect 270 708 302 710
rect 128 663 166 664
rect 136 655 138 663
rect 146 655 148 663
rect 76 641 98 655
rect 128 646 166 655
rect 172 655 178 670
rect 196 663 230 664
rect 204 655 208 663
rect 216 655 218 663
rect 226 655 230 663
rect 196 653 230 655
rect 76 635 94 641
rect 93 633 94 635
rect 102 633 103 641
rect 128 640 134 646
rect 93 631 103 633
rect 93 623 94 631
rect 102 623 103 631
rect 93 621 103 623
rect 93 613 94 621
rect 102 613 103 621
rect 93 611 103 613
rect 93 603 94 611
rect 102 603 103 611
rect 93 601 103 603
rect 93 593 94 601
rect 102 593 103 601
rect 93 591 103 593
rect 93 583 94 591
rect 102 583 103 591
rect 93 581 103 583
rect 93 573 94 581
rect 102 573 103 581
rect 93 571 103 573
rect 93 563 94 571
rect 102 563 103 571
rect 93 561 103 563
rect 93 553 94 561
rect 102 553 103 561
rect 110 639 118 640
rect 86 541 110 547
rect 125 633 134 640
rect 125 625 126 633
rect 125 623 134 625
rect 125 615 126 623
rect 125 613 134 615
rect 125 605 126 613
rect 125 603 134 605
rect 125 595 126 603
rect 125 593 134 595
rect 125 585 126 593
rect 125 583 134 585
rect 125 575 126 583
rect 125 573 134 575
rect 125 565 126 573
rect 125 563 134 565
rect 125 555 126 563
rect 142 639 150 640
rect 118 541 120 549
rect 48 535 54 541
rect 114 539 120 541
rect 157 637 166 646
rect 222 641 230 653
rect 174 640 182 641
rect 157 633 167 637
rect 157 625 158 633
rect 166 625 167 633
rect 157 623 167 625
rect 157 615 158 623
rect 166 615 167 623
rect 157 613 167 615
rect 157 605 158 613
rect 166 605 167 613
rect 157 603 167 605
rect 157 585 158 603
rect 166 585 167 603
rect 157 583 167 585
rect 157 565 158 583
rect 166 565 167 583
rect 157 563 167 565
rect 157 555 158 563
rect 166 555 167 563
rect 157 553 167 555
rect 157 545 158 553
rect 166 545 167 553
rect 142 539 150 541
rect 206 639 214 640
rect 189 633 199 637
rect 189 625 190 633
rect 198 625 199 633
rect 189 623 199 625
rect 189 615 190 623
rect 198 615 199 623
rect 189 613 199 615
rect 189 605 190 613
rect 198 605 199 613
rect 189 603 199 605
rect 189 595 190 603
rect 198 595 199 603
rect 189 593 199 595
rect 189 585 190 593
rect 198 585 199 593
rect 189 583 199 585
rect 189 575 190 583
rect 198 575 199 583
rect 189 573 199 575
rect 189 565 190 573
rect 198 565 199 573
rect 189 563 199 565
rect 189 555 190 563
rect 198 555 199 563
rect 189 553 199 555
rect 189 545 190 553
rect 198 545 199 553
rect 174 539 182 542
rect 222 631 230 633
rect 236 640 242 708
rect 248 695 268 697
rect 256 687 260 695
rect 248 686 268 687
rect 280 678 286 694
rect 254 655 260 670
rect 272 663 296 664
rect 272 655 274 663
rect 282 655 284 663
rect 292 655 296 663
rect 272 653 296 655
rect 302 641 308 708
rect 236 629 238 640
rect 222 621 230 623
rect 222 611 230 613
rect 222 601 230 603
rect 222 591 230 593
rect 222 581 230 583
rect 222 571 230 573
rect 222 561 230 563
rect 206 539 214 541
rect 221 542 238 547
rect 246 634 270 640
rect 270 629 278 632
rect 221 541 246 542
rect 254 623 262 627
rect 270 614 278 621
rect 262 545 286 550
rect 254 543 286 545
rect 294 635 308 641
rect 254 542 294 543
rect 302 619 310 621
rect 221 539 228 541
rect 0 532 16 534
rect 0 524 2 532
rect 10 524 16 532
rect 0 522 16 524
rect 0 514 2 522
rect 10 514 16 522
rect 0 512 16 514
rect 0 4 4 512
rect 12 12 16 512
rect 48 527 50 535
rect 114 533 228 539
rect 254 535 262 542
rect 234 529 262 535
rect 316 532 380 766
rect 436 760 442 767
rect 466 761 474 767
rect 498 767 570 773
rect 386 750 394 752
rect 386 740 394 742
rect 386 730 394 732
rect 386 720 394 722
rect 386 709 394 712
rect 410 754 434 760
rect 402 709 410 712
rect 418 728 426 730
rect 418 717 426 720
rect 388 697 394 709
rect 418 697 426 709
rect 388 693 426 697
rect 388 681 426 685
rect 434 709 442 712
rect 448 753 450 761
rect 448 751 458 753
rect 448 743 450 751
rect 448 741 458 743
rect 448 733 450 741
rect 448 731 458 733
rect 448 723 450 731
rect 448 721 458 723
rect 448 713 450 721
rect 448 709 458 713
rect 466 709 474 713
rect 482 761 490 765
rect 482 751 490 753
rect 482 741 490 743
rect 482 731 490 733
rect 482 721 490 723
rect 482 709 490 713
rect 498 761 506 767
rect 530 761 538 767
rect 562 761 570 767
rect 498 709 506 713
rect 514 751 522 753
rect 514 741 522 743
rect 514 731 522 733
rect 514 721 522 723
rect 434 678 440 709
rect 448 694 454 709
rect 484 697 490 709
rect 514 697 522 713
rect 388 663 426 665
rect 406 655 408 663
rect 416 655 418 663
rect 388 653 426 655
rect 388 637 394 653
rect 22 26 28 527
rect 34 516 72 521
rect 34 502 72 508
rect 34 484 72 486
rect 52 456 72 466
rect 34 454 72 456
rect 52 452 72 454
rect 52 446 64 452
rect 34 444 64 446
rect 52 443 72 444
rect 78 484 84 514
rect 78 472 86 476
rect 52 416 58 443
rect 78 434 84 464
rect 34 414 58 416
rect 52 406 58 414
rect 34 404 58 406
rect 52 376 58 404
rect 34 374 58 376
rect 52 366 58 374
rect 34 364 58 366
rect 52 336 58 364
rect 34 334 58 336
rect 52 326 58 334
rect 34 324 58 326
rect 52 296 58 324
rect 34 294 58 296
rect 52 286 58 294
rect 34 284 58 286
rect 52 256 58 284
rect 34 254 58 256
rect 52 246 58 254
rect 34 244 58 246
rect 52 216 58 244
rect 34 214 58 216
rect 52 206 58 214
rect 34 204 58 206
rect 52 176 58 204
rect 34 174 58 176
rect 52 166 58 174
rect 34 164 58 166
rect 52 136 58 164
rect 34 134 58 136
rect 52 126 58 134
rect 34 124 58 126
rect 52 96 58 124
rect 34 94 58 96
rect 52 86 58 94
rect 72 428 84 434
rect 34 84 58 86
rect 52 75 58 84
rect 52 72 78 75
rect 52 66 64 72
rect 34 64 64 66
rect 72 67 78 72
rect 72 64 86 67
rect 34 58 78 64
rect 42 50 48 58
rect 76 54 86 56
rect 76 50 78 54
rect 34 48 78 50
rect 42 40 48 48
rect 76 44 86 46
rect 76 40 78 44
rect 34 38 78 40
rect 34 32 48 38
rect 46 30 48 32
rect 76 32 86 36
rect 76 30 80 32
rect 46 28 80 30
rect 94 26 100 527
rect 114 526 228 527
rect 114 521 118 526
rect 106 518 118 521
rect 106 514 218 518
rect 106 506 108 514
rect 226 508 228 526
rect 106 502 214 506
rect 234 502 240 529
rect 269 523 380 532
rect 246 492 380 523
rect 386 633 394 637
rect 386 623 394 625
rect 386 613 394 615
rect 386 603 394 605
rect 386 583 394 585
rect 386 563 394 565
rect 386 553 394 555
rect 386 529 394 545
rect 402 633 410 641
rect 418 633 426 653
rect 418 623 426 625
rect 418 613 426 615
rect 418 603 426 605
rect 418 583 426 585
rect 418 563 426 565
rect 418 553 426 555
rect 434 641 440 670
rect 466 655 472 695
rect 484 693 522 697
rect 502 685 504 693
rect 512 685 514 693
rect 544 753 546 761
rect 544 751 554 753
rect 544 743 546 751
rect 544 741 554 743
rect 544 733 546 741
rect 544 731 554 733
rect 544 723 546 731
rect 544 721 554 723
rect 544 713 546 721
rect 484 663 522 665
rect 502 655 504 663
rect 512 655 514 663
rect 448 641 454 655
rect 484 653 522 655
rect 484 641 490 653
rect 434 633 442 641
rect 448 633 458 641
rect 448 625 450 633
rect 448 623 458 625
rect 448 615 450 623
rect 448 613 458 615
rect 448 605 450 613
rect 448 603 458 605
rect 448 585 450 603
rect 448 583 458 585
rect 448 565 450 583
rect 448 563 458 565
rect 448 555 450 563
rect 448 553 458 555
rect 448 545 450 553
rect 466 633 474 641
rect 402 535 410 545
rect 434 535 442 545
rect 466 535 474 545
rect 402 527 474 535
rect 386 516 460 521
rect 386 508 389 516
rect 457 508 460 516
rect 386 502 460 508
rect 386 494 389 502
rect 457 494 460 502
rect 466 500 474 527
rect 482 633 490 641
rect 482 623 490 625
rect 482 613 490 615
rect 482 603 490 605
rect 482 583 490 585
rect 482 563 490 565
rect 482 553 490 555
rect 482 529 490 545
rect 480 519 482 521
rect 498 633 506 641
rect 514 633 522 653
rect 514 623 522 625
rect 514 613 522 615
rect 514 603 522 605
rect 514 583 522 585
rect 514 563 522 565
rect 514 553 522 555
rect 530 641 536 713
rect 544 710 554 713
rect 544 697 550 710
rect 562 709 570 713
rect 578 765 590 773
rect 598 765 600 773
rect 578 763 600 765
rect 578 761 590 763
rect 586 755 590 761
rect 598 755 600 763
rect 586 753 600 755
rect 578 751 590 753
rect 586 745 590 751
rect 598 745 600 753
rect 586 743 600 745
rect 578 741 590 743
rect 586 735 590 741
rect 598 735 600 743
rect 586 733 600 735
rect 578 731 590 733
rect 586 725 590 731
rect 598 725 600 733
rect 586 723 600 725
rect 578 721 590 723
rect 586 715 590 721
rect 598 715 600 723
rect 586 713 600 715
rect 578 709 590 713
rect 580 705 590 709
rect 598 705 600 713
rect 588 703 600 705
rect 542 692 550 697
rect 580 695 590 697
rect 598 695 600 703
rect 542 683 550 684
rect 561 678 567 695
rect 580 693 600 695
rect 598 685 600 693
rect 580 683 600 685
rect 542 663 550 665
rect 561 655 567 670
rect 580 664 600 665
rect 542 653 550 655
rect 544 641 550 653
rect 580 646 590 656
rect 598 646 600 664
rect 580 644 600 646
rect 580 641 590 644
rect 530 633 538 641
rect 544 633 554 641
rect 544 625 546 633
rect 544 623 554 625
rect 544 615 546 623
rect 544 613 554 615
rect 544 605 546 613
rect 544 603 554 605
rect 544 585 546 603
rect 544 583 554 585
rect 544 565 546 583
rect 544 563 554 565
rect 544 555 546 563
rect 544 553 554 555
rect 544 545 546 553
rect 562 633 570 641
rect 498 535 506 545
rect 530 535 538 545
rect 562 535 570 545
rect 498 527 570 535
rect 578 636 590 641
rect 598 636 600 644
rect 578 634 600 636
rect 578 633 590 634
rect 586 626 590 633
rect 598 626 600 634
rect 586 625 600 626
rect 578 624 600 625
rect 578 623 590 624
rect 586 616 590 623
rect 598 616 600 624
rect 586 615 600 616
rect 578 614 600 615
rect 578 613 590 614
rect 586 606 590 613
rect 598 606 600 614
rect 586 605 600 606
rect 578 604 600 605
rect 578 603 590 604
rect 586 596 590 603
rect 598 596 600 604
rect 586 595 600 596
rect 578 594 600 595
rect 578 593 590 594
rect 586 586 590 593
rect 598 586 600 594
rect 586 585 600 586
rect 578 584 600 585
rect 578 583 590 584
rect 586 576 590 583
rect 598 576 600 584
rect 586 575 600 576
rect 578 574 600 575
rect 578 573 590 574
rect 586 566 590 573
rect 598 566 600 574
rect 586 565 600 566
rect 578 564 600 565
rect 578 563 590 564
rect 586 556 590 563
rect 598 556 600 564
rect 586 555 600 556
rect 578 554 600 555
rect 578 553 590 554
rect 586 546 590 553
rect 598 546 600 554
rect 586 545 600 546
rect 578 544 600 545
rect 578 541 590 544
rect 578 533 580 541
rect 598 536 600 544
rect 588 534 600 536
rect 588 533 590 534
rect 578 531 590 533
rect 490 519 508 521
rect 480 507 508 511
rect 466 492 506 500
rect 246 488 352 492
rect 106 458 108 468
rect 126 466 138 468
rect 126 458 128 466
rect 136 458 138 466
rect 156 466 168 468
rect 156 458 158 466
rect 166 458 168 466
rect 186 466 198 468
rect 186 458 188 466
rect 196 458 198 466
rect 216 466 228 468
rect 234 466 240 486
rect 216 458 218 466
rect 226 458 228 466
rect 236 458 240 466
rect 106 454 240 458
rect 106 446 108 454
rect 126 446 128 454
rect 136 446 138 454
rect 156 446 158 454
rect 166 446 168 454
rect 186 446 188 454
rect 196 446 198 454
rect 216 446 218 454
rect 226 446 228 454
rect 236 446 240 454
rect 106 429 240 446
rect 106 421 108 429
rect 236 421 240 429
rect 106 419 240 421
rect 246 411 286 488
rect 106 400 286 411
rect 106 392 112 400
rect 240 392 286 400
rect 106 388 286 392
rect 106 380 112 388
rect 240 380 286 388
rect 106 371 286 380
rect 106 362 240 365
rect 106 354 112 362
rect 106 334 240 354
rect 106 326 110 334
rect 128 326 130 334
rect 138 326 140 334
rect 158 326 160 334
rect 168 326 170 334
rect 188 326 190 334
rect 198 326 200 334
rect 218 326 220 334
rect 228 326 230 334
rect 238 326 240 334
rect 106 322 240 326
rect 106 314 110 322
rect 128 314 130 322
rect 138 314 140 322
rect 158 314 160 322
rect 168 314 170 322
rect 188 314 190 322
rect 198 314 200 322
rect 218 314 220 322
rect 228 314 230 322
rect 238 314 240 322
rect 106 296 240 314
rect 106 288 110 296
rect 238 288 240 296
rect 106 286 240 288
rect 246 278 286 371
rect 112 268 286 278
rect 240 250 286 268
rect 112 241 286 250
rect 106 232 240 234
rect 106 224 110 232
rect 238 224 240 232
rect 106 204 240 224
rect 106 196 109 204
rect 127 196 129 204
rect 137 196 139 204
rect 157 196 159 204
rect 167 196 169 204
rect 187 196 189 204
rect 197 196 199 204
rect 217 196 219 204
rect 227 196 229 204
rect 237 196 240 204
rect 106 192 240 196
rect 106 184 109 192
rect 127 184 129 192
rect 137 184 139 192
rect 157 184 159 192
rect 167 184 169 192
rect 187 184 189 192
rect 197 184 199 192
rect 217 184 219 192
rect 227 184 229 192
rect 237 184 240 192
rect 106 168 240 184
rect 106 160 110 168
rect 238 160 240 168
rect 106 157 240 160
rect 246 148 286 241
rect 106 138 286 148
rect 106 120 112 138
rect 240 120 286 138
rect 106 112 286 120
rect 107 102 238 105
rect 107 94 108 102
rect 236 94 238 102
rect 107 74 238 94
rect 115 66 118 74
rect 236 66 238 74
rect 107 64 238 66
rect 115 62 238 64
rect 115 36 118 62
rect 114 34 118 36
rect 126 34 128 62
rect 136 34 138 62
rect 146 34 148 62
rect 156 34 158 62
rect 166 34 168 62
rect 176 34 178 62
rect 186 34 188 62
rect 196 34 198 62
rect 206 34 208 62
rect 216 34 218 62
rect 226 34 228 62
rect 236 34 238 62
rect 114 28 238 34
rect 246 98 286 112
rect 294 478 306 481
rect 294 460 296 478
rect 304 460 306 478
rect 294 458 306 460
rect 294 450 296 458
rect 304 450 306 458
rect 294 448 306 450
rect 294 430 296 448
rect 304 430 306 448
rect 294 428 306 430
rect 294 420 296 428
rect 304 420 306 428
rect 294 418 306 420
rect 294 400 296 418
rect 304 400 306 418
rect 294 398 306 400
rect 294 390 296 398
rect 304 390 306 398
rect 294 388 306 390
rect 294 370 296 388
rect 304 370 306 388
rect 294 368 306 370
rect 294 360 296 368
rect 304 360 306 368
rect 294 358 306 360
rect 294 340 296 358
rect 304 340 306 358
rect 294 338 306 340
rect 294 330 296 338
rect 304 330 306 338
rect 294 328 306 330
rect 294 310 296 328
rect 304 310 306 328
rect 294 308 306 310
rect 294 300 296 308
rect 304 300 306 308
rect 294 288 306 300
rect 294 280 296 288
rect 304 280 306 288
rect 294 278 306 280
rect 294 270 296 278
rect 304 270 306 278
rect 294 268 306 270
rect 294 250 296 268
rect 304 250 306 268
rect 294 248 306 250
rect 294 240 296 248
rect 304 240 306 248
rect 294 238 306 240
rect 294 220 296 238
rect 304 220 306 238
rect 294 218 306 220
rect 294 210 296 218
rect 304 210 306 218
rect 294 208 306 210
rect 294 190 296 208
rect 304 190 306 208
rect 294 188 306 190
rect 294 180 296 188
rect 304 180 306 188
rect 294 178 306 180
rect 294 170 296 178
rect 304 170 306 178
rect 294 158 306 170
rect 294 150 296 158
rect 304 150 306 158
rect 294 148 306 150
rect 294 130 296 148
rect 304 130 306 148
rect 294 128 306 130
rect 294 120 296 128
rect 304 120 306 128
rect 294 118 306 120
rect 294 110 296 118
rect 304 110 306 118
rect 294 108 306 110
rect 314 411 352 488
rect 359 458 364 486
rect 382 466 394 468
rect 382 458 384 466
rect 392 458 394 466
rect 412 466 424 468
rect 412 458 414 466
rect 422 458 424 466
rect 442 466 454 468
rect 442 458 444 466
rect 452 458 454 466
rect 472 466 484 468
rect 472 458 474 466
rect 482 458 484 466
rect 492 458 494 486
rect 359 454 494 458
rect 359 446 364 454
rect 382 446 384 454
rect 392 446 394 454
rect 412 446 414 454
rect 422 446 424 454
rect 442 446 444 454
rect 452 446 454 454
rect 472 446 474 454
rect 482 446 484 454
rect 492 446 494 454
rect 359 429 494 446
rect 359 421 364 429
rect 492 421 494 429
rect 359 419 494 421
rect 314 400 494 411
rect 314 392 360 400
rect 488 392 494 400
rect 314 388 494 392
rect 314 380 360 388
rect 488 380 494 388
rect 314 371 494 380
rect 314 278 352 371
rect 360 362 494 365
rect 360 354 364 362
rect 492 354 494 362
rect 360 335 494 354
rect 360 327 363 335
rect 381 327 383 335
rect 391 327 393 335
rect 411 327 413 335
rect 421 327 423 335
rect 441 327 443 335
rect 451 327 453 335
rect 471 327 473 335
rect 481 327 483 335
rect 491 327 494 335
rect 360 323 494 327
rect 360 315 363 323
rect 381 315 383 323
rect 391 315 393 323
rect 411 315 413 323
rect 421 315 423 323
rect 441 315 443 323
rect 451 315 453 323
rect 471 315 473 323
rect 481 315 483 323
rect 491 315 494 323
rect 360 296 494 315
rect 360 288 363 296
rect 491 288 494 296
rect 360 286 494 288
rect 314 268 494 278
rect 314 250 360 268
rect 488 250 494 268
rect 314 241 494 250
rect 314 148 352 241
rect 360 231 494 234
rect 360 223 364 231
rect 492 223 494 231
rect 360 204 494 223
rect 360 196 364 204
rect 382 196 384 204
rect 392 196 394 204
rect 412 196 414 204
rect 422 196 424 204
rect 442 196 444 204
rect 452 196 454 204
rect 472 196 474 204
rect 482 196 484 204
rect 492 196 494 204
rect 360 192 494 196
rect 360 184 364 192
rect 382 184 384 192
rect 392 184 394 192
rect 412 184 414 192
rect 422 184 424 192
rect 442 184 444 192
rect 452 184 454 192
rect 472 184 474 192
rect 482 184 484 192
rect 492 184 494 192
rect 360 168 494 184
rect 360 160 364 168
rect 492 160 494 168
rect 360 157 494 160
rect 314 138 494 148
rect 314 120 360 138
rect 488 120 494 138
rect 314 112 494 120
rect 314 98 352 112
rect 246 38 352 98
rect 246 30 256 38
rect 344 30 352 38
rect 246 25 352 30
rect 360 103 494 105
rect 360 95 364 103
rect 492 95 494 103
rect 360 74 494 95
rect 360 66 364 74
rect 492 66 494 74
rect 360 64 494 66
rect 360 62 474 64
rect 360 34 364 62
rect 372 34 374 62
rect 382 34 384 62
rect 392 34 394 62
rect 402 34 404 62
rect 412 34 414 62
rect 422 34 424 62
rect 432 34 434 62
rect 442 34 444 62
rect 452 34 454 62
rect 462 34 464 62
rect 472 36 474 62
rect 482 36 484 64
rect 492 36 494 64
rect 472 34 494 36
rect 360 32 494 34
rect 360 28 482 32
rect 500 26 506 492
rect 514 26 520 527
rect 578 521 580 531
rect 598 526 600 534
rect 588 524 600 526
rect 535 513 540 521
rect 588 516 590 524
rect 598 516 600 524
rect 588 513 600 516
rect 527 512 600 513
rect 527 502 590 512
rect 575 494 580 502
rect 542 484 572 486
rect 527 472 535 476
rect 528 434 535 464
rect 560 466 572 484
rect 542 461 572 466
rect 560 459 572 461
rect 560 453 564 459
rect 542 451 564 453
rect 560 443 564 451
rect 542 441 564 443
rect 560 413 564 441
rect 542 411 564 413
rect 560 403 564 411
rect 542 401 564 403
rect 560 373 564 401
rect 542 371 564 373
rect 560 363 564 371
rect 542 361 564 363
rect 560 333 564 361
rect 542 331 564 333
rect 560 323 564 331
rect 542 321 564 323
rect 560 293 564 321
rect 542 291 564 293
rect 560 283 564 291
rect 542 281 564 283
rect 560 253 564 281
rect 542 251 564 253
rect 560 243 564 251
rect 542 241 564 243
rect 560 213 564 241
rect 542 211 564 213
rect 560 203 564 211
rect 542 201 564 203
rect 560 173 564 201
rect 542 171 564 173
rect 560 163 564 171
rect 542 161 564 163
rect 560 133 564 161
rect 542 131 564 133
rect 560 123 564 131
rect 542 121 564 123
rect 560 93 564 121
rect 542 91 564 93
rect 560 83 564 91
rect 542 81 564 83
rect 526 73 542 75
rect 526 65 528 73
rect 536 65 542 73
rect 526 63 542 65
rect 560 63 564 81
rect 526 58 564 63
rect 544 50 552 58
rect 560 50 564 58
rect 526 48 564 50
rect 526 40 536 48
rect 544 40 552 48
rect 560 40 564 48
rect 534 38 564 40
rect 534 32 552 38
rect 538 30 552 32
rect 560 31 564 38
rect 560 30 572 31
rect 538 28 572 30
rect 578 16 580 494
rect 48 12 82 16
rect 113 12 482 16
rect 538 12 580 16
rect 12 10 56 12
rect 74 10 116 12
rect 0 2 14 4
rect 42 2 46 10
rect 334 4 338 12
rect 476 10 538 12
rect 586 4 590 14
rect 598 4 600 512
rect 54 2 76 4
rect 114 2 478 4
rect 536 2 600 4
rect 0 0 600 2
<< m2contact >>
rect 28 1300 226 1308
rect 28 880 36 1300
rect 40 1282 88 1290
rect 60 1262 88 1282
rect 122 1262 130 1290
rect 152 1262 160 1290
rect 182 1262 190 1290
rect 212 1262 220 1290
rect 40 1242 58 1250
rect 64 1243 72 1251
rect 84 1236 232 1244
rect 40 1202 58 1210
rect 82 1185 100 1233
rect 40 1162 58 1170
rect 40 1122 58 1130
rect 64 1111 72 1179
rect 84 1172 232 1180
rect 83 1144 121 1152
rect 143 1144 151 1152
rect 173 1144 181 1152
rect 203 1144 211 1152
rect 83 1132 121 1140
rect 143 1132 151 1140
rect 173 1132 181 1140
rect 203 1132 211 1140
rect 84 1105 232 1113
rect 40 1082 58 1090
rect 84 1055 102 1105
rect 40 1042 58 1050
rect 40 1002 58 1010
rect 64 981 72 1049
rect 84 1044 232 1052
rect 82 1016 120 1024
rect 142 1016 150 1024
rect 172 1016 180 1024
rect 202 1016 210 1024
rect 82 1004 120 1012
rect 142 1004 150 1012
rect 172 1004 180 1012
rect 202 1004 210 1012
rect 84 978 232 986
rect 40 962 58 970
rect 40 922 58 930
rect 40 882 58 890
rect 84 927 102 975
rect 82 914 230 922
rect 80 886 88 894
rect 91 886 99 894
rect 102 886 110 894
rect 113 886 121 894
rect 143 886 151 894
rect 173 886 181 894
rect 203 886 211 894
rect 93 874 101 882
rect 113 874 121 882
rect 143 874 151 882
rect 173 874 181 882
rect 203 874 211 882
rect 64 862 82 870
rect 30 842 58 850
rect 14 790 22 818
rect 26 810 54 818
rect 78 842 226 850
rect 78 810 216 818
rect 296 1276 304 1284
rect 296 1236 304 1244
rect 296 1196 304 1204
rect 296 1156 304 1164
rect 296 1116 304 1124
rect 296 1076 304 1084
rect 296 1036 304 1044
rect 296 996 304 1004
rect 296 956 304 964
rect 296 916 304 924
rect 296 876 304 884
rect 374 1302 572 1310
rect 376 1262 384 1290
rect 406 1262 414 1290
rect 436 1262 444 1290
rect 466 1262 474 1290
rect 508 1262 536 1290
rect 542 1282 560 1290
rect 368 1236 516 1244
rect 528 1242 536 1250
rect 542 1242 560 1250
rect 498 1181 516 1229
rect 542 1202 560 1210
rect 368 1170 516 1178
rect 388 1144 396 1152
rect 418 1144 426 1152
rect 448 1144 456 1152
rect 478 1144 516 1152
rect 388 1132 396 1140
rect 418 1132 426 1140
rect 448 1132 456 1140
rect 478 1132 516 1140
rect 368 1106 516 1114
rect 528 1108 536 1176
rect 542 1162 560 1170
rect 542 1122 560 1130
rect 498 1055 516 1103
rect 542 1082 560 1090
rect 368 1044 516 1052
rect 387 1016 395 1024
rect 417 1016 425 1024
rect 447 1016 455 1024
rect 477 1016 515 1024
rect 387 1004 395 1012
rect 417 1004 425 1012
rect 447 1004 455 1012
rect 477 1004 515 1012
rect 368 978 516 986
rect 528 981 536 1049
rect 542 1042 560 1050
rect 542 1002 560 1010
rect 296 842 304 850
rect 500 926 518 974
rect 370 914 518 922
rect 389 886 397 894
rect 419 886 427 894
rect 449 886 457 894
rect 479 886 487 894
rect 490 886 498 894
rect 501 886 509 894
rect 512 886 520 894
rect 389 874 397 882
rect 419 874 427 882
rect 449 874 457 882
rect 479 874 487 882
rect 499 874 507 882
rect 518 862 536 870
rect 542 962 560 970
rect 542 922 560 930
rect 542 882 560 890
rect 564 882 572 1302
rect 368 842 576 850
rect 590 815 598 823
rect 14 708 22 786
rect 590 795 598 803
rect 576 776 584 784
rect 590 775 598 783
rect 44 742 52 750
rect 44 722 52 730
rect 94 738 102 746
rect 94 718 102 726
rect 126 738 134 746
rect 126 718 134 726
rect 158 738 166 746
rect 158 718 166 726
rect 190 738 198 746
rect 190 718 198 726
rect 222 738 230 746
rect 222 718 230 726
rect 238 720 246 728
rect 40 670 58 678
rect 2 634 10 642
rect 2 614 10 622
rect 2 594 10 602
rect 2 574 10 582
rect 2 554 10 562
rect 14 548 22 636
rect 2 534 10 542
rect 44 623 52 631
rect 44 603 52 611
rect 44 583 52 591
rect 44 563 52 571
rect 206 687 214 695
rect 270 720 278 728
rect 184 670 202 678
rect 138 655 146 663
rect 208 655 216 663
rect 94 623 102 631
rect 94 603 102 611
rect 94 583 102 591
rect 94 563 102 571
rect 126 615 134 623
rect 126 595 134 603
rect 126 575 134 583
rect 126 555 134 563
rect 158 615 166 623
rect 158 585 166 603
rect 158 555 166 563
rect 190 615 198 623
rect 190 595 198 603
rect 190 575 198 583
rect 190 555 198 563
rect 222 623 230 631
rect 260 687 268 695
rect 248 670 266 678
rect 284 655 292 663
rect 222 603 230 611
rect 222 583 230 591
rect 222 563 230 571
rect 270 621 278 629
rect 302 621 310 629
rect 2 514 10 522
rect 386 742 394 750
rect 386 722 394 730
rect 418 720 426 728
rect 388 673 426 681
rect 450 743 458 751
rect 450 723 458 731
rect 482 743 490 751
rect 482 723 490 731
rect 514 743 522 751
rect 514 723 522 731
rect 434 670 452 678
rect 408 655 416 663
rect 34 494 72 502
rect 34 446 52 454
rect 64 444 72 452
rect 78 476 86 484
rect 78 464 86 472
rect 34 406 52 414
rect 34 366 52 374
rect 34 326 52 334
rect 34 286 52 294
rect 34 246 52 254
rect 34 206 52 214
rect 34 166 52 174
rect 34 126 52 134
rect 34 86 52 94
rect 64 64 72 72
rect 78 48 86 54
rect 34 40 42 48
rect 48 46 86 48
rect 48 40 76 46
rect 106 494 214 502
rect 222 494 240 502
rect 386 615 394 623
rect 386 585 394 603
rect 386 555 394 563
rect 418 615 426 623
rect 418 585 426 603
rect 418 555 426 563
rect 504 685 512 693
rect 546 743 554 751
rect 546 723 554 731
rect 504 655 512 663
rect 450 615 458 623
rect 450 585 458 603
rect 450 555 458 563
rect 389 494 457 502
rect 482 615 490 623
rect 482 585 490 603
rect 482 555 490 563
rect 514 615 522 623
rect 514 585 522 603
rect 514 555 522 563
rect 590 755 598 763
rect 578 743 586 751
rect 590 735 598 743
rect 578 723 586 731
rect 590 715 598 723
rect 580 703 588 705
rect 580 697 598 703
rect 590 695 598 697
rect 555 670 573 678
rect 546 615 554 623
rect 546 585 554 603
rect 546 555 554 563
rect 590 636 598 644
rect 578 615 586 623
rect 590 616 598 624
rect 578 595 586 603
rect 590 596 598 604
rect 578 575 586 583
rect 590 576 598 584
rect 578 555 586 563
rect 590 556 598 564
rect 590 541 598 544
rect 580 536 598 541
rect 580 533 588 536
rect 128 458 136 466
rect 158 458 166 466
rect 188 458 196 466
rect 218 458 226 466
rect 128 446 136 454
rect 158 446 166 454
rect 188 446 196 454
rect 218 446 226 454
rect 108 421 236 429
rect 112 354 240 362
rect 130 326 138 334
rect 160 326 168 334
rect 190 326 198 334
rect 220 326 228 334
rect 130 314 138 322
rect 160 314 168 322
rect 190 314 198 322
rect 220 314 228 322
rect 110 288 238 296
rect 110 224 238 232
rect 129 196 137 204
rect 159 196 167 204
rect 189 196 197 204
rect 219 196 227 204
rect 129 184 137 192
rect 159 184 167 192
rect 189 184 197 192
rect 219 184 227 192
rect 110 160 238 168
rect 108 94 236 102
rect 118 34 126 62
rect 138 34 146 62
rect 158 34 166 62
rect 178 34 186 62
rect 198 34 206 62
rect 218 34 226 62
rect 296 450 304 458
rect 296 420 304 428
rect 296 390 304 398
rect 296 360 304 368
rect 296 330 304 338
rect 296 300 304 308
rect 296 270 304 278
rect 296 240 304 248
rect 296 210 304 218
rect 296 180 304 188
rect 296 150 304 158
rect 296 120 304 128
rect 384 458 392 466
rect 414 458 422 466
rect 444 458 452 466
rect 474 458 482 466
rect 384 446 392 454
rect 414 446 422 454
rect 444 446 452 454
rect 474 446 482 454
rect 364 421 492 429
rect 364 354 492 362
rect 383 327 391 335
rect 413 327 421 335
rect 443 327 451 335
rect 473 327 481 335
rect 383 315 391 323
rect 413 315 421 323
rect 443 315 451 323
rect 473 315 481 323
rect 363 288 491 296
rect 364 223 492 231
rect 384 196 392 204
rect 414 196 422 204
rect 444 196 452 204
rect 474 196 482 204
rect 384 184 392 192
rect 414 184 422 192
rect 444 184 452 192
rect 474 184 482 192
rect 364 160 492 168
rect 256 30 344 38
rect 22 18 40 26
rect 88 18 106 26
rect 364 95 492 103
rect 374 34 382 62
rect 394 34 402 62
rect 414 34 422 62
rect 434 34 442 62
rect 454 34 462 62
rect 474 36 482 64
rect 488 18 506 26
rect 590 516 598 524
rect 527 494 575 502
rect 527 476 535 484
rect 527 464 535 472
rect 542 443 560 451
rect 542 403 560 411
rect 542 363 560 371
rect 542 323 560 331
rect 542 283 560 291
rect 542 243 560 251
rect 542 203 560 211
rect 542 163 560 171
rect 542 123 560 131
rect 542 83 560 91
rect 528 65 536 73
rect 536 40 544 48
rect 552 40 560 48
rect 564 31 572 459
rect 514 18 532 26
<< metal2 >>
rect 0 1310 600 1340
rect 0 1308 374 1310
rect 0 880 28 1308
rect 226 1302 374 1308
rect 226 1300 564 1302
rect 36 1290 564 1300
rect 36 1282 40 1290
rect 36 1262 60 1282
rect 88 1262 122 1290
rect 130 1262 152 1290
rect 160 1262 182 1290
rect 190 1262 212 1290
rect 220 1284 376 1290
rect 220 1276 296 1284
rect 304 1276 376 1284
rect 220 1262 376 1276
rect 384 1262 406 1290
rect 414 1262 436 1290
rect 444 1262 466 1290
rect 474 1262 508 1290
rect 536 1282 542 1290
rect 560 1282 564 1290
rect 536 1262 564 1282
rect 36 1251 564 1262
rect 36 1250 64 1251
rect 36 1242 40 1250
rect 58 1243 64 1250
rect 72 1250 564 1251
rect 72 1244 528 1250
rect 72 1243 84 1244
rect 58 1242 84 1243
rect 36 1236 84 1242
rect 232 1236 296 1244
rect 304 1236 368 1244
rect 516 1242 528 1244
rect 536 1242 542 1250
rect 560 1242 564 1250
rect 516 1236 564 1242
rect 36 1233 564 1236
rect 36 1210 82 1233
rect 36 1202 40 1210
rect 58 1202 82 1210
rect 36 1185 82 1202
rect 100 1229 564 1233
rect 100 1204 498 1229
rect 100 1196 296 1204
rect 304 1196 498 1204
rect 100 1190 498 1196
rect 100 1185 104 1190
rect 36 1180 104 1185
rect 284 1180 316 1190
rect 497 1181 498 1190
rect 516 1210 564 1229
rect 516 1202 542 1210
rect 560 1202 564 1210
rect 516 1181 564 1202
rect 497 1180 564 1181
rect 36 1179 84 1180
rect 36 1170 64 1179
rect 36 1162 40 1170
rect 58 1162 64 1170
rect 36 1130 64 1162
rect 36 1122 40 1130
rect 58 1122 64 1130
rect 36 1111 64 1122
rect 72 1172 84 1179
rect 232 1178 564 1180
rect 232 1172 368 1178
rect 72 1170 368 1172
rect 516 1176 564 1178
rect 516 1170 528 1176
rect 72 1164 528 1170
rect 72 1156 296 1164
rect 304 1156 528 1164
rect 72 1152 528 1156
rect 72 1144 83 1152
rect 121 1144 143 1152
rect 151 1144 173 1152
rect 181 1144 203 1152
rect 211 1144 388 1152
rect 396 1144 418 1152
rect 426 1144 448 1152
rect 456 1144 478 1152
rect 516 1144 528 1152
rect 72 1140 528 1144
rect 72 1132 83 1140
rect 121 1132 143 1140
rect 151 1132 173 1140
rect 181 1132 203 1140
rect 211 1132 388 1140
rect 396 1132 418 1140
rect 426 1132 448 1140
rect 456 1132 478 1140
rect 516 1132 528 1140
rect 72 1124 528 1132
rect 72 1116 296 1124
rect 304 1116 528 1124
rect 72 1114 528 1116
rect 72 1113 368 1114
rect 72 1111 84 1113
rect 36 1090 84 1111
rect 232 1106 368 1113
rect 516 1108 528 1114
rect 536 1170 564 1176
rect 536 1162 542 1170
rect 560 1162 564 1170
rect 536 1130 564 1162
rect 536 1122 542 1130
rect 560 1122 564 1130
rect 536 1108 564 1122
rect 516 1106 564 1108
rect 232 1105 564 1106
rect 36 1082 40 1090
rect 58 1082 84 1090
rect 36 1055 84 1082
rect 102 1103 564 1105
rect 102 1084 498 1103
rect 102 1076 296 1084
rect 304 1076 498 1084
rect 102 1055 498 1076
rect 516 1090 564 1103
rect 516 1082 542 1090
rect 560 1082 564 1090
rect 516 1055 564 1082
rect 36 1052 564 1055
rect 36 1050 84 1052
rect 36 1042 40 1050
rect 58 1049 84 1050
rect 58 1042 64 1049
rect 36 1010 64 1042
rect 36 1002 40 1010
rect 58 1002 64 1010
rect 36 981 64 1002
rect 72 1044 84 1049
rect 232 1044 368 1052
rect 516 1050 564 1052
rect 516 1049 542 1050
rect 516 1044 528 1049
rect 72 1040 296 1044
rect 72 1030 104 1040
rect 284 1036 296 1040
rect 304 1040 528 1044
rect 304 1036 316 1040
rect 284 1030 316 1036
rect 500 1030 528 1040
rect 72 1024 528 1030
rect 72 1016 82 1024
rect 120 1016 142 1024
rect 150 1016 172 1024
rect 180 1016 202 1024
rect 210 1016 387 1024
rect 395 1016 417 1024
rect 425 1016 447 1024
rect 455 1016 477 1024
rect 515 1016 528 1024
rect 72 1012 528 1016
rect 72 1004 82 1012
rect 120 1004 142 1012
rect 150 1004 172 1012
rect 180 1004 202 1012
rect 210 1004 387 1012
rect 395 1004 417 1012
rect 425 1004 447 1012
rect 455 1004 477 1012
rect 515 1004 528 1012
rect 72 996 296 1004
rect 304 996 528 1004
rect 72 986 528 996
rect 72 981 84 986
rect 36 978 84 981
rect 232 978 368 986
rect 516 981 528 986
rect 536 1042 542 1049
rect 560 1042 564 1050
rect 536 1010 564 1042
rect 536 1002 542 1010
rect 560 1002 564 1010
rect 536 981 564 1002
rect 516 978 564 981
rect 36 975 564 978
rect 36 970 84 975
rect 36 962 40 970
rect 58 962 84 970
rect 36 930 84 962
rect 36 922 40 930
rect 58 927 84 930
rect 102 974 564 975
rect 102 964 500 974
rect 102 956 296 964
rect 304 956 500 964
rect 102 927 500 956
rect 58 926 500 927
rect 518 970 564 974
rect 518 962 542 970
rect 560 962 564 970
rect 518 930 564 962
rect 518 926 542 930
rect 58 924 542 926
rect 58 922 296 924
rect 36 914 82 922
rect 230 916 296 922
rect 304 922 542 924
rect 560 922 564 930
rect 304 916 370 922
rect 230 914 370 916
rect 518 914 564 922
rect 36 894 564 914
rect 36 890 80 894
rect 36 882 40 890
rect 58 886 80 890
rect 88 886 91 894
rect 99 886 102 894
rect 110 886 113 894
rect 121 886 143 894
rect 151 886 173 894
rect 181 886 203 894
rect 211 886 389 894
rect 397 886 419 894
rect 427 886 449 894
rect 457 886 479 894
rect 487 886 490 894
rect 498 886 501 894
rect 509 886 512 894
rect 520 890 564 894
rect 520 886 542 890
rect 58 884 542 886
rect 58 882 296 884
rect 36 880 93 882
rect 0 878 58 880
rect 90 874 93 880
rect 101 874 113 882
rect 121 874 143 882
rect 151 874 173 882
rect 181 874 203 882
rect 211 876 296 882
rect 304 882 542 884
rect 560 882 564 890
rect 572 882 600 1310
rect 304 876 389 882
rect 211 874 389 876
rect 397 874 419 882
rect 427 874 449 882
rect 457 874 479 882
rect 487 874 499 882
rect 507 880 600 882
rect 507 874 510 880
rect 542 878 600 880
rect 64 870 82 872
rect 518 870 536 872
rect 82 862 518 866
rect 64 860 536 862
rect 72 858 536 860
rect 20 845 30 850
rect 0 842 30 845
rect 58 842 78 850
rect 226 842 296 850
rect 304 842 368 850
rect 576 842 600 845
rect 0 823 600 842
rect 0 818 590 823
rect 0 790 14 818
rect 22 810 26 818
rect 54 810 78 818
rect 216 815 590 818
rect 598 815 600 823
rect 216 810 600 815
rect 22 803 600 810
rect 22 795 590 803
rect 598 795 600 803
rect 22 790 600 795
rect 0 786 600 790
rect 0 708 14 786
rect 22 784 600 786
rect 22 777 576 784
rect 22 767 68 777
rect 123 767 163 777
rect 238 767 280 777
rect 381 767 421 777
rect 500 776 576 777
rect 584 783 600 784
rect 584 776 590 783
rect 500 775 590 776
rect 598 775 600 783
rect 500 767 600 775
rect 22 763 600 767
rect 22 755 590 763
rect 598 755 600 763
rect 22 751 600 755
rect 22 750 450 751
rect 22 742 44 750
rect 52 746 386 750
rect 52 742 94 746
rect 22 738 94 742
rect 102 738 126 746
rect 134 738 158 746
rect 166 738 190 746
rect 198 738 222 746
rect 230 742 386 746
rect 394 743 450 750
rect 458 743 482 751
rect 490 743 514 751
rect 522 743 546 751
rect 554 743 578 751
rect 586 743 600 751
rect 394 742 590 743
rect 230 738 590 742
rect 22 737 590 738
rect 22 730 230 737
rect 22 722 44 730
rect 52 726 230 730
rect 286 735 590 737
rect 598 735 600 743
rect 286 731 600 735
rect 286 730 450 731
rect 52 722 94 726
rect 22 718 94 722
rect 102 718 126 726
rect 134 718 158 726
rect 166 718 190 726
rect 198 718 222 726
rect 246 720 270 728
rect 286 722 386 730
rect 394 728 450 730
rect 394 722 418 728
rect 286 720 418 722
rect 426 723 450 728
rect 458 723 482 731
rect 490 723 514 731
rect 522 723 546 731
rect 554 723 578 731
rect 586 723 600 731
rect 426 720 590 723
rect 22 710 230 718
rect 286 715 590 720
rect 598 715 600 723
rect 286 710 600 715
rect 22 708 600 710
rect 0 705 600 708
rect 0 697 580 705
rect 588 703 600 705
rect 0 695 590 697
rect 598 695 600 703
rect 0 687 206 695
rect 214 687 260 695
rect 268 693 600 695
rect 268 687 504 693
rect 0 686 504 687
rect 273 683 426 686
rect 484 685 504 686
rect 512 686 600 693
rect 512 685 522 686
rect 388 681 426 683
rect 58 671 184 677
rect 202 671 248 677
rect 452 671 555 677
rect 273 663 426 665
rect 16 662 36 663
rect 62 662 138 663
rect 16 655 138 662
rect 146 662 180 663
rect 206 662 208 663
rect 146 655 208 662
rect 216 655 230 663
rect 16 652 230 655
rect 273 655 284 663
rect 292 655 408 663
rect 416 659 426 663
rect 484 659 504 663
rect 416 655 504 659
rect 512 655 522 663
rect 273 652 522 655
rect 0 644 600 652
rect 0 642 590 644
rect 0 634 2 642
rect 10 637 590 642
rect 10 636 262 637
rect 10 634 14 636
rect 0 622 14 634
rect 0 614 2 622
rect 10 614 14 622
rect 0 602 14 614
rect 0 594 2 602
rect 10 594 14 602
rect 0 582 14 594
rect 0 574 2 582
rect 10 574 14 582
rect 0 562 14 574
rect 0 554 2 562
rect 10 554 14 562
rect 0 548 14 554
rect 22 631 262 636
rect 22 623 44 631
rect 52 623 94 631
rect 102 623 222 631
rect 230 623 262 631
rect 318 636 590 637
rect 598 636 600 644
rect 22 615 126 623
rect 134 615 158 623
rect 166 615 190 623
rect 198 615 262 623
rect 278 621 302 629
rect 318 624 600 636
rect 318 623 590 624
rect 22 612 262 615
rect 318 615 386 623
rect 394 615 418 623
rect 426 615 450 623
rect 458 615 482 623
rect 490 615 514 623
rect 522 615 546 623
rect 554 615 578 623
rect 586 616 590 623
rect 598 616 600 624
rect 586 615 600 616
rect 318 612 600 615
rect 22 611 600 612
rect 22 603 44 611
rect 52 603 94 611
rect 102 603 222 611
rect 230 604 600 611
rect 230 603 590 604
rect 22 595 126 603
rect 134 595 158 603
rect 22 591 158 595
rect 22 583 44 591
rect 52 583 94 591
rect 102 585 158 591
rect 166 595 190 603
rect 198 595 386 603
rect 166 591 386 595
rect 166 585 222 591
rect 102 583 222 585
rect 230 585 386 591
rect 394 585 418 603
rect 426 585 450 603
rect 458 585 482 603
rect 490 585 514 603
rect 522 585 546 603
rect 554 595 578 603
rect 586 596 590 603
rect 598 596 600 604
rect 586 595 600 596
rect 554 585 600 595
rect 230 584 600 585
rect 230 583 590 584
rect 22 582 126 583
rect 22 572 36 582
rect 92 575 126 582
rect 134 582 190 583
rect 134 575 136 582
rect 92 572 136 575
rect 188 575 190 582
rect 198 582 578 583
rect 198 575 232 582
rect 188 572 232 575
rect 336 572 379 582
rect 447 572 490 582
rect 561 575 578 582
rect 586 576 590 583
rect 598 576 600 584
rect 586 575 600 576
rect 561 572 600 575
rect 22 571 600 572
rect 22 563 44 571
rect 52 563 94 571
rect 102 563 222 571
rect 230 564 600 571
rect 230 563 590 564
rect 22 555 126 563
rect 134 555 158 563
rect 166 555 190 563
rect 198 555 386 563
rect 394 555 418 563
rect 426 555 450 563
rect 458 555 482 563
rect 490 555 514 563
rect 522 555 546 563
rect 554 555 578 563
rect 586 556 590 563
rect 598 556 600 564
rect 586 555 600 556
rect 22 548 600 555
rect 0 544 600 548
rect 0 542 590 544
rect 0 534 2 542
rect 10 541 590 542
rect 10 534 580 541
rect 598 536 600 544
rect 0 533 580 534
rect 588 533 600 536
rect 0 524 600 533
rect 0 522 590 524
rect 0 514 2 522
rect 10 516 590 522
rect 598 516 600 524
rect 10 514 600 516
rect 0 510 600 514
rect 0 502 214 510
rect 248 502 600 510
rect 0 494 34 502
rect 72 494 106 502
rect 0 492 214 494
rect 222 484 240 494
rect 248 494 389 502
rect 457 494 527 502
rect 575 494 600 502
rect 248 492 600 494
rect 86 476 527 484
rect 78 472 86 476
rect 527 472 535 476
rect 0 456 70 460
rect 108 458 128 466
rect 136 458 158 466
rect 166 458 188 466
rect 196 458 218 466
rect 226 458 384 466
rect 392 458 414 466
rect 422 458 444 466
rect 452 458 474 466
rect 482 458 492 466
rect 108 456 296 458
rect 0 454 296 456
rect 0 446 34 454
rect 52 452 128 454
rect 52 446 64 452
rect 0 444 64 446
rect 72 446 128 452
rect 136 446 158 454
rect 166 446 188 454
rect 196 446 218 454
rect 226 450 296 454
rect 304 456 492 458
rect 542 459 600 460
rect 542 456 564 459
rect 304 454 564 456
rect 304 450 384 454
rect 226 446 384 450
rect 392 446 414 454
rect 422 446 444 454
rect 452 446 474 454
rect 482 451 564 454
rect 482 446 542 451
rect 72 444 542 446
rect 0 443 542 444
rect 560 443 564 451
rect 0 429 564 443
rect 0 421 108 429
rect 236 428 364 429
rect 236 421 296 428
rect 0 420 296 421
rect 304 421 364 428
rect 492 421 564 429
rect 304 420 564 421
rect 0 414 564 420
rect 0 406 34 414
rect 52 411 564 414
rect 52 406 542 411
rect 0 403 542 406
rect 560 403 564 411
rect 0 398 564 403
rect 0 390 296 398
rect 304 390 564 398
rect 0 374 564 390
rect 0 366 34 374
rect 52 371 564 374
rect 52 368 542 371
rect 52 366 296 368
rect 0 362 296 366
rect 0 354 112 362
rect 240 360 296 362
rect 304 363 542 368
rect 560 363 564 371
rect 304 362 564 363
rect 304 360 364 362
rect 240 354 364 360
rect 492 354 564 362
rect 0 338 564 354
rect 0 334 296 338
rect 0 326 34 334
rect 52 326 130 334
rect 138 326 160 334
rect 168 326 190 334
rect 198 326 220 334
rect 228 330 296 334
rect 304 335 564 338
rect 304 330 383 335
rect 228 327 383 330
rect 391 327 413 335
rect 421 327 443 335
rect 451 327 473 335
rect 481 331 564 335
rect 481 327 542 331
rect 228 326 542 327
rect 0 323 542 326
rect 560 323 564 331
rect 0 322 383 323
rect 0 314 130 322
rect 138 314 160 322
rect 168 314 190 322
rect 198 314 220 322
rect 228 315 383 322
rect 391 315 413 323
rect 421 315 443 323
rect 451 315 473 323
rect 481 315 564 323
rect 228 314 564 315
rect 0 310 564 314
rect 0 300 100 310
rect 286 308 314 310
rect 286 300 296 308
rect 304 300 314 308
rect 500 300 564 310
rect 0 296 564 300
rect 0 294 110 296
rect 0 286 34 294
rect 52 288 110 294
rect 238 288 363 296
rect 491 291 564 296
rect 491 288 542 291
rect 52 286 542 288
rect 0 283 542 286
rect 560 283 564 291
rect 0 278 564 283
rect 0 270 296 278
rect 304 270 564 278
rect 0 254 564 270
rect 0 246 34 254
rect 52 251 564 254
rect 52 248 542 251
rect 52 246 296 248
rect 0 240 296 246
rect 304 243 542 248
rect 560 243 564 251
rect 304 240 564 243
rect 0 232 564 240
rect 0 224 110 232
rect 238 231 564 232
rect 238 224 364 231
rect 0 223 364 224
rect 492 223 564 231
rect 0 218 564 223
rect 0 214 296 218
rect 0 206 34 214
rect 52 210 296 214
rect 304 211 564 218
rect 304 210 542 211
rect 52 206 542 210
rect 0 204 542 206
rect 0 196 129 204
rect 137 196 159 204
rect 167 196 189 204
rect 197 196 219 204
rect 227 196 384 204
rect 392 196 414 204
rect 422 196 444 204
rect 452 196 474 204
rect 482 203 542 204
rect 560 203 564 211
rect 482 196 564 203
rect 0 192 564 196
rect 0 184 129 192
rect 137 184 159 192
rect 167 184 189 192
rect 197 184 219 192
rect 227 188 384 192
rect 227 184 296 188
rect 0 180 296 184
rect 304 184 384 188
rect 392 184 414 192
rect 422 184 444 192
rect 452 184 474 192
rect 482 184 564 192
rect 304 180 564 184
rect 0 174 564 180
rect 0 166 34 174
rect 52 171 564 174
rect 52 168 542 171
rect 52 166 110 168
rect 0 160 110 166
rect 238 160 364 168
rect 492 163 542 168
rect 560 163 564 171
rect 492 160 564 163
rect 0 150 100 160
rect 286 158 314 160
rect 286 150 296 158
rect 304 150 314 158
rect 500 150 564 160
rect 0 134 564 150
rect 0 126 34 134
rect 52 131 564 134
rect 52 128 542 131
rect 52 126 296 128
rect 0 120 296 126
rect 304 123 542 128
rect 560 123 564 131
rect 304 120 564 123
rect 0 103 564 120
rect 0 102 364 103
rect 0 94 108 102
rect 236 95 364 102
rect 492 95 564 103
rect 236 94 564 95
rect 0 86 34 94
rect 52 91 564 94
rect 52 86 542 91
rect 0 83 542 86
rect 560 83 564 91
rect 0 73 564 83
rect 0 72 528 73
rect 0 64 64 72
rect 72 65 528 72
rect 536 65 564 73
rect 72 64 564 65
rect 0 62 474 64
rect 0 54 118 62
rect 0 48 78 54
rect 0 40 34 48
rect 42 40 48 48
rect 86 46 118 54
rect 76 40 118 46
rect 0 38 118 40
rect 0 0 14 38
rect 22 0 40 18
rect 48 0 80 38
rect 114 34 118 38
rect 126 34 138 62
rect 146 34 158 62
rect 166 34 178 62
rect 186 34 198 62
rect 206 34 218 62
rect 226 47 374 62
rect 226 34 246 47
rect 88 0 106 18
rect 114 0 246 34
rect 256 38 344 39
rect 256 0 344 30
rect 352 34 374 47
rect 382 34 394 62
rect 402 34 414 62
rect 422 34 434 62
rect 442 34 454 62
rect 462 36 474 62
rect 482 48 564 64
rect 482 40 536 48
rect 544 40 552 48
rect 560 40 564 48
rect 482 36 564 40
rect 462 35 564 36
rect 462 34 480 35
rect 352 0 480 34
rect 540 31 564 35
rect 572 31 600 459
rect 488 0 506 18
rect 514 0 532 18
rect 540 0 600 31
use PadBox  PadBox_0
timestamp 1570494029
transform 1 0 40 0 1 1480
box 0 0 520 520
<< labels >>
flabel nwell 600 -6 600 -6 6 FreeSans 16 0 0 0 VddNW
flabel nwell 0 -6 0 -6 4 FreeSans 16 0 0 0 VddNW
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 VddAct
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 VddAct
flabel psubstratepdiff 0 686 0 686 4 FreeSans 16 0 0 0 GndAct
flabel psubstratepdiff 600 686 600 686 6 FreeSans 16 0 0 0 GndAct
flabel metal1 466 682 466 682 4 FreeSans 64 0 0 0 DIunbuf
flabel metal1 434 682 434 682 6 FreeSans 64 0 0 0 DIB
flabel metal1 530 682 530 682 4 FreeSans 64 0 0 0 DI
flabel space 30 682 30 682 6 FreeSans 50 0 0 0 OEN
flabel metal1 54 682 54 682 6 FreeSans 50 0 0 0 OEB
flabel metal1 68 666 68 666 2 FreeSans 50 0 0 0 OE
flabel metal2 88 0 88 0 2 FreeSans 64 0 0 0 DO
flabel metal2 256 0 256 0 2 FreeSans 64 0 0 0 DATA
flabel metal2 22 0 22 0 4 FreeSans 64 0 0 0 OEN
flabel metal2 514 0 514 0 2 FreeSans 64 0 0 0 DI
flabel metal2 488 0 488 0 8 FreeSans 64 0 0 0 DIB
flabel metal2 256 0 256 0 4 FreeSans 64 0 0 0 DATA
flabel metal2 514 0 514 0 6 FreeSans 64 0 0 0 DI
flabel metal2 488 0 488 0 6 FreeSans 64 0 0 0 DIB
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 688 600 688 6 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 688 0 688 4 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 880 0 880 4 FreeSans 16 0 0 0 VddM2A
flabel metal2 600 880 600 880 6 FreeSans 16 0 0 0 VddM2A
flabel metal2 0 492 0 492 4 FreeSans 16 0 0 0 VddM2B
flabel metal2 600 492 600 492 6 FreeSans 16 0 0 0 VddM2B
flabel metal2 88 0 88 0 4 FreeSans 52 0 0 0 DO
<< properties >>
string path 1278.000 4630.500 1422.000 4630.500 1422.000 5539.500 1278.000 5539.500 1278.000 4630.500 
<< end >>
