../../lef/amic5n_std_cell.lef