`celldefine
module inv_d (z, a);
  output z;
  input  a;

  not G1 (z, a);
endmodule
`endcelldefine
