magic
tech scmos
timestamp 1592705592
<< nwell >>
rect 14 541 346 770
rect -3 507 363 524
rect -3 462 363 479
rect -3 233 14 462
rect 346 233 363 462
rect -3 216 363 233
rect 12 1 19 53
rect 341 1 348 53
<< ntransistor >>
rect 38 433 159 436
rect 38 389 159 392
rect 38 368 159 371
rect 38 324 159 327
rect 38 303 159 306
rect 38 259 159 262
rect 201 433 322 436
rect 201 389 322 392
rect 201 368 322 371
rect 201 324 322 327
rect 201 303 322 306
rect 201 259 322 262
<< ptransistor >>
rect 38 741 166 744
rect 38 697 166 700
rect 38 676 166 679
rect 38 632 166 635
rect 38 611 166 614
rect 38 567 166 570
rect 194 741 322 744
rect 194 697 322 700
rect 194 676 322 679
rect 194 632 322 635
rect 194 611 322 614
rect 194 567 322 570
<< ndiffusion >>
rect 36 439 161 445
rect 199 439 324 445
rect 38 436 159 439
rect 38 392 159 433
rect 38 371 159 389
rect 38 327 159 368
rect 38 306 159 324
rect 38 262 159 303
rect 38 256 159 259
rect 201 436 322 439
rect 201 392 322 433
rect 201 371 322 389
rect 201 327 322 368
rect 201 306 322 324
rect 201 262 322 303
rect 201 256 322 259
rect 36 250 161 256
rect 199 250 324 256
<< pdiffusion >>
rect 36 747 168 753
rect 192 747 324 753
rect 38 744 166 747
rect 38 700 166 741
rect 38 679 166 697
rect 38 635 166 676
rect 38 614 166 632
rect 38 570 166 611
rect 38 564 166 567
rect 194 744 322 747
rect 194 700 322 741
rect 194 679 322 697
rect 194 635 322 676
rect 194 614 322 632
rect 194 570 322 611
rect 194 564 322 567
rect 36 558 168 564
rect 192 558 324 564
<< psubstratepdiff >>
rect 0 773 360 784
rect 0 538 11 773
rect 349 538 360 773
rect 0 527 360 538
rect 0 482 360 493
rect 19 445 341 457
rect 19 439 36 445
rect 161 439 199 445
rect 324 439 341 445
rect 19 256 30 439
rect 167 256 193 439
rect 330 256 341 439
rect 19 250 36 256
rect 161 250 199 256
rect 324 250 341 256
rect 19 238 341 250
rect 0 202 360 213
rect 0 100 11 202
rect 349 100 360 202
rect 0 89 360 100
<< nsubstratendiff >>
rect 19 753 341 765
rect 19 747 36 753
rect 168 747 192 753
rect 324 747 341 753
rect 19 564 30 747
rect 174 564 186 747
rect 330 564 341 747
rect 19 558 36 564
rect 168 558 192 564
rect 324 558 341 564
rect 19 546 341 558
rect 0 510 360 521
rect 0 465 360 476
rect 0 230 11 465
rect 349 230 360 465
rect 0 219 360 230
rect 81 160 279 171
rect 81 125 279 136
<< polysilicon >>
rect 31 741 38 744
rect 166 741 173 744
rect 31 700 37 741
rect 167 700 173 741
rect 31 697 38 700
rect 166 697 173 700
rect 31 679 37 697
rect 167 679 173 697
rect 31 676 38 679
rect 166 676 173 679
rect 31 635 37 676
rect 167 635 173 676
rect 31 632 38 635
rect 166 632 173 635
rect 31 614 37 632
rect 167 614 173 632
rect 31 611 38 614
rect 166 611 173 614
rect 31 570 37 611
rect 167 570 173 611
rect 31 567 38 570
rect 166 567 173 570
rect 187 741 194 744
rect 322 741 329 744
rect 187 700 193 741
rect 323 700 329 741
rect 187 697 194 700
rect 322 697 329 700
rect 187 679 193 697
rect 323 679 329 697
rect 187 676 194 679
rect 322 676 329 679
rect 187 635 193 676
rect 323 635 329 676
rect 187 632 194 635
rect 322 632 329 635
rect 187 614 193 632
rect 323 614 329 632
rect 187 611 194 614
rect 322 611 329 614
rect 187 570 193 611
rect 323 570 329 611
rect 187 567 194 570
rect 322 567 329 570
rect 31 433 38 436
rect 159 433 166 436
rect 31 392 37 433
rect 160 392 166 433
rect 31 389 38 392
rect 159 389 166 392
rect 31 371 37 389
rect 160 371 166 389
rect 31 368 38 371
rect 159 368 166 371
rect 31 327 37 368
rect 160 327 166 368
rect 31 324 38 327
rect 159 324 166 327
rect 31 306 37 324
rect 160 306 166 324
rect 31 303 38 306
rect 159 303 166 306
rect 31 262 37 303
rect 160 262 166 303
rect 31 259 38 262
rect 159 259 166 262
rect 194 433 201 436
rect 322 433 329 436
rect 194 392 200 433
rect 323 392 329 433
rect 194 389 201 392
rect 322 389 329 392
rect 194 371 200 389
rect 323 371 329 389
rect 194 368 201 371
rect 322 368 329 371
rect 194 327 200 368
rect 323 327 329 368
rect 194 324 201 327
rect 322 324 329 327
rect 194 306 200 324
rect 323 306 329 324
rect 194 303 201 306
rect 322 303 329 306
rect 194 262 200 303
rect 323 262 329 303
rect 194 259 201 262
rect 322 259 329 262
<< genericcontact >>
rect 9 780 11 782
rect 17 780 19 782
rect 25 780 27 782
rect 33 780 35 782
rect 41 780 43 782
rect 49 780 51 782
rect 57 780 59 782
rect 65 780 67 782
rect 73 780 75 782
rect 81 780 83 782
rect 89 780 91 782
rect 97 780 99 782
rect 105 780 107 782
rect 113 780 115 782
rect 151 780 153 782
rect 159 780 161 782
rect 167 780 169 782
rect 175 780 177 782
rect 183 780 185 782
rect 191 780 193 782
rect 199 780 201 782
rect 207 780 209 782
rect 245 780 247 782
rect 253 780 255 782
rect 261 780 263 782
rect 269 780 271 782
rect 277 780 279 782
rect 285 780 287 782
rect 293 780 295 782
rect 301 780 303 782
rect 309 780 311 782
rect 317 780 319 782
rect 325 780 327 782
rect 333 780 335 782
rect 341 780 343 782
rect 349 780 351 782
rect 9 775 11 777
rect 17 775 19 777
rect 25 775 27 777
rect 33 775 35 777
rect 41 775 43 777
rect 49 775 51 777
rect 57 775 59 777
rect 65 775 67 777
rect 73 775 75 777
rect 81 775 83 777
rect 89 775 91 777
rect 97 775 99 777
rect 105 775 107 777
rect 113 775 115 777
rect 151 775 153 777
rect 159 775 161 777
rect 167 775 169 777
rect 175 775 177 777
rect 183 775 185 777
rect 191 775 193 777
rect 199 775 201 777
rect 207 775 209 777
rect 245 775 247 777
rect 253 775 255 777
rect 261 775 263 777
rect 269 775 271 777
rect 277 775 279 777
rect 285 775 287 777
rect 293 775 295 777
rect 301 775 303 777
rect 309 775 311 777
rect 317 775 319 777
rect 325 775 327 777
rect 333 775 335 777
rect 341 775 343 777
rect 349 775 351 777
rect 2 767 4 769
rect 7 767 9 769
rect 351 767 353 769
rect 356 767 358 769
rect 2 759 4 761
rect 7 759 9 761
rect 351 759 353 761
rect 356 759 358 761
rect 30 757 32 759
rect 41 757 43 759
rect 51 757 53 759
rect 61 757 63 759
rect 71 757 73 759
rect 81 757 83 759
rect 91 757 93 759
rect 101 757 103 759
rect 111 757 113 759
rect 150 757 152 759
rect 160 757 162 759
rect 198 757 200 759
rect 208 757 210 759
rect 247 757 249 759
rect 257 757 259 759
rect 267 757 269 759
rect 277 757 279 759
rect 287 757 289 759
rect 297 757 299 759
rect 307 757 309 759
rect 317 757 319 759
rect 327 757 329 759
rect 2 751 4 753
rect 7 751 9 753
rect 30 752 32 754
rect 41 752 43 754
rect 51 752 53 754
rect 61 752 63 754
rect 71 752 73 754
rect 81 752 83 754
rect 91 752 93 754
rect 101 752 103 754
rect 111 752 113 754
rect 150 752 152 754
rect 160 752 162 754
rect 198 752 200 754
rect 208 752 210 754
rect 247 752 249 754
rect 257 752 259 754
rect 267 752 269 754
rect 277 752 279 754
rect 287 752 289 754
rect 297 752 299 754
rect 307 752 309 754
rect 317 752 319 754
rect 327 752 329 754
rect 351 751 353 753
rect 356 751 358 753
rect 41 747 43 749
rect 51 747 53 749
rect 61 747 63 749
rect 71 747 73 749
rect 81 747 83 749
rect 91 747 93 749
rect 101 747 103 749
rect 111 747 113 749
rect 150 747 152 749
rect 160 747 162 749
rect 198 747 200 749
rect 208 747 210 749
rect 247 747 249 749
rect 257 747 259 749
rect 267 747 269 749
rect 277 747 279 749
rect 287 747 289 749
rect 297 747 299 749
rect 307 747 309 749
rect 317 747 319 749
rect 2 743 4 745
rect 7 743 9 745
rect 20 742 22 744
rect 25 742 27 744
rect 177 742 179 744
rect 182 742 184 744
rect 333 742 335 744
rect 338 742 340 744
rect 351 743 353 745
rect 356 743 358 745
rect 33 739 35 741
rect 169 739 171 741
rect 189 739 191 741
rect 325 739 327 741
rect 20 737 22 739
rect 25 737 27 739
rect 42 737 44 739
rect 47 737 49 739
rect 52 737 54 739
rect 57 737 59 739
rect 62 737 64 739
rect 67 737 69 739
rect 72 737 74 739
rect 77 737 79 739
rect 82 737 84 739
rect 87 737 89 739
rect 92 737 94 739
rect 97 737 99 739
rect 102 737 104 739
rect 107 737 109 739
rect 112 737 114 739
rect 117 737 119 739
rect 122 737 124 739
rect 127 737 129 739
rect 132 737 134 739
rect 137 737 139 739
rect 142 737 144 739
rect 147 737 149 739
rect 152 737 154 739
rect 157 737 159 739
rect 162 737 164 739
rect 177 737 179 739
rect 182 737 184 739
rect 196 737 198 739
rect 201 737 203 739
rect 206 737 208 739
rect 211 737 213 739
rect 216 737 218 739
rect 221 737 223 739
rect 226 737 228 739
rect 231 737 233 739
rect 236 737 238 739
rect 241 737 243 739
rect 246 737 248 739
rect 251 737 253 739
rect 256 737 258 739
rect 261 737 263 739
rect 266 737 268 739
rect 271 737 273 739
rect 276 737 278 739
rect 281 737 283 739
rect 286 737 288 739
rect 291 737 293 739
rect 296 737 298 739
rect 301 737 303 739
rect 306 737 308 739
rect 311 737 313 739
rect 316 737 318 739
rect 333 737 335 739
rect 338 737 340 739
rect 2 735 4 737
rect 7 735 9 737
rect 33 734 35 736
rect 169 734 171 736
rect 189 734 191 736
rect 325 734 327 736
rect 351 735 353 737
rect 356 735 358 737
rect 20 732 22 734
rect 25 732 27 734
rect 42 732 44 734
rect 47 732 49 734
rect 52 732 54 734
rect 57 732 59 734
rect 62 732 64 734
rect 67 732 69 734
rect 72 732 74 734
rect 77 732 79 734
rect 82 732 84 734
rect 87 732 89 734
rect 92 732 94 734
rect 97 732 99 734
rect 102 732 104 734
rect 107 732 109 734
rect 112 732 114 734
rect 117 732 119 734
rect 122 732 124 734
rect 127 732 129 734
rect 132 732 134 734
rect 137 732 139 734
rect 142 732 144 734
rect 147 732 149 734
rect 152 732 154 734
rect 157 732 159 734
rect 162 732 164 734
rect 177 732 179 734
rect 182 732 184 734
rect 196 732 198 734
rect 201 732 203 734
rect 206 732 208 734
rect 211 732 213 734
rect 216 732 218 734
rect 221 732 223 734
rect 226 732 228 734
rect 231 732 233 734
rect 236 732 238 734
rect 241 732 243 734
rect 246 732 248 734
rect 251 732 253 734
rect 256 732 258 734
rect 261 732 263 734
rect 266 732 268 734
rect 271 732 273 734
rect 276 732 278 734
rect 281 732 283 734
rect 286 732 288 734
rect 291 732 293 734
rect 296 732 298 734
rect 301 732 303 734
rect 306 732 308 734
rect 311 732 313 734
rect 316 732 318 734
rect 333 732 335 734
rect 338 732 340 734
rect 33 729 35 731
rect 169 729 171 731
rect 189 729 191 731
rect 325 729 327 731
rect 2 727 4 729
rect 7 727 9 729
rect 20 727 22 729
rect 25 727 27 729
rect 42 727 44 729
rect 47 727 49 729
rect 52 727 54 729
rect 57 727 59 729
rect 62 727 64 729
rect 67 727 69 729
rect 72 727 74 729
rect 77 727 79 729
rect 82 727 84 729
rect 87 727 89 729
rect 92 727 94 729
rect 97 727 99 729
rect 102 727 104 729
rect 107 727 109 729
rect 112 727 114 729
rect 117 727 119 729
rect 122 727 124 729
rect 127 727 129 729
rect 132 727 134 729
rect 137 727 139 729
rect 142 727 144 729
rect 147 727 149 729
rect 152 727 154 729
rect 157 727 159 729
rect 162 727 164 729
rect 177 727 179 729
rect 182 727 184 729
rect 196 727 198 729
rect 201 727 203 729
rect 206 727 208 729
rect 211 727 213 729
rect 216 727 218 729
rect 221 727 223 729
rect 226 727 228 729
rect 231 727 233 729
rect 236 727 238 729
rect 241 727 243 729
rect 246 727 248 729
rect 251 727 253 729
rect 256 727 258 729
rect 261 727 263 729
rect 266 727 268 729
rect 271 727 273 729
rect 276 727 278 729
rect 281 727 283 729
rect 286 727 288 729
rect 291 727 293 729
rect 296 727 298 729
rect 301 727 303 729
rect 306 727 308 729
rect 311 727 313 729
rect 316 727 318 729
rect 333 727 335 729
rect 338 727 340 729
rect 351 727 353 729
rect 356 727 358 729
rect 33 724 35 726
rect 169 724 171 726
rect 189 724 191 726
rect 325 724 327 726
rect 20 722 22 724
rect 25 722 27 724
rect 42 722 44 724
rect 47 722 49 724
rect 52 722 54 724
rect 57 722 59 724
rect 62 722 64 724
rect 67 722 69 724
rect 72 722 74 724
rect 77 722 79 724
rect 82 722 84 724
rect 87 722 89 724
rect 92 722 94 724
rect 97 722 99 724
rect 102 722 104 724
rect 107 722 109 724
rect 112 722 114 724
rect 117 722 119 724
rect 122 722 124 724
rect 127 722 129 724
rect 132 722 134 724
rect 137 722 139 724
rect 142 722 144 724
rect 147 722 149 724
rect 152 722 154 724
rect 157 722 159 724
rect 162 722 164 724
rect 177 722 179 724
rect 182 722 184 724
rect 196 722 198 724
rect 201 722 203 724
rect 206 722 208 724
rect 211 722 213 724
rect 216 722 218 724
rect 221 722 223 724
rect 226 722 228 724
rect 231 722 233 724
rect 236 722 238 724
rect 241 722 243 724
rect 246 722 248 724
rect 251 722 253 724
rect 256 722 258 724
rect 261 722 263 724
rect 266 722 268 724
rect 271 722 273 724
rect 276 722 278 724
rect 281 722 283 724
rect 286 722 288 724
rect 291 722 293 724
rect 296 722 298 724
rect 301 722 303 724
rect 306 722 308 724
rect 311 722 313 724
rect 316 722 318 724
rect 333 722 335 724
rect 338 722 340 724
rect 2 719 4 721
rect 7 719 9 721
rect 33 719 35 721
rect 169 719 171 721
rect 189 719 191 721
rect 325 719 327 721
rect 351 719 353 721
rect 356 719 358 721
rect 20 717 22 719
rect 25 717 27 719
rect 42 717 44 719
rect 47 717 49 719
rect 52 717 54 719
rect 57 717 59 719
rect 62 717 64 719
rect 67 717 69 719
rect 72 717 74 719
rect 77 717 79 719
rect 82 717 84 719
rect 87 717 89 719
rect 92 717 94 719
rect 97 717 99 719
rect 102 717 104 719
rect 107 717 109 719
rect 112 717 114 719
rect 117 717 119 719
rect 122 717 124 719
rect 127 717 129 719
rect 132 717 134 719
rect 137 717 139 719
rect 142 717 144 719
rect 147 717 149 719
rect 152 717 154 719
rect 157 717 159 719
rect 162 717 164 719
rect 177 717 179 719
rect 182 717 184 719
rect 196 717 198 719
rect 201 717 203 719
rect 206 717 208 719
rect 211 717 213 719
rect 216 717 218 719
rect 221 717 223 719
rect 226 717 228 719
rect 231 717 233 719
rect 236 717 238 719
rect 241 717 243 719
rect 246 717 248 719
rect 251 717 253 719
rect 256 717 258 719
rect 261 717 263 719
rect 266 717 268 719
rect 271 717 273 719
rect 276 717 278 719
rect 281 717 283 719
rect 286 717 288 719
rect 291 717 293 719
rect 296 717 298 719
rect 301 717 303 719
rect 306 717 308 719
rect 311 717 313 719
rect 316 717 318 719
rect 333 717 335 719
rect 338 717 340 719
rect 33 714 35 716
rect 169 714 171 716
rect 189 714 191 716
rect 325 714 327 716
rect 2 711 4 713
rect 7 711 9 713
rect 20 712 22 714
rect 25 712 27 714
rect 42 712 44 714
rect 47 712 49 714
rect 52 712 54 714
rect 57 712 59 714
rect 62 712 64 714
rect 67 712 69 714
rect 72 712 74 714
rect 77 712 79 714
rect 82 712 84 714
rect 87 712 89 714
rect 92 712 94 714
rect 97 712 99 714
rect 102 712 104 714
rect 107 712 109 714
rect 112 712 114 714
rect 117 712 119 714
rect 122 712 124 714
rect 127 712 129 714
rect 132 712 134 714
rect 137 712 139 714
rect 142 712 144 714
rect 147 712 149 714
rect 152 712 154 714
rect 157 712 159 714
rect 162 712 164 714
rect 177 712 179 714
rect 182 712 184 714
rect 196 712 198 714
rect 201 712 203 714
rect 206 712 208 714
rect 211 712 213 714
rect 216 712 218 714
rect 221 712 223 714
rect 226 712 228 714
rect 231 712 233 714
rect 236 712 238 714
rect 241 712 243 714
rect 246 712 248 714
rect 251 712 253 714
rect 256 712 258 714
rect 261 712 263 714
rect 266 712 268 714
rect 271 712 273 714
rect 276 712 278 714
rect 281 712 283 714
rect 286 712 288 714
rect 291 712 293 714
rect 296 712 298 714
rect 301 712 303 714
rect 306 712 308 714
rect 311 712 313 714
rect 316 712 318 714
rect 333 712 335 714
rect 338 712 340 714
rect 351 711 353 713
rect 356 711 358 713
rect 33 709 35 711
rect 169 709 171 711
rect 189 709 191 711
rect 325 709 327 711
rect 20 707 22 709
rect 25 707 27 709
rect 42 707 44 709
rect 47 707 49 709
rect 52 707 54 709
rect 57 707 59 709
rect 62 707 64 709
rect 67 707 69 709
rect 72 707 74 709
rect 77 707 79 709
rect 82 707 84 709
rect 87 707 89 709
rect 92 707 94 709
rect 97 707 99 709
rect 102 707 104 709
rect 107 707 109 709
rect 112 707 114 709
rect 117 707 119 709
rect 122 707 124 709
rect 127 707 129 709
rect 132 707 134 709
rect 137 707 139 709
rect 142 707 144 709
rect 147 707 149 709
rect 152 707 154 709
rect 157 707 159 709
rect 162 707 164 709
rect 177 707 179 709
rect 182 707 184 709
rect 196 707 198 709
rect 201 707 203 709
rect 206 707 208 709
rect 211 707 213 709
rect 216 707 218 709
rect 221 707 223 709
rect 226 707 228 709
rect 231 707 233 709
rect 236 707 238 709
rect 241 707 243 709
rect 246 707 248 709
rect 251 707 253 709
rect 256 707 258 709
rect 261 707 263 709
rect 266 707 268 709
rect 271 707 273 709
rect 276 707 278 709
rect 281 707 283 709
rect 286 707 288 709
rect 291 707 293 709
rect 296 707 298 709
rect 301 707 303 709
rect 306 707 308 709
rect 311 707 313 709
rect 316 707 318 709
rect 333 707 335 709
rect 338 707 340 709
rect 2 703 4 705
rect 7 703 9 705
rect 33 704 35 706
rect 169 704 171 706
rect 189 704 191 706
rect 325 704 327 706
rect 20 702 22 704
rect 25 702 27 704
rect 42 702 44 704
rect 47 702 49 704
rect 52 702 54 704
rect 57 702 59 704
rect 62 702 64 704
rect 67 702 69 704
rect 72 702 74 704
rect 77 702 79 704
rect 82 702 84 704
rect 87 702 89 704
rect 92 702 94 704
rect 97 702 99 704
rect 102 702 104 704
rect 107 702 109 704
rect 112 702 114 704
rect 117 702 119 704
rect 122 702 124 704
rect 127 702 129 704
rect 132 702 134 704
rect 137 702 139 704
rect 142 702 144 704
rect 147 702 149 704
rect 152 702 154 704
rect 157 702 159 704
rect 162 702 164 704
rect 177 702 179 704
rect 182 702 184 704
rect 196 702 198 704
rect 201 702 203 704
rect 206 702 208 704
rect 211 702 213 704
rect 216 702 218 704
rect 221 702 223 704
rect 226 702 228 704
rect 231 702 233 704
rect 236 702 238 704
rect 241 702 243 704
rect 246 702 248 704
rect 251 702 253 704
rect 256 702 258 704
rect 261 702 263 704
rect 266 702 268 704
rect 271 702 273 704
rect 276 702 278 704
rect 281 702 283 704
rect 286 702 288 704
rect 291 702 293 704
rect 296 702 298 704
rect 301 702 303 704
rect 306 702 308 704
rect 311 702 313 704
rect 316 702 318 704
rect 333 702 335 704
rect 338 702 340 704
rect 351 703 353 705
rect 356 703 358 705
rect 33 699 35 701
rect 169 699 171 701
rect 189 699 191 701
rect 325 699 327 701
rect 20 697 22 699
rect 25 697 27 699
rect 177 697 179 699
rect 182 697 184 699
rect 333 697 335 699
rect 338 697 340 699
rect 2 695 4 697
rect 7 695 9 697
rect 33 694 35 696
rect 169 694 171 696
rect 189 694 191 696
rect 325 694 327 696
rect 351 695 353 697
rect 356 695 358 697
rect 41 692 43 694
rect 51 692 53 694
rect 61 692 63 694
rect 71 692 73 694
rect 81 692 83 694
rect 91 692 93 694
rect 101 692 103 694
rect 111 692 113 694
rect 150 692 152 694
rect 160 692 162 694
rect 198 692 200 694
rect 208 692 210 694
rect 247 692 249 694
rect 257 692 259 694
rect 267 692 269 694
rect 277 692 279 694
rect 287 692 289 694
rect 297 692 299 694
rect 307 692 309 694
rect 317 692 319 694
rect 33 689 35 691
rect 169 689 171 691
rect 189 689 191 691
rect 325 689 327 691
rect 2 687 4 689
rect 7 687 9 689
rect 41 687 43 689
rect 51 687 53 689
rect 61 687 63 689
rect 71 687 73 689
rect 81 687 83 689
rect 91 687 93 689
rect 101 687 103 689
rect 111 687 113 689
rect 150 687 152 689
rect 160 687 162 689
rect 198 687 200 689
rect 208 687 210 689
rect 247 687 249 689
rect 257 687 259 689
rect 267 687 269 689
rect 277 687 279 689
rect 287 687 289 689
rect 297 687 299 689
rect 307 687 309 689
rect 317 687 319 689
rect 351 687 353 689
rect 356 687 358 689
rect 33 684 35 686
rect 169 684 171 686
rect 189 684 191 686
rect 325 684 327 686
rect 41 682 43 684
rect 51 682 53 684
rect 61 682 63 684
rect 71 682 73 684
rect 81 682 83 684
rect 91 682 93 684
rect 101 682 103 684
rect 111 682 113 684
rect 150 682 152 684
rect 160 682 162 684
rect 198 682 200 684
rect 208 682 210 684
rect 247 682 249 684
rect 257 682 259 684
rect 267 682 269 684
rect 277 682 279 684
rect 287 682 289 684
rect 297 682 299 684
rect 307 682 309 684
rect 317 682 319 684
rect 2 679 4 681
rect 7 679 9 681
rect 33 679 35 681
rect 169 679 171 681
rect 189 679 191 681
rect 325 679 327 681
rect 351 679 353 681
rect 356 679 358 681
rect 20 677 22 679
rect 25 677 27 679
rect 177 677 179 679
rect 182 677 184 679
rect 333 677 335 679
rect 338 677 340 679
rect 33 674 35 676
rect 169 674 171 676
rect 189 674 191 676
rect 325 674 327 676
rect 2 671 4 673
rect 7 671 9 673
rect 20 672 22 674
rect 25 672 27 674
rect 42 672 44 674
rect 47 672 49 674
rect 52 672 54 674
rect 57 672 59 674
rect 62 672 64 674
rect 67 672 69 674
rect 72 672 74 674
rect 77 672 79 674
rect 82 672 84 674
rect 87 672 89 674
rect 92 672 94 674
rect 97 672 99 674
rect 102 672 104 674
rect 107 672 109 674
rect 112 672 114 674
rect 117 672 119 674
rect 122 672 124 674
rect 127 672 129 674
rect 132 672 134 674
rect 137 672 139 674
rect 142 672 144 674
rect 147 672 149 674
rect 152 672 154 674
rect 157 672 159 674
rect 162 672 164 674
rect 177 672 179 674
rect 182 672 184 674
rect 196 672 198 674
rect 201 672 203 674
rect 206 672 208 674
rect 211 672 213 674
rect 216 672 218 674
rect 221 672 223 674
rect 226 672 228 674
rect 231 672 233 674
rect 236 672 238 674
rect 241 672 243 674
rect 246 672 248 674
rect 251 672 253 674
rect 256 672 258 674
rect 261 672 263 674
rect 266 672 268 674
rect 271 672 273 674
rect 276 672 278 674
rect 281 672 283 674
rect 286 672 288 674
rect 291 672 293 674
rect 296 672 298 674
rect 301 672 303 674
rect 306 672 308 674
rect 311 672 313 674
rect 316 672 318 674
rect 333 672 335 674
rect 338 672 340 674
rect 351 671 353 673
rect 356 671 358 673
rect 33 669 35 671
rect 169 669 171 671
rect 189 669 191 671
rect 325 669 327 671
rect 20 667 22 669
rect 25 667 27 669
rect 42 667 44 669
rect 47 667 49 669
rect 52 667 54 669
rect 57 667 59 669
rect 62 667 64 669
rect 67 667 69 669
rect 72 667 74 669
rect 77 667 79 669
rect 82 667 84 669
rect 87 667 89 669
rect 92 667 94 669
rect 97 667 99 669
rect 102 667 104 669
rect 107 667 109 669
rect 112 667 114 669
rect 117 667 119 669
rect 122 667 124 669
rect 127 667 129 669
rect 132 667 134 669
rect 137 667 139 669
rect 142 667 144 669
rect 147 667 149 669
rect 152 667 154 669
rect 157 667 159 669
rect 162 667 164 669
rect 177 667 179 669
rect 182 667 184 669
rect 196 667 198 669
rect 201 667 203 669
rect 206 667 208 669
rect 211 667 213 669
rect 216 667 218 669
rect 221 667 223 669
rect 226 667 228 669
rect 231 667 233 669
rect 236 667 238 669
rect 241 667 243 669
rect 246 667 248 669
rect 251 667 253 669
rect 256 667 258 669
rect 261 667 263 669
rect 266 667 268 669
rect 271 667 273 669
rect 276 667 278 669
rect 281 667 283 669
rect 286 667 288 669
rect 291 667 293 669
rect 296 667 298 669
rect 301 667 303 669
rect 306 667 308 669
rect 311 667 313 669
rect 316 667 318 669
rect 333 667 335 669
rect 338 667 340 669
rect 2 663 4 665
rect 7 663 9 665
rect 33 664 35 666
rect 169 664 171 666
rect 189 664 191 666
rect 325 664 327 666
rect 20 662 22 664
rect 25 662 27 664
rect 42 662 44 664
rect 47 662 49 664
rect 52 662 54 664
rect 57 662 59 664
rect 62 662 64 664
rect 67 662 69 664
rect 72 662 74 664
rect 77 662 79 664
rect 82 662 84 664
rect 87 662 89 664
rect 92 662 94 664
rect 97 662 99 664
rect 102 662 104 664
rect 107 662 109 664
rect 112 662 114 664
rect 117 662 119 664
rect 122 662 124 664
rect 127 662 129 664
rect 132 662 134 664
rect 137 662 139 664
rect 142 662 144 664
rect 147 662 149 664
rect 152 662 154 664
rect 157 662 159 664
rect 162 662 164 664
rect 177 662 179 664
rect 182 662 184 664
rect 196 662 198 664
rect 201 662 203 664
rect 206 662 208 664
rect 211 662 213 664
rect 216 662 218 664
rect 221 662 223 664
rect 226 662 228 664
rect 231 662 233 664
rect 236 662 238 664
rect 241 662 243 664
rect 246 662 248 664
rect 251 662 253 664
rect 256 662 258 664
rect 261 662 263 664
rect 266 662 268 664
rect 271 662 273 664
rect 276 662 278 664
rect 281 662 283 664
rect 286 662 288 664
rect 291 662 293 664
rect 296 662 298 664
rect 301 662 303 664
rect 306 662 308 664
rect 311 662 313 664
rect 316 662 318 664
rect 333 662 335 664
rect 338 662 340 664
rect 351 663 353 665
rect 356 663 358 665
rect 33 659 35 661
rect 169 659 171 661
rect 189 659 191 661
rect 325 659 327 661
rect 20 657 22 659
rect 25 657 27 659
rect 42 657 44 659
rect 47 657 49 659
rect 52 657 54 659
rect 57 657 59 659
rect 62 657 64 659
rect 67 657 69 659
rect 72 657 74 659
rect 77 657 79 659
rect 82 657 84 659
rect 87 657 89 659
rect 92 657 94 659
rect 97 657 99 659
rect 102 657 104 659
rect 107 657 109 659
rect 112 657 114 659
rect 117 657 119 659
rect 122 657 124 659
rect 127 657 129 659
rect 132 657 134 659
rect 137 657 139 659
rect 142 657 144 659
rect 147 657 149 659
rect 152 657 154 659
rect 157 657 159 659
rect 162 657 164 659
rect 177 657 179 659
rect 182 657 184 659
rect 196 657 198 659
rect 201 657 203 659
rect 206 657 208 659
rect 211 657 213 659
rect 216 657 218 659
rect 221 657 223 659
rect 226 657 228 659
rect 231 657 233 659
rect 236 657 238 659
rect 241 657 243 659
rect 246 657 248 659
rect 251 657 253 659
rect 256 657 258 659
rect 261 657 263 659
rect 266 657 268 659
rect 271 657 273 659
rect 276 657 278 659
rect 281 657 283 659
rect 286 657 288 659
rect 291 657 293 659
rect 296 657 298 659
rect 301 657 303 659
rect 306 657 308 659
rect 311 657 313 659
rect 316 657 318 659
rect 333 657 335 659
rect 338 657 340 659
rect 2 655 4 657
rect 7 655 9 657
rect 351 655 353 657
rect 356 655 358 657
rect 20 652 22 654
rect 25 652 27 654
rect 33 653 35 655
rect 42 652 44 654
rect 47 652 49 654
rect 52 652 54 654
rect 57 652 59 654
rect 62 652 64 654
rect 67 652 69 654
rect 72 652 74 654
rect 77 652 79 654
rect 82 652 84 654
rect 87 652 89 654
rect 92 652 94 654
rect 97 652 99 654
rect 102 652 104 654
rect 107 652 109 654
rect 112 652 114 654
rect 117 652 119 654
rect 122 652 124 654
rect 127 652 129 654
rect 132 652 134 654
rect 137 652 139 654
rect 142 652 144 654
rect 147 652 149 654
rect 152 652 154 654
rect 157 652 159 654
rect 162 652 164 654
rect 169 653 171 655
rect 177 652 179 654
rect 182 652 184 654
rect 189 653 191 655
rect 196 652 198 654
rect 201 652 203 654
rect 206 652 208 654
rect 211 652 213 654
rect 216 652 218 654
rect 221 652 223 654
rect 226 652 228 654
rect 231 652 233 654
rect 236 652 238 654
rect 241 652 243 654
rect 246 652 248 654
rect 251 652 253 654
rect 256 652 258 654
rect 261 652 263 654
rect 266 652 268 654
rect 271 652 273 654
rect 276 652 278 654
rect 281 652 283 654
rect 286 652 288 654
rect 291 652 293 654
rect 296 652 298 654
rect 301 652 303 654
rect 306 652 308 654
rect 311 652 313 654
rect 316 652 318 654
rect 325 653 327 655
rect 333 652 335 654
rect 338 652 340 654
rect 2 647 4 649
rect 7 647 9 649
rect 20 647 22 649
rect 25 647 27 649
rect 33 648 35 650
rect 42 647 44 649
rect 47 647 49 649
rect 52 647 54 649
rect 57 647 59 649
rect 62 647 64 649
rect 67 647 69 649
rect 72 647 74 649
rect 77 647 79 649
rect 82 647 84 649
rect 87 647 89 649
rect 92 647 94 649
rect 97 647 99 649
rect 102 647 104 649
rect 107 647 109 649
rect 112 647 114 649
rect 117 647 119 649
rect 122 647 124 649
rect 127 647 129 649
rect 132 647 134 649
rect 137 647 139 649
rect 142 647 144 649
rect 147 647 149 649
rect 152 647 154 649
rect 157 647 159 649
rect 162 647 164 649
rect 169 648 171 650
rect 177 647 179 649
rect 182 647 184 649
rect 189 648 191 650
rect 196 647 198 649
rect 201 647 203 649
rect 206 647 208 649
rect 211 647 213 649
rect 216 647 218 649
rect 221 647 223 649
rect 226 647 228 649
rect 231 647 233 649
rect 236 647 238 649
rect 241 647 243 649
rect 246 647 248 649
rect 251 647 253 649
rect 256 647 258 649
rect 261 647 263 649
rect 266 647 268 649
rect 271 647 273 649
rect 276 647 278 649
rect 281 647 283 649
rect 286 647 288 649
rect 291 647 293 649
rect 296 647 298 649
rect 301 647 303 649
rect 306 647 308 649
rect 311 647 313 649
rect 316 647 318 649
rect 325 648 327 650
rect 333 647 335 649
rect 338 647 340 649
rect 351 647 353 649
rect 356 647 358 649
rect 20 642 22 644
rect 25 642 27 644
rect 33 643 35 645
rect 42 642 44 644
rect 47 642 49 644
rect 52 642 54 644
rect 57 642 59 644
rect 62 642 64 644
rect 67 642 69 644
rect 72 642 74 644
rect 77 642 79 644
rect 82 642 84 644
rect 87 642 89 644
rect 92 642 94 644
rect 97 642 99 644
rect 102 642 104 644
rect 107 642 109 644
rect 112 642 114 644
rect 117 642 119 644
rect 122 642 124 644
rect 127 642 129 644
rect 132 642 134 644
rect 137 642 139 644
rect 142 642 144 644
rect 147 642 149 644
rect 152 642 154 644
rect 157 642 159 644
rect 162 642 164 644
rect 169 643 171 645
rect 177 642 179 644
rect 182 642 184 644
rect 189 643 191 645
rect 196 642 198 644
rect 201 642 203 644
rect 206 642 208 644
rect 211 642 213 644
rect 216 642 218 644
rect 221 642 223 644
rect 226 642 228 644
rect 231 642 233 644
rect 236 642 238 644
rect 241 642 243 644
rect 246 642 248 644
rect 251 642 253 644
rect 256 642 258 644
rect 261 642 263 644
rect 266 642 268 644
rect 271 642 273 644
rect 276 642 278 644
rect 281 642 283 644
rect 286 642 288 644
rect 291 642 293 644
rect 296 642 298 644
rect 301 642 303 644
rect 306 642 308 644
rect 311 642 313 644
rect 316 642 318 644
rect 325 643 327 645
rect 333 642 335 644
rect 338 642 340 644
rect 2 638 4 640
rect 7 638 9 640
rect 20 637 22 639
rect 25 637 27 639
rect 33 638 35 640
rect 42 637 44 639
rect 47 637 49 639
rect 52 637 54 639
rect 57 637 59 639
rect 62 637 64 639
rect 67 637 69 639
rect 72 637 74 639
rect 77 637 79 639
rect 82 637 84 639
rect 87 637 89 639
rect 92 637 94 639
rect 97 637 99 639
rect 102 637 104 639
rect 107 637 109 639
rect 112 637 114 639
rect 117 637 119 639
rect 122 637 124 639
rect 127 637 129 639
rect 132 637 134 639
rect 137 637 139 639
rect 142 637 144 639
rect 147 637 149 639
rect 152 637 154 639
rect 157 637 159 639
rect 162 637 164 639
rect 169 638 171 640
rect 177 637 179 639
rect 182 637 184 639
rect 189 638 191 640
rect 196 637 198 639
rect 201 637 203 639
rect 206 637 208 639
rect 211 637 213 639
rect 216 637 218 639
rect 221 637 223 639
rect 226 637 228 639
rect 231 637 233 639
rect 236 637 238 639
rect 241 637 243 639
rect 246 637 248 639
rect 251 637 253 639
rect 256 637 258 639
rect 261 637 263 639
rect 266 637 268 639
rect 271 637 273 639
rect 276 637 278 639
rect 281 637 283 639
rect 286 637 288 639
rect 291 637 293 639
rect 296 637 298 639
rect 301 637 303 639
rect 306 637 308 639
rect 311 637 313 639
rect 316 637 318 639
rect 325 638 327 640
rect 333 637 335 639
rect 338 637 340 639
rect 351 638 353 640
rect 356 638 358 640
rect 20 632 22 634
rect 25 632 27 634
rect 33 633 35 635
rect 169 633 171 635
rect 177 632 179 634
rect 182 632 184 634
rect 189 633 191 635
rect 325 633 327 635
rect 333 632 335 634
rect 338 632 340 634
rect 2 630 4 632
rect 7 630 9 632
rect 351 630 353 632
rect 356 630 358 632
rect 33 628 35 630
rect 41 627 43 629
rect 51 627 53 629
rect 61 627 63 629
rect 71 627 73 629
rect 81 627 83 629
rect 91 627 93 629
rect 101 627 103 629
rect 111 627 113 629
rect 150 627 152 629
rect 160 627 162 629
rect 169 628 171 630
rect 189 628 191 630
rect 198 627 200 629
rect 208 627 210 629
rect 247 627 249 629
rect 257 627 259 629
rect 267 627 269 629
rect 277 627 279 629
rect 287 627 289 629
rect 297 627 299 629
rect 307 627 309 629
rect 317 627 319 629
rect 325 628 327 630
rect 2 622 4 624
rect 7 622 9 624
rect 33 623 35 625
rect 41 622 43 624
rect 51 622 53 624
rect 61 622 63 624
rect 71 622 73 624
rect 81 622 83 624
rect 91 622 93 624
rect 101 622 103 624
rect 111 622 113 624
rect 150 622 152 624
rect 160 622 162 624
rect 169 623 171 625
rect 189 623 191 625
rect 198 622 200 624
rect 208 622 210 624
rect 247 622 249 624
rect 257 622 259 624
rect 267 622 269 624
rect 277 622 279 624
rect 287 622 289 624
rect 297 622 299 624
rect 307 622 309 624
rect 317 622 319 624
rect 325 623 327 625
rect 351 622 353 624
rect 356 622 358 624
rect 33 618 35 620
rect 41 617 43 619
rect 51 617 53 619
rect 61 617 63 619
rect 71 617 73 619
rect 81 617 83 619
rect 91 617 93 619
rect 101 617 103 619
rect 111 617 113 619
rect 150 617 152 619
rect 160 617 162 619
rect 169 618 171 620
rect 189 618 191 620
rect 198 617 200 619
rect 208 617 210 619
rect 247 617 249 619
rect 257 617 259 619
rect 267 617 269 619
rect 277 617 279 619
rect 287 617 289 619
rect 297 617 299 619
rect 307 617 309 619
rect 317 617 319 619
rect 325 618 327 620
rect 2 614 4 616
rect 7 614 9 616
rect 20 612 22 614
rect 25 612 27 614
rect 33 613 35 615
rect 169 613 171 615
rect 177 612 179 614
rect 182 612 184 614
rect 189 613 191 615
rect 325 613 327 615
rect 351 614 353 616
rect 356 614 358 616
rect 333 612 335 614
rect 338 612 340 614
rect 2 606 4 608
rect 7 606 9 608
rect 20 607 22 609
rect 25 607 27 609
rect 33 608 35 610
rect 42 607 44 609
rect 47 607 49 609
rect 52 607 54 609
rect 57 607 59 609
rect 62 607 64 609
rect 67 607 69 609
rect 72 607 74 609
rect 77 607 79 609
rect 82 607 84 609
rect 87 607 89 609
rect 92 607 94 609
rect 97 607 99 609
rect 102 607 104 609
rect 107 607 109 609
rect 112 607 114 609
rect 117 607 119 609
rect 122 607 124 609
rect 127 607 129 609
rect 132 607 134 609
rect 137 607 139 609
rect 142 607 144 609
rect 147 607 149 609
rect 152 607 154 609
rect 157 607 159 609
rect 162 607 164 609
rect 169 608 171 610
rect 177 607 179 609
rect 182 607 184 609
rect 189 608 191 610
rect 196 607 198 609
rect 201 607 203 609
rect 206 607 208 609
rect 211 607 213 609
rect 216 607 218 609
rect 221 607 223 609
rect 226 607 228 609
rect 231 607 233 609
rect 236 607 238 609
rect 241 607 243 609
rect 246 607 248 609
rect 251 607 253 609
rect 256 607 258 609
rect 261 607 263 609
rect 266 607 268 609
rect 271 607 273 609
rect 276 607 278 609
rect 281 607 283 609
rect 286 607 288 609
rect 291 607 293 609
rect 296 607 298 609
rect 301 607 303 609
rect 306 607 308 609
rect 311 607 313 609
rect 316 607 318 609
rect 325 608 327 610
rect 333 607 335 609
rect 338 607 340 609
rect 351 606 353 608
rect 356 606 358 608
rect 20 602 22 604
rect 25 602 27 604
rect 33 603 35 605
rect 42 602 44 604
rect 47 602 49 604
rect 52 602 54 604
rect 57 602 59 604
rect 62 602 64 604
rect 67 602 69 604
rect 72 602 74 604
rect 77 602 79 604
rect 82 602 84 604
rect 87 602 89 604
rect 92 602 94 604
rect 97 602 99 604
rect 102 602 104 604
rect 107 602 109 604
rect 112 602 114 604
rect 117 602 119 604
rect 122 602 124 604
rect 127 602 129 604
rect 132 602 134 604
rect 137 602 139 604
rect 142 602 144 604
rect 147 602 149 604
rect 152 602 154 604
rect 157 602 159 604
rect 162 602 164 604
rect 169 603 171 605
rect 177 602 179 604
rect 182 602 184 604
rect 189 603 191 605
rect 196 602 198 604
rect 201 602 203 604
rect 206 602 208 604
rect 211 602 213 604
rect 216 602 218 604
rect 221 602 223 604
rect 226 602 228 604
rect 231 602 233 604
rect 236 602 238 604
rect 241 602 243 604
rect 246 602 248 604
rect 251 602 253 604
rect 256 602 258 604
rect 261 602 263 604
rect 266 602 268 604
rect 271 602 273 604
rect 276 602 278 604
rect 281 602 283 604
rect 286 602 288 604
rect 291 602 293 604
rect 296 602 298 604
rect 301 602 303 604
rect 306 602 308 604
rect 311 602 313 604
rect 316 602 318 604
rect 325 603 327 605
rect 333 602 335 604
rect 338 602 340 604
rect 2 598 4 600
rect 7 598 9 600
rect 20 597 22 599
rect 25 597 27 599
rect 33 598 35 600
rect 42 597 44 599
rect 47 597 49 599
rect 52 597 54 599
rect 57 597 59 599
rect 62 597 64 599
rect 67 597 69 599
rect 72 597 74 599
rect 77 597 79 599
rect 82 597 84 599
rect 87 597 89 599
rect 92 597 94 599
rect 97 597 99 599
rect 102 597 104 599
rect 107 597 109 599
rect 112 597 114 599
rect 117 597 119 599
rect 122 597 124 599
rect 127 597 129 599
rect 132 597 134 599
rect 137 597 139 599
rect 142 597 144 599
rect 147 597 149 599
rect 152 597 154 599
rect 157 597 159 599
rect 162 597 164 599
rect 169 598 171 600
rect 177 597 179 599
rect 182 597 184 599
rect 189 598 191 600
rect 196 597 198 599
rect 201 597 203 599
rect 206 597 208 599
rect 211 597 213 599
rect 216 597 218 599
rect 221 597 223 599
rect 226 597 228 599
rect 231 597 233 599
rect 236 597 238 599
rect 241 597 243 599
rect 246 597 248 599
rect 251 597 253 599
rect 256 597 258 599
rect 261 597 263 599
rect 266 597 268 599
rect 271 597 273 599
rect 276 597 278 599
rect 281 597 283 599
rect 286 597 288 599
rect 291 597 293 599
rect 296 597 298 599
rect 301 597 303 599
rect 306 597 308 599
rect 311 597 313 599
rect 316 597 318 599
rect 325 598 327 600
rect 333 597 335 599
rect 338 597 340 599
rect 351 598 353 600
rect 356 598 358 600
rect 20 592 22 594
rect 25 592 27 594
rect 33 593 35 595
rect 42 592 44 594
rect 47 592 49 594
rect 52 592 54 594
rect 57 592 59 594
rect 62 592 64 594
rect 67 592 69 594
rect 72 592 74 594
rect 77 592 79 594
rect 82 592 84 594
rect 87 592 89 594
rect 92 592 94 594
rect 97 592 99 594
rect 102 592 104 594
rect 107 592 109 594
rect 112 592 114 594
rect 117 592 119 594
rect 122 592 124 594
rect 127 592 129 594
rect 132 592 134 594
rect 137 592 139 594
rect 142 592 144 594
rect 147 592 149 594
rect 152 592 154 594
rect 157 592 159 594
rect 162 592 164 594
rect 169 593 171 595
rect 177 592 179 594
rect 182 592 184 594
rect 189 593 191 595
rect 196 592 198 594
rect 201 592 203 594
rect 206 592 208 594
rect 211 592 213 594
rect 216 592 218 594
rect 221 592 223 594
rect 226 592 228 594
rect 231 592 233 594
rect 236 592 238 594
rect 241 592 243 594
rect 246 592 248 594
rect 251 592 253 594
rect 256 592 258 594
rect 261 592 263 594
rect 266 592 268 594
rect 271 592 273 594
rect 276 592 278 594
rect 281 592 283 594
rect 286 592 288 594
rect 291 592 293 594
rect 296 592 298 594
rect 301 592 303 594
rect 306 592 308 594
rect 311 592 313 594
rect 316 592 318 594
rect 325 593 327 595
rect 333 592 335 594
rect 338 592 340 594
rect 2 590 4 592
rect 7 590 9 592
rect 351 590 353 592
rect 356 590 358 592
rect 20 587 22 589
rect 25 587 27 589
rect 33 588 35 590
rect 42 587 44 589
rect 47 587 49 589
rect 52 587 54 589
rect 57 587 59 589
rect 62 587 64 589
rect 67 587 69 589
rect 72 587 74 589
rect 77 587 79 589
rect 82 587 84 589
rect 87 587 89 589
rect 92 587 94 589
rect 97 587 99 589
rect 102 587 104 589
rect 107 587 109 589
rect 112 587 114 589
rect 117 587 119 589
rect 122 587 124 589
rect 127 587 129 589
rect 132 587 134 589
rect 137 587 139 589
rect 142 587 144 589
rect 147 587 149 589
rect 152 587 154 589
rect 157 587 159 589
rect 162 587 164 589
rect 169 588 171 590
rect 177 587 179 589
rect 182 587 184 589
rect 189 588 191 590
rect 196 587 198 589
rect 201 587 203 589
rect 206 587 208 589
rect 211 587 213 589
rect 216 587 218 589
rect 221 587 223 589
rect 226 587 228 589
rect 231 587 233 589
rect 236 587 238 589
rect 241 587 243 589
rect 246 587 248 589
rect 251 587 253 589
rect 256 587 258 589
rect 261 587 263 589
rect 266 587 268 589
rect 271 587 273 589
rect 276 587 278 589
rect 281 587 283 589
rect 286 587 288 589
rect 291 587 293 589
rect 296 587 298 589
rect 301 587 303 589
rect 306 587 308 589
rect 311 587 313 589
rect 316 587 318 589
rect 325 588 327 590
rect 333 587 335 589
rect 338 587 340 589
rect 2 582 4 584
rect 7 582 9 584
rect 20 582 22 584
rect 25 582 27 584
rect 33 583 35 585
rect 42 582 44 584
rect 47 582 49 584
rect 52 582 54 584
rect 57 582 59 584
rect 62 582 64 584
rect 67 582 69 584
rect 72 582 74 584
rect 77 582 79 584
rect 82 582 84 584
rect 87 582 89 584
rect 92 582 94 584
rect 97 582 99 584
rect 102 582 104 584
rect 107 582 109 584
rect 112 582 114 584
rect 117 582 119 584
rect 122 582 124 584
rect 127 582 129 584
rect 132 582 134 584
rect 137 582 139 584
rect 142 582 144 584
rect 147 582 149 584
rect 152 582 154 584
rect 157 582 159 584
rect 162 582 164 584
rect 169 583 171 585
rect 177 582 179 584
rect 182 582 184 584
rect 189 583 191 585
rect 196 582 198 584
rect 201 582 203 584
rect 206 582 208 584
rect 211 582 213 584
rect 216 582 218 584
rect 221 582 223 584
rect 226 582 228 584
rect 231 582 233 584
rect 236 582 238 584
rect 241 582 243 584
rect 246 582 248 584
rect 251 582 253 584
rect 256 582 258 584
rect 261 582 263 584
rect 266 582 268 584
rect 271 582 273 584
rect 276 582 278 584
rect 281 582 283 584
rect 286 582 288 584
rect 291 582 293 584
rect 296 582 298 584
rect 301 582 303 584
rect 306 582 308 584
rect 311 582 313 584
rect 316 582 318 584
rect 325 583 327 585
rect 333 582 335 584
rect 338 582 340 584
rect 351 582 353 584
rect 356 582 358 584
rect 20 577 22 579
rect 25 577 27 579
rect 33 578 35 580
rect 42 577 44 579
rect 47 577 49 579
rect 52 577 54 579
rect 57 577 59 579
rect 62 577 64 579
rect 67 577 69 579
rect 72 577 74 579
rect 77 577 79 579
rect 82 577 84 579
rect 87 577 89 579
rect 92 577 94 579
rect 97 577 99 579
rect 102 577 104 579
rect 107 577 109 579
rect 112 577 114 579
rect 117 577 119 579
rect 122 577 124 579
rect 127 577 129 579
rect 132 577 134 579
rect 137 577 139 579
rect 142 577 144 579
rect 147 577 149 579
rect 152 577 154 579
rect 157 577 159 579
rect 162 577 164 579
rect 169 578 171 580
rect 177 577 179 579
rect 182 577 184 579
rect 189 578 191 580
rect 196 577 198 579
rect 201 577 203 579
rect 206 577 208 579
rect 211 577 213 579
rect 216 577 218 579
rect 221 577 223 579
rect 226 577 228 579
rect 231 577 233 579
rect 236 577 238 579
rect 241 577 243 579
rect 246 577 248 579
rect 251 577 253 579
rect 256 577 258 579
rect 261 577 263 579
rect 266 577 268 579
rect 271 577 273 579
rect 276 577 278 579
rect 281 577 283 579
rect 286 577 288 579
rect 291 577 293 579
rect 296 577 298 579
rect 301 577 303 579
rect 306 577 308 579
rect 311 577 313 579
rect 316 577 318 579
rect 325 578 327 580
rect 333 577 335 579
rect 338 577 340 579
rect 2 574 4 576
rect 7 574 9 576
rect 20 572 22 574
rect 25 572 27 574
rect 33 573 35 575
rect 42 572 44 574
rect 47 572 49 574
rect 52 572 54 574
rect 57 572 59 574
rect 62 572 64 574
rect 67 572 69 574
rect 72 572 74 574
rect 77 572 79 574
rect 82 572 84 574
rect 87 572 89 574
rect 92 572 94 574
rect 97 572 99 574
rect 102 572 104 574
rect 107 572 109 574
rect 112 572 114 574
rect 117 572 119 574
rect 122 572 124 574
rect 127 572 129 574
rect 132 572 134 574
rect 137 572 139 574
rect 142 572 144 574
rect 147 572 149 574
rect 152 572 154 574
rect 157 572 159 574
rect 162 572 164 574
rect 169 573 171 575
rect 177 572 179 574
rect 182 572 184 574
rect 189 573 191 575
rect 196 572 198 574
rect 201 572 203 574
rect 206 572 208 574
rect 211 572 213 574
rect 216 572 218 574
rect 221 572 223 574
rect 226 572 228 574
rect 231 572 233 574
rect 236 572 238 574
rect 241 572 243 574
rect 246 572 248 574
rect 251 572 253 574
rect 256 572 258 574
rect 261 572 263 574
rect 266 572 268 574
rect 271 572 273 574
rect 276 572 278 574
rect 281 572 283 574
rect 286 572 288 574
rect 291 572 293 574
rect 296 572 298 574
rect 301 572 303 574
rect 306 572 308 574
rect 311 572 313 574
rect 316 572 318 574
rect 325 573 327 575
rect 351 574 353 576
rect 356 574 358 576
rect 333 572 335 574
rect 338 572 340 574
rect 2 566 4 568
rect 7 566 9 568
rect 20 567 22 569
rect 25 567 27 569
rect 33 568 35 570
rect 169 568 171 570
rect 177 567 179 569
rect 182 567 184 569
rect 189 568 191 570
rect 325 568 327 570
rect 333 567 335 569
rect 338 567 340 569
rect 351 566 353 568
rect 356 566 358 568
rect 41 562 43 564
rect 51 562 53 564
rect 61 562 63 564
rect 71 562 73 564
rect 81 562 83 564
rect 91 562 93 564
rect 101 562 103 564
rect 111 562 113 564
rect 150 562 152 564
rect 160 562 162 564
rect 198 562 200 564
rect 208 562 210 564
rect 247 562 249 564
rect 257 562 259 564
rect 267 562 269 564
rect 277 562 279 564
rect 287 562 289 564
rect 297 562 299 564
rect 307 562 309 564
rect 317 562 319 564
rect 2 558 4 560
rect 7 558 9 560
rect 41 557 43 559
rect 51 557 53 559
rect 61 557 63 559
rect 71 557 73 559
rect 81 557 83 559
rect 91 557 93 559
rect 101 557 103 559
rect 111 557 113 559
rect 150 557 152 559
rect 160 557 162 559
rect 198 557 200 559
rect 208 557 210 559
rect 247 557 249 559
rect 257 557 259 559
rect 267 557 269 559
rect 277 557 279 559
rect 287 557 289 559
rect 297 557 299 559
rect 307 557 309 559
rect 317 557 319 559
rect 351 558 353 560
rect 356 558 358 560
rect 41 552 43 554
rect 51 552 53 554
rect 61 552 63 554
rect 71 552 73 554
rect 81 552 83 554
rect 91 552 93 554
rect 101 552 103 554
rect 111 552 113 554
rect 150 552 152 554
rect 160 552 162 554
rect 198 552 200 554
rect 208 552 210 554
rect 247 552 249 554
rect 257 552 259 554
rect 267 552 269 554
rect 277 552 279 554
rect 287 552 289 554
rect 297 552 299 554
rect 307 552 309 554
rect 317 552 319 554
rect 2 550 4 552
rect 7 550 9 552
rect 351 550 353 552
rect 356 550 358 552
rect 2 542 4 544
rect 7 542 9 544
rect 351 542 353 544
rect 356 542 358 544
rect 9 534 11 536
rect 17 534 19 536
rect 25 534 27 536
rect 41 534 43 536
rect 49 534 51 536
rect 57 534 59 536
rect 65 534 67 536
rect 73 534 75 536
rect 81 534 83 536
rect 89 534 91 536
rect 97 534 99 536
rect 105 534 107 536
rect 113 534 115 536
rect 150 534 152 536
rect 158 534 160 536
rect 181 534 183 536
rect 198 534 200 536
rect 206 534 208 536
rect 245 534 247 536
rect 253 534 255 536
rect 261 534 263 536
rect 269 534 271 536
rect 277 534 279 536
rect 285 534 287 536
rect 293 534 295 536
rect 301 534 303 536
rect 309 534 311 536
rect 317 534 319 536
rect 333 534 335 536
rect 341 534 343 536
rect 349 534 351 536
rect 9 529 11 531
rect 17 529 19 531
rect 25 529 27 531
rect 41 529 43 531
rect 49 529 51 531
rect 57 529 59 531
rect 65 529 67 531
rect 73 529 75 531
rect 81 529 83 531
rect 89 529 91 531
rect 97 529 99 531
rect 105 529 107 531
rect 113 529 115 531
rect 150 529 152 531
rect 158 529 160 531
rect 181 529 183 531
rect 198 529 200 531
rect 206 529 208 531
rect 245 529 247 531
rect 253 529 255 531
rect 261 529 263 531
rect 269 529 271 531
rect 277 529 279 531
rect 285 529 287 531
rect 293 529 295 531
rect 301 529 303 531
rect 309 529 311 531
rect 317 529 319 531
rect 333 529 335 531
rect 341 529 343 531
rect 349 529 351 531
rect 9 517 11 519
rect 17 517 19 519
rect 25 517 27 519
rect 41 517 43 519
rect 49 517 51 519
rect 57 517 59 519
rect 65 517 67 519
rect 73 517 75 519
rect 81 517 83 519
rect 89 517 91 519
rect 97 517 99 519
rect 105 517 107 519
rect 113 517 115 519
rect 150 517 152 519
rect 158 517 160 519
rect 181 517 183 519
rect 198 517 200 519
rect 206 517 208 519
rect 245 517 247 519
rect 253 517 255 519
rect 261 517 263 519
rect 269 517 271 519
rect 277 517 279 519
rect 285 517 287 519
rect 293 517 295 519
rect 301 517 303 519
rect 309 517 311 519
rect 317 517 319 519
rect 333 517 335 519
rect 341 517 343 519
rect 349 517 351 519
rect 9 512 11 514
rect 17 512 19 514
rect 25 512 27 514
rect 41 512 43 514
rect 49 512 51 514
rect 57 512 59 514
rect 65 512 67 514
rect 73 512 75 514
rect 81 512 83 514
rect 89 512 91 514
rect 97 512 99 514
rect 105 512 107 514
rect 113 512 115 514
rect 150 512 152 514
rect 158 512 160 514
rect 181 512 183 514
rect 198 512 200 514
rect 206 512 208 514
rect 245 512 247 514
rect 253 512 255 514
rect 261 512 263 514
rect 269 512 271 514
rect 277 512 279 514
rect 285 512 287 514
rect 293 512 295 514
rect 301 512 303 514
rect 309 512 311 514
rect 317 512 319 514
rect 333 512 335 514
rect 341 512 343 514
rect 349 512 351 514
rect 9 489 11 491
rect 17 489 19 491
rect 25 489 27 491
rect 33 489 35 491
rect 41 489 43 491
rect 49 489 51 491
rect 57 489 59 491
rect 65 489 67 491
rect 73 489 75 491
rect 81 489 83 491
rect 89 489 91 491
rect 97 489 99 491
rect 105 489 107 491
rect 113 489 115 491
rect 150 489 152 491
rect 158 489 160 491
rect 181 489 183 491
rect 198 489 200 491
rect 206 489 208 491
rect 245 489 247 491
rect 253 489 255 491
rect 261 489 263 491
rect 269 489 271 491
rect 277 489 279 491
rect 285 489 287 491
rect 293 489 295 491
rect 301 489 303 491
rect 309 489 311 491
rect 317 489 319 491
rect 325 489 327 491
rect 333 489 335 491
rect 341 489 343 491
rect 349 489 351 491
rect 9 484 11 486
rect 17 484 19 486
rect 25 484 27 486
rect 33 484 35 486
rect 41 484 43 486
rect 49 484 51 486
rect 57 484 59 486
rect 65 484 67 486
rect 73 484 75 486
rect 81 484 83 486
rect 89 484 91 486
rect 97 484 99 486
rect 105 484 107 486
rect 113 484 115 486
rect 150 484 152 486
rect 158 484 160 486
rect 181 484 183 486
rect 198 484 200 486
rect 206 484 208 486
rect 245 484 247 486
rect 253 484 255 486
rect 261 484 263 486
rect 269 484 271 486
rect 277 484 279 486
rect 285 484 287 486
rect 293 484 295 486
rect 301 484 303 486
rect 309 484 311 486
rect 317 484 319 486
rect 325 484 327 486
rect 333 484 335 486
rect 341 484 343 486
rect 349 484 351 486
rect 9 472 11 474
rect 17 472 19 474
rect 25 472 27 474
rect 33 472 35 474
rect 41 472 43 474
rect 49 472 51 474
rect 57 472 59 474
rect 65 472 67 474
rect 73 472 75 474
rect 81 472 83 474
rect 89 472 91 474
rect 97 472 99 474
rect 105 472 107 474
rect 113 472 115 474
rect 150 472 152 474
rect 158 472 160 474
rect 181 472 183 474
rect 198 472 200 474
rect 206 472 208 474
rect 245 472 247 474
rect 253 472 255 474
rect 261 472 263 474
rect 269 472 271 474
rect 277 472 279 474
rect 285 472 287 474
rect 293 472 295 474
rect 301 472 303 474
rect 309 472 311 474
rect 317 472 319 474
rect 325 472 327 474
rect 333 472 335 474
rect 341 472 343 474
rect 349 472 351 474
rect 357 472 359 474
rect 9 467 11 469
rect 17 467 19 469
rect 25 467 27 469
rect 33 467 35 469
rect 41 467 43 469
rect 49 467 51 469
rect 57 467 59 469
rect 65 467 67 469
rect 73 467 75 469
rect 81 467 83 469
rect 89 467 91 469
rect 97 467 99 469
rect 105 467 107 469
rect 113 467 115 469
rect 150 467 152 469
rect 158 467 160 469
rect 181 467 183 469
rect 198 467 200 469
rect 206 467 208 469
rect 245 467 247 469
rect 253 467 255 469
rect 261 467 263 469
rect 269 467 271 469
rect 277 467 279 469
rect 285 467 287 469
rect 293 467 295 469
rect 301 467 303 469
rect 309 467 311 469
rect 317 467 319 469
rect 325 467 327 469
rect 333 467 335 469
rect 341 467 343 469
rect 349 467 351 469
rect 357 467 359 469
rect 2 459 4 461
rect 7 459 9 461
rect 351 459 353 461
rect 356 459 358 461
rect 2 451 4 453
rect 7 451 9 453
rect 351 451 353 453
rect 356 451 358 453
rect 41 449 43 451
rect 51 449 53 451
rect 61 449 63 451
rect 71 449 73 451
rect 81 449 83 451
rect 91 449 93 451
rect 101 449 103 451
rect 111 449 113 451
rect 154 449 156 451
rect 204 449 206 451
rect 247 449 249 451
rect 257 449 259 451
rect 267 449 269 451
rect 277 449 279 451
rect 287 449 289 451
rect 297 449 299 451
rect 307 449 309 451
rect 317 449 319 451
rect 2 443 4 445
rect 7 443 9 445
rect 41 444 43 446
rect 51 444 53 446
rect 61 444 63 446
rect 71 444 73 446
rect 81 444 83 446
rect 91 444 93 446
rect 101 444 103 446
rect 111 444 113 446
rect 154 444 156 446
rect 204 444 206 446
rect 247 444 249 446
rect 257 444 259 446
rect 267 444 269 446
rect 277 444 279 446
rect 287 444 289 446
rect 297 444 299 446
rect 307 444 309 446
rect 317 444 319 446
rect 351 443 353 445
rect 356 443 358 445
rect 41 439 43 441
rect 51 439 53 441
rect 61 439 63 441
rect 71 439 73 441
rect 81 439 83 441
rect 91 439 93 441
rect 101 439 103 441
rect 111 439 113 441
rect 154 439 156 441
rect 204 439 206 441
rect 247 439 249 441
rect 257 439 259 441
rect 267 439 269 441
rect 277 439 279 441
rect 287 439 289 441
rect 297 439 299 441
rect 307 439 309 441
rect 317 439 319 441
rect 2 435 4 437
rect 7 435 9 437
rect 20 434 22 436
rect 25 434 27 436
rect 177 434 179 436
rect 182 434 184 436
rect 333 434 335 436
rect 338 434 340 436
rect 351 435 353 437
rect 356 435 358 437
rect 33 431 35 433
rect 162 431 164 433
rect 196 431 198 433
rect 325 431 327 433
rect 20 429 22 431
rect 25 429 27 431
rect 42 429 44 431
rect 47 429 49 431
rect 52 429 54 431
rect 57 429 59 431
rect 62 429 64 431
rect 67 429 69 431
rect 72 429 74 431
rect 77 429 79 431
rect 82 429 84 431
rect 87 429 89 431
rect 92 429 94 431
rect 97 429 99 431
rect 102 429 104 431
rect 107 429 109 431
rect 112 429 114 431
rect 117 429 119 431
rect 122 429 124 431
rect 127 429 129 431
rect 132 429 134 431
rect 137 429 139 431
rect 142 429 144 431
rect 147 429 149 431
rect 152 429 154 431
rect 177 429 179 431
rect 182 429 184 431
rect 206 429 208 431
rect 211 429 213 431
rect 216 429 218 431
rect 221 429 223 431
rect 226 429 228 431
rect 231 429 233 431
rect 236 429 238 431
rect 241 429 243 431
rect 246 429 248 431
rect 251 429 253 431
rect 256 429 258 431
rect 261 429 263 431
rect 266 429 268 431
rect 271 429 273 431
rect 276 429 278 431
rect 281 429 283 431
rect 286 429 288 431
rect 291 429 293 431
rect 296 429 298 431
rect 301 429 303 431
rect 306 429 308 431
rect 311 429 313 431
rect 316 429 318 431
rect 333 429 335 431
rect 338 429 340 431
rect 2 427 4 429
rect 7 427 9 429
rect 33 426 35 428
rect 162 426 164 428
rect 196 426 198 428
rect 325 426 327 428
rect 351 427 353 429
rect 356 427 358 429
rect 20 424 22 426
rect 25 424 27 426
rect 42 424 44 426
rect 47 424 49 426
rect 52 424 54 426
rect 57 424 59 426
rect 62 424 64 426
rect 67 424 69 426
rect 72 424 74 426
rect 77 424 79 426
rect 82 424 84 426
rect 87 424 89 426
rect 92 424 94 426
rect 97 424 99 426
rect 102 424 104 426
rect 107 424 109 426
rect 112 424 114 426
rect 117 424 119 426
rect 122 424 124 426
rect 127 424 129 426
rect 132 424 134 426
rect 137 424 139 426
rect 142 424 144 426
rect 147 424 149 426
rect 152 424 154 426
rect 177 424 179 426
rect 182 424 184 426
rect 206 424 208 426
rect 211 424 213 426
rect 216 424 218 426
rect 221 424 223 426
rect 226 424 228 426
rect 231 424 233 426
rect 236 424 238 426
rect 241 424 243 426
rect 246 424 248 426
rect 251 424 253 426
rect 256 424 258 426
rect 261 424 263 426
rect 266 424 268 426
rect 271 424 273 426
rect 276 424 278 426
rect 281 424 283 426
rect 286 424 288 426
rect 291 424 293 426
rect 296 424 298 426
rect 301 424 303 426
rect 306 424 308 426
rect 311 424 313 426
rect 316 424 318 426
rect 333 424 335 426
rect 338 424 340 426
rect 33 421 35 423
rect 162 421 164 423
rect 196 421 198 423
rect 325 421 327 423
rect 2 419 4 421
rect 7 419 9 421
rect 20 419 22 421
rect 25 419 27 421
rect 42 419 44 421
rect 47 419 49 421
rect 52 419 54 421
rect 57 419 59 421
rect 62 419 64 421
rect 67 419 69 421
rect 72 419 74 421
rect 77 419 79 421
rect 82 419 84 421
rect 87 419 89 421
rect 92 419 94 421
rect 97 419 99 421
rect 102 419 104 421
rect 107 419 109 421
rect 112 419 114 421
rect 117 419 119 421
rect 122 419 124 421
rect 127 419 129 421
rect 132 419 134 421
rect 137 419 139 421
rect 142 419 144 421
rect 147 419 149 421
rect 152 419 154 421
rect 177 419 179 421
rect 182 419 184 421
rect 206 419 208 421
rect 211 419 213 421
rect 216 419 218 421
rect 221 419 223 421
rect 226 419 228 421
rect 231 419 233 421
rect 236 419 238 421
rect 241 419 243 421
rect 246 419 248 421
rect 251 419 253 421
rect 256 419 258 421
rect 261 419 263 421
rect 266 419 268 421
rect 271 419 273 421
rect 276 419 278 421
rect 281 419 283 421
rect 286 419 288 421
rect 291 419 293 421
rect 296 419 298 421
rect 301 419 303 421
rect 306 419 308 421
rect 311 419 313 421
rect 316 419 318 421
rect 333 419 335 421
rect 338 419 340 421
rect 351 419 353 421
rect 356 419 358 421
rect 33 416 35 418
rect 162 416 164 418
rect 196 416 198 418
rect 325 416 327 418
rect 20 414 22 416
rect 25 414 27 416
rect 42 414 44 416
rect 47 414 49 416
rect 52 414 54 416
rect 57 414 59 416
rect 62 414 64 416
rect 67 414 69 416
rect 72 414 74 416
rect 77 414 79 416
rect 82 414 84 416
rect 87 414 89 416
rect 92 414 94 416
rect 97 414 99 416
rect 102 414 104 416
rect 107 414 109 416
rect 112 414 114 416
rect 117 414 119 416
rect 122 414 124 416
rect 127 414 129 416
rect 132 414 134 416
rect 137 414 139 416
rect 142 414 144 416
rect 147 414 149 416
rect 152 414 154 416
rect 177 414 179 416
rect 182 414 184 416
rect 206 414 208 416
rect 211 414 213 416
rect 216 414 218 416
rect 221 414 223 416
rect 226 414 228 416
rect 231 414 233 416
rect 236 414 238 416
rect 241 414 243 416
rect 246 414 248 416
rect 251 414 253 416
rect 256 414 258 416
rect 261 414 263 416
rect 266 414 268 416
rect 271 414 273 416
rect 276 414 278 416
rect 281 414 283 416
rect 286 414 288 416
rect 291 414 293 416
rect 296 414 298 416
rect 301 414 303 416
rect 306 414 308 416
rect 311 414 313 416
rect 316 414 318 416
rect 333 414 335 416
rect 338 414 340 416
rect 2 411 4 413
rect 7 411 9 413
rect 33 411 35 413
rect 162 411 164 413
rect 196 411 198 413
rect 325 411 327 413
rect 351 411 353 413
rect 356 411 358 413
rect 20 409 22 411
rect 25 409 27 411
rect 42 409 44 411
rect 47 409 49 411
rect 52 409 54 411
rect 57 409 59 411
rect 62 409 64 411
rect 67 409 69 411
rect 72 409 74 411
rect 77 409 79 411
rect 82 409 84 411
rect 87 409 89 411
rect 92 409 94 411
rect 97 409 99 411
rect 102 409 104 411
rect 107 409 109 411
rect 112 409 114 411
rect 117 409 119 411
rect 122 409 124 411
rect 127 409 129 411
rect 132 409 134 411
rect 137 409 139 411
rect 142 409 144 411
rect 147 409 149 411
rect 152 409 154 411
rect 177 409 179 411
rect 182 409 184 411
rect 206 409 208 411
rect 211 409 213 411
rect 216 409 218 411
rect 221 409 223 411
rect 226 409 228 411
rect 231 409 233 411
rect 236 409 238 411
rect 241 409 243 411
rect 246 409 248 411
rect 251 409 253 411
rect 256 409 258 411
rect 261 409 263 411
rect 266 409 268 411
rect 271 409 273 411
rect 276 409 278 411
rect 281 409 283 411
rect 286 409 288 411
rect 291 409 293 411
rect 296 409 298 411
rect 301 409 303 411
rect 306 409 308 411
rect 311 409 313 411
rect 316 409 318 411
rect 333 409 335 411
rect 338 409 340 411
rect 33 406 35 408
rect 162 406 164 408
rect 196 406 198 408
rect 325 406 327 408
rect 2 403 4 405
rect 7 403 9 405
rect 20 404 22 406
rect 25 404 27 406
rect 42 404 44 406
rect 47 404 49 406
rect 52 404 54 406
rect 57 404 59 406
rect 62 404 64 406
rect 67 404 69 406
rect 72 404 74 406
rect 77 404 79 406
rect 82 404 84 406
rect 87 404 89 406
rect 92 404 94 406
rect 97 404 99 406
rect 102 404 104 406
rect 107 404 109 406
rect 112 404 114 406
rect 117 404 119 406
rect 122 404 124 406
rect 127 404 129 406
rect 132 404 134 406
rect 137 404 139 406
rect 142 404 144 406
rect 147 404 149 406
rect 152 404 154 406
rect 177 404 179 406
rect 182 404 184 406
rect 206 404 208 406
rect 211 404 213 406
rect 216 404 218 406
rect 221 404 223 406
rect 226 404 228 406
rect 231 404 233 406
rect 236 404 238 406
rect 241 404 243 406
rect 246 404 248 406
rect 251 404 253 406
rect 256 404 258 406
rect 261 404 263 406
rect 266 404 268 406
rect 271 404 273 406
rect 276 404 278 406
rect 281 404 283 406
rect 286 404 288 406
rect 291 404 293 406
rect 296 404 298 406
rect 301 404 303 406
rect 306 404 308 406
rect 311 404 313 406
rect 316 404 318 406
rect 333 404 335 406
rect 338 404 340 406
rect 351 403 353 405
rect 356 403 358 405
rect 33 401 35 403
rect 162 401 164 403
rect 196 401 198 403
rect 325 401 327 403
rect 20 399 22 401
rect 25 399 27 401
rect 42 399 44 401
rect 47 399 49 401
rect 52 399 54 401
rect 57 399 59 401
rect 62 399 64 401
rect 67 399 69 401
rect 72 399 74 401
rect 77 399 79 401
rect 82 399 84 401
rect 87 399 89 401
rect 92 399 94 401
rect 97 399 99 401
rect 102 399 104 401
rect 107 399 109 401
rect 112 399 114 401
rect 117 399 119 401
rect 122 399 124 401
rect 127 399 129 401
rect 132 399 134 401
rect 137 399 139 401
rect 142 399 144 401
rect 147 399 149 401
rect 152 399 154 401
rect 177 399 179 401
rect 182 399 184 401
rect 206 399 208 401
rect 211 399 213 401
rect 216 399 218 401
rect 221 399 223 401
rect 226 399 228 401
rect 231 399 233 401
rect 236 399 238 401
rect 241 399 243 401
rect 246 399 248 401
rect 251 399 253 401
rect 256 399 258 401
rect 261 399 263 401
rect 266 399 268 401
rect 271 399 273 401
rect 276 399 278 401
rect 281 399 283 401
rect 286 399 288 401
rect 291 399 293 401
rect 296 399 298 401
rect 301 399 303 401
rect 306 399 308 401
rect 311 399 313 401
rect 316 399 318 401
rect 333 399 335 401
rect 338 399 340 401
rect 2 395 4 397
rect 7 395 9 397
rect 33 396 35 398
rect 162 396 164 398
rect 196 396 198 398
rect 325 396 327 398
rect 20 394 22 396
rect 25 394 27 396
rect 42 394 44 396
rect 47 394 49 396
rect 52 394 54 396
rect 57 394 59 396
rect 62 394 64 396
rect 67 394 69 396
rect 72 394 74 396
rect 77 394 79 396
rect 82 394 84 396
rect 87 394 89 396
rect 92 394 94 396
rect 97 394 99 396
rect 102 394 104 396
rect 107 394 109 396
rect 112 394 114 396
rect 117 394 119 396
rect 122 394 124 396
rect 127 394 129 396
rect 132 394 134 396
rect 137 394 139 396
rect 142 394 144 396
rect 147 394 149 396
rect 152 394 154 396
rect 177 394 179 396
rect 182 394 184 396
rect 206 394 208 396
rect 211 394 213 396
rect 216 394 218 396
rect 221 394 223 396
rect 226 394 228 396
rect 231 394 233 396
rect 236 394 238 396
rect 241 394 243 396
rect 246 394 248 396
rect 251 394 253 396
rect 256 394 258 396
rect 261 394 263 396
rect 266 394 268 396
rect 271 394 273 396
rect 276 394 278 396
rect 281 394 283 396
rect 286 394 288 396
rect 291 394 293 396
rect 296 394 298 396
rect 301 394 303 396
rect 306 394 308 396
rect 311 394 313 396
rect 316 394 318 396
rect 333 394 335 396
rect 338 394 340 396
rect 351 395 353 397
rect 356 395 358 397
rect 33 391 35 393
rect 162 391 164 393
rect 196 391 198 393
rect 325 391 327 393
rect 20 389 22 391
rect 25 389 27 391
rect 177 389 179 391
rect 182 389 184 391
rect 333 389 335 391
rect 338 389 340 391
rect 2 387 4 389
rect 7 387 9 389
rect 33 386 35 388
rect 162 386 164 388
rect 196 386 198 388
rect 325 386 327 388
rect 351 387 353 389
rect 356 387 358 389
rect 41 384 43 386
rect 51 384 53 386
rect 61 384 63 386
rect 71 384 73 386
rect 81 384 83 386
rect 91 384 93 386
rect 101 384 103 386
rect 111 384 113 386
rect 154 384 156 386
rect 204 384 206 386
rect 247 384 249 386
rect 257 384 259 386
rect 267 384 269 386
rect 277 384 279 386
rect 287 384 289 386
rect 297 384 299 386
rect 307 384 309 386
rect 317 384 319 386
rect 33 381 35 383
rect 162 381 164 383
rect 196 381 198 383
rect 325 381 327 383
rect 2 379 4 381
rect 7 379 9 381
rect 41 379 43 381
rect 51 379 53 381
rect 61 379 63 381
rect 71 379 73 381
rect 81 379 83 381
rect 91 379 93 381
rect 101 379 103 381
rect 111 379 113 381
rect 154 379 156 381
rect 204 379 206 381
rect 247 379 249 381
rect 257 379 259 381
rect 267 379 269 381
rect 277 379 279 381
rect 287 379 289 381
rect 297 379 299 381
rect 307 379 309 381
rect 317 379 319 381
rect 351 379 353 381
rect 356 379 358 381
rect 33 376 35 378
rect 162 376 164 378
rect 196 376 198 378
rect 325 376 327 378
rect 41 374 43 376
rect 51 374 53 376
rect 61 374 63 376
rect 71 374 73 376
rect 81 374 83 376
rect 91 374 93 376
rect 101 374 103 376
rect 111 374 113 376
rect 154 374 156 376
rect 204 374 206 376
rect 247 374 249 376
rect 257 374 259 376
rect 267 374 269 376
rect 277 374 279 376
rect 287 374 289 376
rect 297 374 299 376
rect 307 374 309 376
rect 317 374 319 376
rect 2 371 4 373
rect 7 371 9 373
rect 33 371 35 373
rect 162 371 164 373
rect 196 371 198 373
rect 325 371 327 373
rect 351 371 353 373
rect 356 371 358 373
rect 20 369 22 371
rect 25 369 27 371
rect 177 369 179 371
rect 182 369 184 371
rect 333 369 335 371
rect 338 369 340 371
rect 33 366 35 368
rect 162 366 164 368
rect 196 366 198 368
rect 325 366 327 368
rect 2 363 4 365
rect 7 363 9 365
rect 20 364 22 366
rect 25 364 27 366
rect 42 364 44 366
rect 47 364 49 366
rect 52 364 54 366
rect 57 364 59 366
rect 62 364 64 366
rect 67 364 69 366
rect 72 364 74 366
rect 77 364 79 366
rect 82 364 84 366
rect 87 364 89 366
rect 92 364 94 366
rect 97 364 99 366
rect 102 364 104 366
rect 107 364 109 366
rect 112 364 114 366
rect 117 364 119 366
rect 122 364 124 366
rect 127 364 129 366
rect 132 364 134 366
rect 137 364 139 366
rect 142 364 144 366
rect 147 364 149 366
rect 152 364 154 366
rect 177 364 179 366
rect 182 364 184 366
rect 206 364 208 366
rect 211 364 213 366
rect 216 364 218 366
rect 221 364 223 366
rect 226 364 228 366
rect 231 364 233 366
rect 236 364 238 366
rect 241 364 243 366
rect 246 364 248 366
rect 251 364 253 366
rect 256 364 258 366
rect 261 364 263 366
rect 266 364 268 366
rect 271 364 273 366
rect 276 364 278 366
rect 281 364 283 366
rect 286 364 288 366
rect 291 364 293 366
rect 296 364 298 366
rect 301 364 303 366
rect 306 364 308 366
rect 311 364 313 366
rect 316 364 318 366
rect 333 364 335 366
rect 338 364 340 366
rect 351 363 353 365
rect 356 363 358 365
rect 33 361 35 363
rect 162 361 164 363
rect 196 361 198 363
rect 325 361 327 363
rect 20 359 22 361
rect 25 359 27 361
rect 42 359 44 361
rect 47 359 49 361
rect 52 359 54 361
rect 57 359 59 361
rect 62 359 64 361
rect 67 359 69 361
rect 72 359 74 361
rect 77 359 79 361
rect 82 359 84 361
rect 87 359 89 361
rect 92 359 94 361
rect 97 359 99 361
rect 102 359 104 361
rect 107 359 109 361
rect 112 359 114 361
rect 117 359 119 361
rect 122 359 124 361
rect 127 359 129 361
rect 132 359 134 361
rect 137 359 139 361
rect 142 359 144 361
rect 147 359 149 361
rect 152 359 154 361
rect 177 359 179 361
rect 182 359 184 361
rect 206 359 208 361
rect 211 359 213 361
rect 216 359 218 361
rect 221 359 223 361
rect 226 359 228 361
rect 231 359 233 361
rect 236 359 238 361
rect 241 359 243 361
rect 246 359 248 361
rect 251 359 253 361
rect 256 359 258 361
rect 261 359 263 361
rect 266 359 268 361
rect 271 359 273 361
rect 276 359 278 361
rect 281 359 283 361
rect 286 359 288 361
rect 291 359 293 361
rect 296 359 298 361
rect 301 359 303 361
rect 306 359 308 361
rect 311 359 313 361
rect 316 359 318 361
rect 333 359 335 361
rect 338 359 340 361
rect 2 355 4 357
rect 7 355 9 357
rect 33 356 35 358
rect 162 356 164 358
rect 196 356 198 358
rect 325 356 327 358
rect 20 354 22 356
rect 25 354 27 356
rect 42 354 44 356
rect 47 354 49 356
rect 52 354 54 356
rect 57 354 59 356
rect 62 354 64 356
rect 67 354 69 356
rect 72 354 74 356
rect 77 354 79 356
rect 82 354 84 356
rect 87 354 89 356
rect 92 354 94 356
rect 97 354 99 356
rect 102 354 104 356
rect 107 354 109 356
rect 112 354 114 356
rect 117 354 119 356
rect 122 354 124 356
rect 127 354 129 356
rect 132 354 134 356
rect 137 354 139 356
rect 142 354 144 356
rect 147 354 149 356
rect 152 354 154 356
rect 177 354 179 356
rect 182 354 184 356
rect 206 354 208 356
rect 211 354 213 356
rect 216 354 218 356
rect 221 354 223 356
rect 226 354 228 356
rect 231 354 233 356
rect 236 354 238 356
rect 241 354 243 356
rect 246 354 248 356
rect 251 354 253 356
rect 256 354 258 356
rect 261 354 263 356
rect 266 354 268 356
rect 271 354 273 356
rect 276 354 278 356
rect 281 354 283 356
rect 286 354 288 356
rect 291 354 293 356
rect 296 354 298 356
rect 301 354 303 356
rect 306 354 308 356
rect 311 354 313 356
rect 316 354 318 356
rect 333 354 335 356
rect 338 354 340 356
rect 351 355 353 357
rect 356 355 358 357
rect 33 351 35 353
rect 162 351 164 353
rect 196 351 198 353
rect 325 351 327 353
rect 20 349 22 351
rect 25 349 27 351
rect 42 349 44 351
rect 47 349 49 351
rect 52 349 54 351
rect 57 349 59 351
rect 62 349 64 351
rect 67 349 69 351
rect 72 349 74 351
rect 77 349 79 351
rect 82 349 84 351
rect 87 349 89 351
rect 92 349 94 351
rect 97 349 99 351
rect 102 349 104 351
rect 107 349 109 351
rect 112 349 114 351
rect 117 349 119 351
rect 122 349 124 351
rect 127 349 129 351
rect 132 349 134 351
rect 137 349 139 351
rect 142 349 144 351
rect 147 349 149 351
rect 152 349 154 351
rect 177 349 179 351
rect 182 349 184 351
rect 206 349 208 351
rect 211 349 213 351
rect 216 349 218 351
rect 221 349 223 351
rect 226 349 228 351
rect 231 349 233 351
rect 236 349 238 351
rect 241 349 243 351
rect 246 349 248 351
rect 251 349 253 351
rect 256 349 258 351
rect 261 349 263 351
rect 266 349 268 351
rect 271 349 273 351
rect 276 349 278 351
rect 281 349 283 351
rect 286 349 288 351
rect 291 349 293 351
rect 296 349 298 351
rect 301 349 303 351
rect 306 349 308 351
rect 311 349 313 351
rect 316 349 318 351
rect 333 349 335 351
rect 338 349 340 351
rect 2 347 4 349
rect 7 347 9 349
rect 351 347 353 349
rect 356 347 358 349
rect 20 344 22 346
rect 25 344 27 346
rect 33 345 35 347
rect 42 344 44 346
rect 47 344 49 346
rect 52 344 54 346
rect 57 344 59 346
rect 62 344 64 346
rect 67 344 69 346
rect 72 344 74 346
rect 77 344 79 346
rect 82 344 84 346
rect 87 344 89 346
rect 92 344 94 346
rect 97 344 99 346
rect 102 344 104 346
rect 107 344 109 346
rect 112 344 114 346
rect 117 344 119 346
rect 122 344 124 346
rect 127 344 129 346
rect 132 344 134 346
rect 137 344 139 346
rect 142 344 144 346
rect 147 344 149 346
rect 152 344 154 346
rect 162 345 164 347
rect 177 344 179 346
rect 182 344 184 346
rect 196 345 198 347
rect 206 344 208 346
rect 211 344 213 346
rect 216 344 218 346
rect 221 344 223 346
rect 226 344 228 346
rect 231 344 233 346
rect 236 344 238 346
rect 241 344 243 346
rect 246 344 248 346
rect 251 344 253 346
rect 256 344 258 346
rect 261 344 263 346
rect 266 344 268 346
rect 271 344 273 346
rect 276 344 278 346
rect 281 344 283 346
rect 286 344 288 346
rect 291 344 293 346
rect 296 344 298 346
rect 301 344 303 346
rect 306 344 308 346
rect 311 344 313 346
rect 316 344 318 346
rect 325 345 327 347
rect 333 344 335 346
rect 338 344 340 346
rect 2 339 4 341
rect 7 339 9 341
rect 20 339 22 341
rect 25 339 27 341
rect 33 340 35 342
rect 42 339 44 341
rect 47 339 49 341
rect 52 339 54 341
rect 57 339 59 341
rect 62 339 64 341
rect 67 339 69 341
rect 72 339 74 341
rect 77 339 79 341
rect 82 339 84 341
rect 87 339 89 341
rect 92 339 94 341
rect 97 339 99 341
rect 102 339 104 341
rect 107 339 109 341
rect 112 339 114 341
rect 117 339 119 341
rect 122 339 124 341
rect 127 339 129 341
rect 132 339 134 341
rect 137 339 139 341
rect 142 339 144 341
rect 147 339 149 341
rect 152 339 154 341
rect 162 340 164 342
rect 177 339 179 341
rect 182 339 184 341
rect 196 340 198 342
rect 206 339 208 341
rect 211 339 213 341
rect 216 339 218 341
rect 221 339 223 341
rect 226 339 228 341
rect 231 339 233 341
rect 236 339 238 341
rect 241 339 243 341
rect 246 339 248 341
rect 251 339 253 341
rect 256 339 258 341
rect 261 339 263 341
rect 266 339 268 341
rect 271 339 273 341
rect 276 339 278 341
rect 281 339 283 341
rect 286 339 288 341
rect 291 339 293 341
rect 296 339 298 341
rect 301 339 303 341
rect 306 339 308 341
rect 311 339 313 341
rect 316 339 318 341
rect 325 340 327 342
rect 333 339 335 341
rect 338 339 340 341
rect 351 339 353 341
rect 356 339 358 341
rect 20 334 22 336
rect 25 334 27 336
rect 33 335 35 337
rect 42 334 44 336
rect 47 334 49 336
rect 52 334 54 336
rect 57 334 59 336
rect 62 334 64 336
rect 67 334 69 336
rect 72 334 74 336
rect 77 334 79 336
rect 82 334 84 336
rect 87 334 89 336
rect 92 334 94 336
rect 97 334 99 336
rect 102 334 104 336
rect 107 334 109 336
rect 112 334 114 336
rect 117 334 119 336
rect 122 334 124 336
rect 127 334 129 336
rect 132 334 134 336
rect 137 334 139 336
rect 142 334 144 336
rect 147 334 149 336
rect 152 334 154 336
rect 162 335 164 337
rect 177 334 179 336
rect 182 334 184 336
rect 196 335 198 337
rect 206 334 208 336
rect 211 334 213 336
rect 216 334 218 336
rect 221 334 223 336
rect 226 334 228 336
rect 231 334 233 336
rect 236 334 238 336
rect 241 334 243 336
rect 246 334 248 336
rect 251 334 253 336
rect 256 334 258 336
rect 261 334 263 336
rect 266 334 268 336
rect 271 334 273 336
rect 276 334 278 336
rect 281 334 283 336
rect 286 334 288 336
rect 291 334 293 336
rect 296 334 298 336
rect 301 334 303 336
rect 306 334 308 336
rect 311 334 313 336
rect 316 334 318 336
rect 325 335 327 337
rect 333 334 335 336
rect 338 334 340 336
rect 2 330 4 332
rect 7 330 9 332
rect 20 329 22 331
rect 25 329 27 331
rect 33 330 35 332
rect 42 329 44 331
rect 47 329 49 331
rect 52 329 54 331
rect 57 329 59 331
rect 62 329 64 331
rect 67 329 69 331
rect 72 329 74 331
rect 77 329 79 331
rect 82 329 84 331
rect 87 329 89 331
rect 92 329 94 331
rect 97 329 99 331
rect 102 329 104 331
rect 107 329 109 331
rect 112 329 114 331
rect 117 329 119 331
rect 122 329 124 331
rect 127 329 129 331
rect 132 329 134 331
rect 137 329 139 331
rect 142 329 144 331
rect 147 329 149 331
rect 152 329 154 331
rect 162 330 164 332
rect 177 329 179 331
rect 182 329 184 331
rect 196 330 198 332
rect 206 329 208 331
rect 211 329 213 331
rect 216 329 218 331
rect 221 329 223 331
rect 226 329 228 331
rect 231 329 233 331
rect 236 329 238 331
rect 241 329 243 331
rect 246 329 248 331
rect 251 329 253 331
rect 256 329 258 331
rect 261 329 263 331
rect 266 329 268 331
rect 271 329 273 331
rect 276 329 278 331
rect 281 329 283 331
rect 286 329 288 331
rect 291 329 293 331
rect 296 329 298 331
rect 301 329 303 331
rect 306 329 308 331
rect 311 329 313 331
rect 316 329 318 331
rect 325 330 327 332
rect 333 329 335 331
rect 338 329 340 331
rect 351 330 353 332
rect 356 330 358 332
rect 20 324 22 326
rect 25 324 27 326
rect 33 325 35 327
rect 162 325 164 327
rect 177 324 179 326
rect 182 324 184 326
rect 196 325 198 327
rect 325 325 327 327
rect 333 324 335 326
rect 338 324 340 326
rect 2 322 4 324
rect 7 322 9 324
rect 351 322 353 324
rect 356 322 358 324
rect 33 320 35 322
rect 41 319 43 321
rect 51 319 53 321
rect 61 319 63 321
rect 71 319 73 321
rect 81 319 83 321
rect 91 319 93 321
rect 101 319 103 321
rect 111 319 113 321
rect 154 319 156 321
rect 162 320 164 322
rect 196 320 198 322
rect 204 319 206 321
rect 247 319 249 321
rect 257 319 259 321
rect 267 319 269 321
rect 277 319 279 321
rect 287 319 289 321
rect 297 319 299 321
rect 307 319 309 321
rect 317 319 319 321
rect 325 320 327 322
rect 2 314 4 316
rect 7 314 9 316
rect 33 315 35 317
rect 41 314 43 316
rect 51 314 53 316
rect 61 314 63 316
rect 71 314 73 316
rect 81 314 83 316
rect 91 314 93 316
rect 101 314 103 316
rect 111 314 113 316
rect 154 314 156 316
rect 162 315 164 317
rect 196 315 198 317
rect 204 314 206 316
rect 247 314 249 316
rect 257 314 259 316
rect 267 314 269 316
rect 277 314 279 316
rect 287 314 289 316
rect 297 314 299 316
rect 307 314 309 316
rect 317 314 319 316
rect 325 315 327 317
rect 351 314 353 316
rect 356 314 358 316
rect 33 310 35 312
rect 41 309 43 311
rect 51 309 53 311
rect 61 309 63 311
rect 71 309 73 311
rect 81 309 83 311
rect 91 309 93 311
rect 101 309 103 311
rect 111 309 113 311
rect 154 309 156 311
rect 162 310 164 312
rect 196 310 198 312
rect 204 309 206 311
rect 247 309 249 311
rect 257 309 259 311
rect 267 309 269 311
rect 277 309 279 311
rect 287 309 289 311
rect 297 309 299 311
rect 307 309 309 311
rect 317 309 319 311
rect 325 310 327 312
rect 2 306 4 308
rect 7 306 9 308
rect 20 304 22 306
rect 25 304 27 306
rect 33 305 35 307
rect 162 305 164 307
rect 177 304 179 306
rect 182 304 184 306
rect 196 305 198 307
rect 325 305 327 307
rect 351 306 353 308
rect 356 306 358 308
rect 333 304 335 306
rect 338 304 340 306
rect 2 298 4 300
rect 7 298 9 300
rect 20 299 22 301
rect 25 299 27 301
rect 33 300 35 302
rect 42 299 44 301
rect 47 299 49 301
rect 52 299 54 301
rect 57 299 59 301
rect 62 299 64 301
rect 67 299 69 301
rect 72 299 74 301
rect 77 299 79 301
rect 82 299 84 301
rect 87 299 89 301
rect 92 299 94 301
rect 97 299 99 301
rect 102 299 104 301
rect 107 299 109 301
rect 112 299 114 301
rect 117 299 119 301
rect 122 299 124 301
rect 127 299 129 301
rect 132 299 134 301
rect 137 299 139 301
rect 142 299 144 301
rect 147 299 149 301
rect 152 299 154 301
rect 162 300 164 302
rect 177 299 179 301
rect 182 299 184 301
rect 196 300 198 302
rect 206 299 208 301
rect 211 299 213 301
rect 216 299 218 301
rect 221 299 223 301
rect 226 299 228 301
rect 231 299 233 301
rect 236 299 238 301
rect 241 299 243 301
rect 246 299 248 301
rect 251 299 253 301
rect 256 299 258 301
rect 261 299 263 301
rect 266 299 268 301
rect 271 299 273 301
rect 276 299 278 301
rect 281 299 283 301
rect 286 299 288 301
rect 291 299 293 301
rect 296 299 298 301
rect 301 299 303 301
rect 306 299 308 301
rect 311 299 313 301
rect 316 299 318 301
rect 325 300 327 302
rect 333 299 335 301
rect 338 299 340 301
rect 351 298 353 300
rect 356 298 358 300
rect 20 294 22 296
rect 25 294 27 296
rect 33 295 35 297
rect 42 294 44 296
rect 47 294 49 296
rect 52 294 54 296
rect 57 294 59 296
rect 62 294 64 296
rect 67 294 69 296
rect 72 294 74 296
rect 77 294 79 296
rect 82 294 84 296
rect 87 294 89 296
rect 92 294 94 296
rect 97 294 99 296
rect 102 294 104 296
rect 107 294 109 296
rect 112 294 114 296
rect 117 294 119 296
rect 122 294 124 296
rect 127 294 129 296
rect 132 294 134 296
rect 137 294 139 296
rect 142 294 144 296
rect 147 294 149 296
rect 152 294 154 296
rect 162 295 164 297
rect 177 294 179 296
rect 182 294 184 296
rect 196 295 198 297
rect 206 294 208 296
rect 211 294 213 296
rect 216 294 218 296
rect 221 294 223 296
rect 226 294 228 296
rect 231 294 233 296
rect 236 294 238 296
rect 241 294 243 296
rect 246 294 248 296
rect 251 294 253 296
rect 256 294 258 296
rect 261 294 263 296
rect 266 294 268 296
rect 271 294 273 296
rect 276 294 278 296
rect 281 294 283 296
rect 286 294 288 296
rect 291 294 293 296
rect 296 294 298 296
rect 301 294 303 296
rect 306 294 308 296
rect 311 294 313 296
rect 316 294 318 296
rect 325 295 327 297
rect 333 294 335 296
rect 338 294 340 296
rect 2 290 4 292
rect 7 290 9 292
rect 20 289 22 291
rect 25 289 27 291
rect 33 290 35 292
rect 42 289 44 291
rect 47 289 49 291
rect 52 289 54 291
rect 57 289 59 291
rect 62 289 64 291
rect 67 289 69 291
rect 72 289 74 291
rect 77 289 79 291
rect 82 289 84 291
rect 87 289 89 291
rect 92 289 94 291
rect 97 289 99 291
rect 102 289 104 291
rect 107 289 109 291
rect 112 289 114 291
rect 117 289 119 291
rect 122 289 124 291
rect 127 289 129 291
rect 132 289 134 291
rect 137 289 139 291
rect 142 289 144 291
rect 147 289 149 291
rect 152 289 154 291
rect 162 290 164 292
rect 177 289 179 291
rect 182 289 184 291
rect 196 290 198 292
rect 206 289 208 291
rect 211 289 213 291
rect 216 289 218 291
rect 221 289 223 291
rect 226 289 228 291
rect 231 289 233 291
rect 236 289 238 291
rect 241 289 243 291
rect 246 289 248 291
rect 251 289 253 291
rect 256 289 258 291
rect 261 289 263 291
rect 266 289 268 291
rect 271 289 273 291
rect 276 289 278 291
rect 281 289 283 291
rect 286 289 288 291
rect 291 289 293 291
rect 296 289 298 291
rect 301 289 303 291
rect 306 289 308 291
rect 311 289 313 291
rect 316 289 318 291
rect 325 290 327 292
rect 333 289 335 291
rect 338 289 340 291
rect 351 290 353 292
rect 356 290 358 292
rect 20 284 22 286
rect 25 284 27 286
rect 33 285 35 287
rect 42 284 44 286
rect 47 284 49 286
rect 52 284 54 286
rect 57 284 59 286
rect 62 284 64 286
rect 67 284 69 286
rect 72 284 74 286
rect 77 284 79 286
rect 82 284 84 286
rect 87 284 89 286
rect 92 284 94 286
rect 97 284 99 286
rect 102 284 104 286
rect 107 284 109 286
rect 112 284 114 286
rect 117 284 119 286
rect 122 284 124 286
rect 127 284 129 286
rect 132 284 134 286
rect 137 284 139 286
rect 142 284 144 286
rect 147 284 149 286
rect 152 284 154 286
rect 162 285 164 287
rect 177 284 179 286
rect 182 284 184 286
rect 196 285 198 287
rect 206 284 208 286
rect 211 284 213 286
rect 216 284 218 286
rect 221 284 223 286
rect 226 284 228 286
rect 231 284 233 286
rect 236 284 238 286
rect 241 284 243 286
rect 246 284 248 286
rect 251 284 253 286
rect 256 284 258 286
rect 261 284 263 286
rect 266 284 268 286
rect 271 284 273 286
rect 276 284 278 286
rect 281 284 283 286
rect 286 284 288 286
rect 291 284 293 286
rect 296 284 298 286
rect 301 284 303 286
rect 306 284 308 286
rect 311 284 313 286
rect 316 284 318 286
rect 325 285 327 287
rect 333 284 335 286
rect 338 284 340 286
rect 2 282 4 284
rect 7 282 9 284
rect 351 282 353 284
rect 356 282 358 284
rect 20 279 22 281
rect 25 279 27 281
rect 33 280 35 282
rect 42 279 44 281
rect 47 279 49 281
rect 52 279 54 281
rect 57 279 59 281
rect 62 279 64 281
rect 67 279 69 281
rect 72 279 74 281
rect 77 279 79 281
rect 82 279 84 281
rect 87 279 89 281
rect 92 279 94 281
rect 97 279 99 281
rect 102 279 104 281
rect 107 279 109 281
rect 112 279 114 281
rect 117 279 119 281
rect 122 279 124 281
rect 127 279 129 281
rect 132 279 134 281
rect 137 279 139 281
rect 142 279 144 281
rect 147 279 149 281
rect 152 279 154 281
rect 162 280 164 282
rect 177 279 179 281
rect 182 279 184 281
rect 196 280 198 282
rect 206 279 208 281
rect 211 279 213 281
rect 216 279 218 281
rect 221 279 223 281
rect 226 279 228 281
rect 231 279 233 281
rect 236 279 238 281
rect 241 279 243 281
rect 246 279 248 281
rect 251 279 253 281
rect 256 279 258 281
rect 261 279 263 281
rect 266 279 268 281
rect 271 279 273 281
rect 276 279 278 281
rect 281 279 283 281
rect 286 279 288 281
rect 291 279 293 281
rect 296 279 298 281
rect 301 279 303 281
rect 306 279 308 281
rect 311 279 313 281
rect 316 279 318 281
rect 325 280 327 282
rect 333 279 335 281
rect 338 279 340 281
rect 2 274 4 276
rect 7 274 9 276
rect 20 274 22 276
rect 25 274 27 276
rect 33 275 35 277
rect 42 274 44 276
rect 47 274 49 276
rect 52 274 54 276
rect 57 274 59 276
rect 62 274 64 276
rect 67 274 69 276
rect 72 274 74 276
rect 77 274 79 276
rect 82 274 84 276
rect 87 274 89 276
rect 92 274 94 276
rect 97 274 99 276
rect 102 274 104 276
rect 107 274 109 276
rect 112 274 114 276
rect 117 274 119 276
rect 122 274 124 276
rect 127 274 129 276
rect 132 274 134 276
rect 137 274 139 276
rect 142 274 144 276
rect 147 274 149 276
rect 152 274 154 276
rect 162 275 164 277
rect 177 274 179 276
rect 182 274 184 276
rect 196 275 198 277
rect 206 274 208 276
rect 211 274 213 276
rect 216 274 218 276
rect 221 274 223 276
rect 226 274 228 276
rect 231 274 233 276
rect 236 274 238 276
rect 241 274 243 276
rect 246 274 248 276
rect 251 274 253 276
rect 256 274 258 276
rect 261 274 263 276
rect 266 274 268 276
rect 271 274 273 276
rect 276 274 278 276
rect 281 274 283 276
rect 286 274 288 276
rect 291 274 293 276
rect 296 274 298 276
rect 301 274 303 276
rect 306 274 308 276
rect 311 274 313 276
rect 316 274 318 276
rect 325 275 327 277
rect 333 274 335 276
rect 338 274 340 276
rect 351 274 353 276
rect 356 274 358 276
rect 20 269 22 271
rect 25 269 27 271
rect 33 270 35 272
rect 42 269 44 271
rect 47 269 49 271
rect 52 269 54 271
rect 57 269 59 271
rect 62 269 64 271
rect 67 269 69 271
rect 72 269 74 271
rect 77 269 79 271
rect 82 269 84 271
rect 87 269 89 271
rect 92 269 94 271
rect 97 269 99 271
rect 102 269 104 271
rect 107 269 109 271
rect 112 269 114 271
rect 117 269 119 271
rect 122 269 124 271
rect 127 269 129 271
rect 132 269 134 271
rect 137 269 139 271
rect 142 269 144 271
rect 147 269 149 271
rect 152 269 154 271
rect 162 270 164 272
rect 177 269 179 271
rect 182 269 184 271
rect 196 270 198 272
rect 206 269 208 271
rect 211 269 213 271
rect 216 269 218 271
rect 221 269 223 271
rect 226 269 228 271
rect 231 269 233 271
rect 236 269 238 271
rect 241 269 243 271
rect 246 269 248 271
rect 251 269 253 271
rect 256 269 258 271
rect 261 269 263 271
rect 266 269 268 271
rect 271 269 273 271
rect 276 269 278 271
rect 281 269 283 271
rect 286 269 288 271
rect 291 269 293 271
rect 296 269 298 271
rect 301 269 303 271
rect 306 269 308 271
rect 311 269 313 271
rect 316 269 318 271
rect 325 270 327 272
rect 333 269 335 271
rect 338 269 340 271
rect 2 266 4 268
rect 7 266 9 268
rect 20 264 22 266
rect 25 264 27 266
rect 33 265 35 267
rect 42 264 44 266
rect 47 264 49 266
rect 52 264 54 266
rect 57 264 59 266
rect 62 264 64 266
rect 67 264 69 266
rect 72 264 74 266
rect 77 264 79 266
rect 82 264 84 266
rect 87 264 89 266
rect 92 264 94 266
rect 97 264 99 266
rect 102 264 104 266
rect 107 264 109 266
rect 112 264 114 266
rect 117 264 119 266
rect 122 264 124 266
rect 127 264 129 266
rect 132 264 134 266
rect 137 264 139 266
rect 142 264 144 266
rect 147 264 149 266
rect 152 264 154 266
rect 162 265 164 267
rect 177 264 179 266
rect 182 264 184 266
rect 196 265 198 267
rect 206 264 208 266
rect 211 264 213 266
rect 216 264 218 266
rect 221 264 223 266
rect 226 264 228 266
rect 231 264 233 266
rect 236 264 238 266
rect 241 264 243 266
rect 246 264 248 266
rect 251 264 253 266
rect 256 264 258 266
rect 261 264 263 266
rect 266 264 268 266
rect 271 264 273 266
rect 276 264 278 266
rect 281 264 283 266
rect 286 264 288 266
rect 291 264 293 266
rect 296 264 298 266
rect 301 264 303 266
rect 306 264 308 266
rect 311 264 313 266
rect 316 264 318 266
rect 325 265 327 267
rect 351 266 353 268
rect 356 266 358 268
rect 333 264 335 266
rect 338 264 340 266
rect 2 258 4 260
rect 7 258 9 260
rect 20 259 22 261
rect 25 259 27 261
rect 33 260 35 262
rect 162 260 164 262
rect 177 259 179 261
rect 182 259 184 261
rect 196 260 198 262
rect 325 260 327 262
rect 333 259 335 261
rect 338 259 340 261
rect 351 258 353 260
rect 356 258 358 260
rect 41 254 43 256
rect 51 254 53 256
rect 61 254 63 256
rect 71 254 73 256
rect 81 254 83 256
rect 91 254 93 256
rect 101 254 103 256
rect 111 254 113 256
rect 154 254 156 256
rect 204 254 206 256
rect 247 254 249 256
rect 257 254 259 256
rect 267 254 269 256
rect 277 254 279 256
rect 287 254 289 256
rect 297 254 299 256
rect 307 254 309 256
rect 317 254 319 256
rect 2 250 4 252
rect 7 250 9 252
rect 41 249 43 251
rect 51 249 53 251
rect 61 249 63 251
rect 71 249 73 251
rect 81 249 83 251
rect 91 249 93 251
rect 101 249 103 251
rect 111 249 113 251
rect 154 249 156 251
rect 204 249 206 251
rect 247 249 249 251
rect 257 249 259 251
rect 267 249 269 251
rect 277 249 279 251
rect 287 249 289 251
rect 297 249 299 251
rect 307 249 309 251
rect 317 249 319 251
rect 351 250 353 252
rect 356 250 358 252
rect 41 244 43 246
rect 51 244 53 246
rect 61 244 63 246
rect 71 244 73 246
rect 81 244 83 246
rect 91 244 93 246
rect 101 244 103 246
rect 111 244 113 246
rect 154 244 156 246
rect 204 244 206 246
rect 247 244 249 246
rect 257 244 259 246
rect 267 244 269 246
rect 277 244 279 246
rect 287 244 289 246
rect 297 244 299 246
rect 307 244 309 246
rect 317 244 319 246
rect 2 242 4 244
rect 7 242 9 244
rect 351 242 353 244
rect 356 242 358 244
rect 2 234 4 236
rect 7 234 9 236
rect 351 234 353 236
rect 356 234 358 236
rect 9 226 11 228
rect 17 226 19 228
rect 25 226 27 228
rect 41 226 43 228
rect 49 226 51 228
rect 57 226 59 228
rect 65 226 67 228
rect 73 226 75 228
rect 81 226 83 228
rect 89 226 91 228
rect 97 226 99 228
rect 105 226 107 228
rect 113 226 115 228
rect 153 226 155 228
rect 177 226 179 228
rect 205 226 207 228
rect 245 226 247 228
rect 253 226 255 228
rect 261 226 263 228
rect 269 226 271 228
rect 277 226 279 228
rect 285 226 287 228
rect 293 226 295 228
rect 301 226 303 228
rect 309 226 311 228
rect 317 226 319 228
rect 333 226 335 228
rect 341 226 343 228
rect 349 226 351 228
rect 9 221 11 223
rect 17 221 19 223
rect 25 221 27 223
rect 41 221 43 223
rect 49 221 51 223
rect 57 221 59 223
rect 65 221 67 223
rect 73 221 75 223
rect 81 221 83 223
rect 89 221 91 223
rect 97 221 99 223
rect 105 221 107 223
rect 113 221 115 223
rect 153 221 155 223
rect 177 221 179 223
rect 205 221 207 223
rect 245 221 247 223
rect 253 221 255 223
rect 261 221 263 223
rect 269 221 271 223
rect 277 221 279 223
rect 285 221 287 223
rect 293 221 295 223
rect 301 221 303 223
rect 309 221 311 223
rect 317 221 319 223
rect 333 221 335 223
rect 341 221 343 223
rect 349 221 351 223
rect 9 209 11 211
rect 17 209 19 211
rect 25 209 27 211
rect 41 209 43 211
rect 49 209 51 211
rect 57 209 59 211
rect 65 209 67 211
rect 73 209 75 211
rect 81 209 83 211
rect 89 209 91 211
rect 97 209 99 211
rect 105 209 107 211
rect 113 209 115 211
rect 153 209 155 211
rect 177 209 179 211
rect 205 209 207 211
rect 245 209 247 211
rect 253 209 255 211
rect 261 209 263 211
rect 269 209 271 211
rect 277 209 279 211
rect 285 209 287 211
rect 293 209 295 211
rect 301 209 303 211
rect 309 209 311 211
rect 317 209 319 211
rect 333 209 335 211
rect 341 209 343 211
rect 349 209 351 211
rect 9 204 11 206
rect 17 204 19 206
rect 25 204 27 206
rect 41 204 43 206
rect 49 204 51 206
rect 57 204 59 206
rect 65 204 67 206
rect 73 204 75 206
rect 81 204 83 206
rect 89 204 91 206
rect 97 204 99 206
rect 105 204 107 206
rect 113 204 115 206
rect 153 204 155 206
rect 177 204 179 206
rect 205 204 207 206
rect 245 204 247 206
rect 253 204 255 206
rect 261 204 263 206
rect 269 204 271 206
rect 277 204 279 206
rect 285 204 287 206
rect 293 204 295 206
rect 301 204 303 206
rect 309 204 311 206
rect 317 204 319 206
rect 333 204 335 206
rect 341 204 343 206
rect 349 204 351 206
rect 86 167 88 169
rect 91 167 93 169
rect 96 167 98 169
rect 101 167 103 169
rect 106 167 108 169
rect 111 167 113 169
rect 116 167 118 169
rect 121 167 123 169
rect 126 167 128 169
rect 131 167 133 169
rect 136 167 138 169
rect 141 167 143 169
rect 146 167 148 169
rect 151 167 153 169
rect 156 167 158 169
rect 161 167 163 169
rect 166 167 168 169
rect 171 167 173 169
rect 176 167 178 169
rect 181 167 183 169
rect 186 167 188 169
rect 191 167 193 169
rect 196 167 198 169
rect 201 167 203 169
rect 206 167 208 169
rect 211 167 213 169
rect 216 167 218 169
rect 221 167 223 169
rect 226 167 228 169
rect 231 167 233 169
rect 236 167 238 169
rect 241 167 243 169
rect 246 167 248 169
rect 251 167 253 169
rect 256 167 258 169
rect 261 167 263 169
rect 266 167 268 169
rect 271 167 273 169
rect 276 167 278 169
rect 86 162 88 164
rect 91 162 93 164
rect 96 162 98 164
rect 101 162 103 164
rect 106 162 108 164
rect 111 162 113 164
rect 116 162 118 164
rect 121 162 123 164
rect 126 162 128 164
rect 131 162 133 164
rect 136 162 138 164
rect 141 162 143 164
rect 146 162 148 164
rect 151 162 153 164
rect 156 162 158 164
rect 161 162 163 164
rect 166 162 168 164
rect 171 162 173 164
rect 176 162 178 164
rect 181 162 183 164
rect 186 162 188 164
rect 191 162 193 164
rect 196 162 198 164
rect 201 162 203 164
rect 206 162 208 164
rect 211 162 213 164
rect 216 162 218 164
rect 221 162 223 164
rect 226 162 228 164
rect 231 162 233 164
rect 236 162 238 164
rect 241 162 243 164
rect 246 162 248 164
rect 251 162 253 164
rect 256 162 258 164
rect 261 162 263 164
rect 266 162 268 164
rect 271 162 273 164
rect 276 162 278 164
rect 86 132 88 134
rect 91 132 93 134
rect 96 132 98 134
rect 101 132 103 134
rect 106 132 108 134
rect 111 132 113 134
rect 116 132 118 134
rect 121 132 123 134
rect 126 132 128 134
rect 131 132 133 134
rect 136 132 138 134
rect 141 132 143 134
rect 146 132 148 134
rect 151 132 153 134
rect 156 132 158 134
rect 161 132 163 134
rect 166 132 168 134
rect 171 132 173 134
rect 176 132 178 134
rect 181 132 183 134
rect 186 132 188 134
rect 191 132 193 134
rect 196 132 198 134
rect 201 132 203 134
rect 206 132 208 134
rect 211 132 213 134
rect 216 132 218 134
rect 221 132 223 134
rect 226 132 228 134
rect 231 132 233 134
rect 236 132 238 134
rect 241 132 243 134
rect 246 132 248 134
rect 251 132 253 134
rect 256 132 258 134
rect 261 132 263 134
rect 266 132 268 134
rect 271 132 273 134
rect 276 132 278 134
rect 86 127 88 129
rect 91 127 93 129
rect 96 127 98 129
rect 101 127 103 129
rect 106 127 108 129
rect 111 127 113 129
rect 116 127 118 129
rect 121 127 123 129
rect 126 127 128 129
rect 131 127 133 129
rect 136 127 138 129
rect 141 127 143 129
rect 146 127 148 129
rect 151 127 153 129
rect 156 127 158 129
rect 161 127 163 129
rect 166 127 168 129
rect 171 127 173 129
rect 176 127 178 129
rect 181 127 183 129
rect 186 127 188 129
rect 191 127 193 129
rect 196 127 198 129
rect 201 127 203 129
rect 206 127 208 129
rect 211 127 213 129
rect 216 127 218 129
rect 221 127 223 129
rect 226 127 228 129
rect 231 127 233 129
rect 236 127 238 129
rect 241 127 243 129
rect 246 127 248 129
rect 251 127 253 129
rect 256 127 258 129
rect 261 127 263 129
rect 266 127 268 129
rect 271 127 273 129
rect 276 127 278 129
rect 7 96 9 98
rect 41 96 43 98
rect 49 96 51 98
rect 57 96 59 98
rect 65 96 67 98
rect 73 96 75 98
rect 81 96 83 98
rect 89 96 91 98
rect 97 96 99 98
rect 105 96 107 98
rect 113 96 115 98
rect 121 96 123 98
rect 129 96 131 98
rect 137 96 139 98
rect 145 96 147 98
rect 153 96 155 98
rect 161 96 163 98
rect 197 96 199 98
rect 205 96 207 98
rect 213 96 215 98
rect 221 96 223 98
rect 229 96 231 98
rect 237 96 239 98
rect 245 96 247 98
rect 253 96 255 98
rect 261 96 263 98
rect 269 96 271 98
rect 277 96 279 98
rect 285 96 287 98
rect 293 96 295 98
rect 301 96 303 98
rect 309 96 311 98
rect 317 96 319 98
rect 351 96 353 98
rect 7 91 9 93
rect 41 91 43 93
rect 49 91 51 93
rect 57 91 59 93
rect 65 91 67 93
rect 73 91 75 93
rect 81 91 83 93
rect 89 91 91 93
rect 97 91 99 93
rect 105 91 107 93
rect 113 91 115 93
rect 121 91 123 93
rect 129 91 131 93
rect 137 91 139 93
rect 145 91 147 93
rect 153 91 155 93
rect 161 91 163 93
rect 197 91 199 93
rect 205 91 207 93
rect 213 91 215 93
rect 221 91 223 93
rect 229 91 231 93
rect 237 91 239 93
rect 245 91 247 93
rect 253 91 255 93
rect 261 91 263 93
rect 269 91 271 93
rect 277 91 279 93
rect 285 91 287 93
rect 293 91 295 93
rect 301 91 303 93
rect 309 91 311 93
rect 317 91 319 93
rect 351 91 353 93
<< metal1 >>
rect 45 856 315 1126
rect 62 816 298 856
rect 102 806 258 816
rect 112 796 248 806
rect 120 793 240 796
rect 0 773 117 784
rect 0 538 11 773
rect 18 745 115 761
rect 18 550 29 745
rect 0 527 29 538
rect 0 510 29 521
rect 32 506 36 742
rect 120 740 143 793
rect 149 773 211 784
rect 168 765 192 769
rect 148 745 164 761
rect 41 701 165 740
rect 39 680 115 696
rect 120 675 143 701
rect 148 680 164 696
rect 41 636 165 675
rect 39 615 115 631
rect 120 610 143 636
rect 148 615 164 631
rect 41 571 165 610
rect 39 550 115 566
rect 39 527 117 538
rect 39 510 117 521
rect 31 497 42 506
rect 0 482 117 493
rect 0 465 117 476
rect 0 230 11 465
rect 18 437 115 453
rect 18 242 29 437
rect 0 219 29 230
rect 0 202 29 213
rect 0 89 11 202
rect 32 198 36 434
rect 120 432 143 571
rect 148 550 164 566
rect 168 546 172 765
rect 175 550 185 761
rect 188 546 192 765
rect 196 745 212 761
rect 217 740 240 793
rect 243 773 360 784
rect 245 745 342 761
rect 195 701 319 740
rect 196 680 212 696
rect 217 675 240 701
rect 245 680 321 696
rect 195 636 319 675
rect 196 615 212 631
rect 217 610 240 636
rect 245 615 321 631
rect 195 571 319 610
rect 196 550 212 566
rect 168 542 192 546
rect 148 527 162 538
rect 148 510 162 521
rect 168 506 172 542
rect 175 527 185 538
rect 175 510 185 521
rect 188 506 192 542
rect 196 527 210 538
rect 196 510 210 521
rect 167 497 193 506
rect 148 482 162 493
rect 148 465 162 476
rect 168 461 172 497
rect 175 482 185 493
rect 175 465 185 476
rect 188 461 192 497
rect 196 482 210 493
rect 196 465 210 476
rect 168 457 192 461
rect 148 437 157 453
rect 41 393 155 432
rect 39 372 115 388
rect 120 367 143 393
rect 148 372 157 388
rect 41 328 155 367
rect 39 307 115 323
rect 120 302 143 328
rect 148 307 157 323
rect 41 263 155 302
rect 39 242 115 258
rect 39 219 116 230
rect 39 202 117 213
rect 15 189 42 198
rect 120 189 143 263
rect 148 242 157 258
rect 148 219 156 230
rect 148 202 156 213
rect 161 198 165 436
rect 155 189 165 198
rect 15 89 19 189
rect 117 186 143 189
rect 111 183 143 186
rect 168 184 172 457
rect 175 242 185 453
rect 176 219 184 230
rect 176 202 184 213
rect 188 184 192 457
rect 203 437 212 453
rect 195 198 199 436
rect 217 432 240 571
rect 245 550 321 566
rect 243 527 321 538
rect 243 510 321 521
rect 324 506 328 742
rect 331 550 342 745
rect 349 538 360 773
rect 331 527 360 538
rect 331 510 360 521
rect 318 497 329 506
rect 243 482 360 493
rect 243 465 360 476
rect 245 437 342 453
rect 205 393 319 432
rect 203 372 212 388
rect 217 367 240 393
rect 245 372 321 388
rect 205 328 319 367
rect 203 307 212 323
rect 217 302 240 328
rect 245 307 321 323
rect 205 263 319 302
rect 203 242 212 258
rect 204 219 212 230
rect 204 202 212 213
rect 195 189 205 198
rect 217 189 240 263
rect 245 242 321 258
rect 244 219 321 230
rect 243 202 321 213
rect 324 198 328 434
rect 331 242 342 437
rect 349 230 360 465
rect 331 219 360 230
rect 331 202 360 213
rect 318 189 329 198
rect 217 186 243 189
rect 105 180 146 183
rect 99 177 152 180
rect 93 174 158 177
rect 167 175 193 184
rect 217 183 249 186
rect 214 180 255 183
rect 208 177 261 180
rect 202 174 267 177
rect 318 175 345 184
rect 87 171 163 174
rect 197 171 273 174
rect 81 160 279 171
rect 81 125 279 136
rect 87 122 273 125
rect 99 119 261 122
rect 111 116 249 119
rect 123 113 237 116
rect 135 110 225 113
rect 147 107 213 110
rect 159 104 201 107
rect 23 89 170 100
rect 175 89 187 104
rect 192 89 321 100
rect 341 89 345 175
rect 349 89 360 202
rect 0 82 11 85
rect 8 79 11 82
rect 15 48 19 85
rect 23 82 170 85
rect 235 82 337 85
rect 39 79 170 82
rect 82 66 84 68
rect 341 48 345 85
rect 349 79 360 85
rect 15 44 25 48
rect 335 44 345 48
rect 8 3 23 6
rect 40 3 360 6
rect 0 0 360 3
<< metal2 >>
rect 47 858 313 1124
rect 0 773 360 784
rect 0 745 360 761
rect 0 707 360 734
rect 0 680 360 696
rect 0 647 360 674
rect 0 615 360 631
rect 0 582 360 609
rect 0 550 360 566
rect 0 527 360 538
rect 0 510 360 521
rect 31 497 329 506
rect 0 482 360 493
rect 0 465 360 476
rect 0 437 360 453
rect 0 399 360 426
rect 0 372 360 388
rect 0 339 360 366
rect 0 307 360 323
rect 0 274 360 301
rect 0 242 360 258
rect 0 219 360 230
rect 0 202 360 213
rect 31 189 329 198
rect 167 175 329 184
rect -16 89 360 100
rect -16 6 -8 89
rect 0 79 360 85
rect 95 72 168 76
rect 41 65 85 69
rect 41 55 45 65
rect 95 62 99 72
rect 206 65 265 69
rect 261 62 265 65
rect 104 58 256 62
rect 104 51 108 58
rect 118 51 242 55
rect 252 51 256 58
rect 84 44 116 48
rect 245 44 276 48
rect 315 41 319 51
rect 276 37 319 41
rect -16 0 360 6
<< gv1 >>
rect 59 1110 61 1112
rect 69 1110 71 1112
rect 79 1110 81 1112
rect 89 1110 91 1112
rect 99 1110 101 1112
rect 109 1110 111 1112
rect 119 1110 121 1112
rect 129 1110 131 1112
rect 139 1110 141 1112
rect 149 1110 151 1112
rect 159 1110 161 1112
rect 169 1110 171 1112
rect 179 1110 181 1112
rect 189 1110 191 1112
rect 199 1110 201 1112
rect 209 1110 211 1112
rect 219 1110 221 1112
rect 229 1110 231 1112
rect 239 1110 241 1112
rect 249 1110 251 1112
rect 259 1110 261 1112
rect 269 1110 271 1112
rect 279 1110 281 1112
rect 289 1110 291 1112
rect 299 1110 301 1112
rect 59 1100 61 1102
rect 69 1100 71 1102
rect 79 1100 81 1102
rect 89 1100 91 1102
rect 99 1100 101 1102
rect 109 1100 111 1102
rect 119 1100 121 1102
rect 129 1100 131 1102
rect 139 1100 141 1102
rect 149 1100 151 1102
rect 159 1100 161 1102
rect 169 1100 171 1102
rect 179 1100 181 1102
rect 189 1100 191 1102
rect 199 1100 201 1102
rect 209 1100 211 1102
rect 219 1100 221 1102
rect 229 1100 231 1102
rect 239 1100 241 1102
rect 249 1100 251 1102
rect 259 1100 261 1102
rect 269 1100 271 1102
rect 279 1100 281 1102
rect 289 1100 291 1102
rect 299 1100 301 1102
rect 59 1090 61 1092
rect 69 1090 71 1092
rect 79 1090 81 1092
rect 89 1090 91 1092
rect 99 1090 101 1092
rect 109 1090 111 1092
rect 119 1090 121 1092
rect 129 1090 131 1092
rect 139 1090 141 1092
rect 149 1090 151 1092
rect 159 1090 161 1092
rect 169 1090 171 1092
rect 179 1090 181 1092
rect 189 1090 191 1092
rect 199 1090 201 1092
rect 209 1090 211 1092
rect 219 1090 221 1092
rect 229 1090 231 1092
rect 239 1090 241 1092
rect 249 1090 251 1092
rect 259 1090 261 1092
rect 269 1090 271 1092
rect 279 1090 281 1092
rect 289 1090 291 1092
rect 299 1090 301 1092
rect 59 1080 61 1082
rect 69 1080 71 1082
rect 79 1080 81 1082
rect 89 1080 91 1082
rect 99 1080 101 1082
rect 109 1080 111 1082
rect 119 1080 121 1082
rect 129 1080 131 1082
rect 139 1080 141 1082
rect 149 1080 151 1082
rect 159 1080 161 1082
rect 169 1080 171 1082
rect 179 1080 181 1082
rect 189 1080 191 1082
rect 199 1080 201 1082
rect 209 1080 211 1082
rect 219 1080 221 1082
rect 229 1080 231 1082
rect 239 1080 241 1082
rect 249 1080 251 1082
rect 259 1080 261 1082
rect 269 1080 271 1082
rect 279 1080 281 1082
rect 289 1080 291 1082
rect 299 1080 301 1082
rect 59 1070 61 1072
rect 69 1070 71 1072
rect 79 1070 81 1072
rect 89 1070 91 1072
rect 99 1070 101 1072
rect 109 1070 111 1072
rect 119 1070 121 1072
rect 129 1070 131 1072
rect 139 1070 141 1072
rect 149 1070 151 1072
rect 159 1070 161 1072
rect 169 1070 171 1072
rect 179 1070 181 1072
rect 189 1070 191 1072
rect 199 1070 201 1072
rect 209 1070 211 1072
rect 219 1070 221 1072
rect 229 1070 231 1072
rect 239 1070 241 1072
rect 249 1070 251 1072
rect 259 1070 261 1072
rect 269 1070 271 1072
rect 279 1070 281 1072
rect 289 1070 291 1072
rect 299 1070 301 1072
rect 59 1060 61 1062
rect 69 1060 71 1062
rect 79 1060 81 1062
rect 89 1060 91 1062
rect 99 1060 101 1062
rect 109 1060 111 1062
rect 119 1060 121 1062
rect 129 1060 131 1062
rect 139 1060 141 1062
rect 149 1060 151 1062
rect 159 1060 161 1062
rect 169 1060 171 1062
rect 179 1060 181 1062
rect 189 1060 191 1062
rect 199 1060 201 1062
rect 209 1060 211 1062
rect 219 1060 221 1062
rect 229 1060 231 1062
rect 239 1060 241 1062
rect 249 1060 251 1062
rect 259 1060 261 1062
rect 269 1060 271 1062
rect 279 1060 281 1062
rect 289 1060 291 1062
rect 299 1060 301 1062
rect 59 1050 61 1052
rect 69 1050 71 1052
rect 79 1050 81 1052
rect 89 1050 91 1052
rect 99 1050 101 1052
rect 109 1050 111 1052
rect 119 1050 121 1052
rect 129 1050 131 1052
rect 139 1050 141 1052
rect 149 1050 151 1052
rect 159 1050 161 1052
rect 169 1050 171 1052
rect 179 1050 181 1052
rect 189 1050 191 1052
rect 199 1050 201 1052
rect 209 1050 211 1052
rect 219 1050 221 1052
rect 229 1050 231 1052
rect 239 1050 241 1052
rect 249 1050 251 1052
rect 259 1050 261 1052
rect 269 1050 271 1052
rect 279 1050 281 1052
rect 289 1050 291 1052
rect 299 1050 301 1052
rect 59 1040 61 1042
rect 69 1040 71 1042
rect 79 1040 81 1042
rect 89 1040 91 1042
rect 99 1040 101 1042
rect 109 1040 111 1042
rect 119 1040 121 1042
rect 129 1040 131 1042
rect 139 1040 141 1042
rect 149 1040 151 1042
rect 159 1040 161 1042
rect 169 1040 171 1042
rect 179 1040 181 1042
rect 189 1040 191 1042
rect 199 1040 201 1042
rect 209 1040 211 1042
rect 219 1040 221 1042
rect 229 1040 231 1042
rect 239 1040 241 1042
rect 249 1040 251 1042
rect 259 1040 261 1042
rect 269 1040 271 1042
rect 279 1040 281 1042
rect 289 1040 291 1042
rect 299 1040 301 1042
rect 59 1030 61 1032
rect 69 1030 71 1032
rect 79 1030 81 1032
rect 89 1030 91 1032
rect 99 1030 101 1032
rect 109 1030 111 1032
rect 119 1030 121 1032
rect 129 1030 131 1032
rect 139 1030 141 1032
rect 149 1030 151 1032
rect 159 1030 161 1032
rect 169 1030 171 1032
rect 179 1030 181 1032
rect 189 1030 191 1032
rect 199 1030 201 1032
rect 209 1030 211 1032
rect 219 1030 221 1032
rect 229 1030 231 1032
rect 239 1030 241 1032
rect 249 1030 251 1032
rect 259 1030 261 1032
rect 269 1030 271 1032
rect 279 1030 281 1032
rect 289 1030 291 1032
rect 299 1030 301 1032
rect 59 1020 61 1022
rect 69 1020 71 1022
rect 79 1020 81 1022
rect 89 1020 91 1022
rect 99 1020 101 1022
rect 109 1020 111 1022
rect 119 1020 121 1022
rect 129 1020 131 1022
rect 139 1020 141 1022
rect 149 1020 151 1022
rect 159 1020 161 1022
rect 169 1020 171 1022
rect 179 1020 181 1022
rect 189 1020 191 1022
rect 199 1020 201 1022
rect 209 1020 211 1022
rect 219 1020 221 1022
rect 229 1020 231 1022
rect 239 1020 241 1022
rect 249 1020 251 1022
rect 259 1020 261 1022
rect 269 1020 271 1022
rect 279 1020 281 1022
rect 289 1020 291 1022
rect 299 1020 301 1022
rect 59 1010 61 1012
rect 69 1010 71 1012
rect 79 1010 81 1012
rect 89 1010 91 1012
rect 99 1010 101 1012
rect 109 1010 111 1012
rect 119 1010 121 1012
rect 129 1010 131 1012
rect 139 1010 141 1012
rect 149 1010 151 1012
rect 159 1010 161 1012
rect 169 1010 171 1012
rect 179 1010 181 1012
rect 189 1010 191 1012
rect 199 1010 201 1012
rect 209 1010 211 1012
rect 219 1010 221 1012
rect 229 1010 231 1012
rect 239 1010 241 1012
rect 249 1010 251 1012
rect 259 1010 261 1012
rect 269 1010 271 1012
rect 279 1010 281 1012
rect 289 1010 291 1012
rect 299 1010 301 1012
rect 59 1000 61 1002
rect 69 1000 71 1002
rect 79 1000 81 1002
rect 89 1000 91 1002
rect 99 1000 101 1002
rect 109 1000 111 1002
rect 119 1000 121 1002
rect 129 1000 131 1002
rect 139 1000 141 1002
rect 149 1000 151 1002
rect 159 1000 161 1002
rect 169 1000 171 1002
rect 179 1000 181 1002
rect 189 1000 191 1002
rect 199 1000 201 1002
rect 209 1000 211 1002
rect 219 1000 221 1002
rect 229 1000 231 1002
rect 239 1000 241 1002
rect 249 1000 251 1002
rect 259 1000 261 1002
rect 269 1000 271 1002
rect 279 1000 281 1002
rect 289 1000 291 1002
rect 299 1000 301 1002
rect 59 990 61 992
rect 69 990 71 992
rect 79 990 81 992
rect 89 990 91 992
rect 99 990 101 992
rect 109 990 111 992
rect 119 990 121 992
rect 129 990 131 992
rect 139 990 141 992
rect 149 990 151 992
rect 159 990 161 992
rect 169 990 171 992
rect 179 990 181 992
rect 189 990 191 992
rect 199 990 201 992
rect 209 990 211 992
rect 219 990 221 992
rect 229 990 231 992
rect 239 990 241 992
rect 249 990 251 992
rect 259 990 261 992
rect 269 990 271 992
rect 279 990 281 992
rect 289 990 291 992
rect 299 990 301 992
rect 59 980 61 982
rect 69 980 71 982
rect 79 980 81 982
rect 89 980 91 982
rect 99 980 101 982
rect 109 980 111 982
rect 119 980 121 982
rect 129 980 131 982
rect 139 980 141 982
rect 149 980 151 982
rect 159 980 161 982
rect 169 980 171 982
rect 179 980 181 982
rect 189 980 191 982
rect 199 980 201 982
rect 209 980 211 982
rect 219 980 221 982
rect 229 980 231 982
rect 239 980 241 982
rect 249 980 251 982
rect 259 980 261 982
rect 269 980 271 982
rect 279 980 281 982
rect 289 980 291 982
rect 299 980 301 982
rect 59 970 61 972
rect 69 970 71 972
rect 79 970 81 972
rect 89 970 91 972
rect 99 970 101 972
rect 109 970 111 972
rect 119 970 121 972
rect 129 970 131 972
rect 139 970 141 972
rect 149 970 151 972
rect 159 970 161 972
rect 169 970 171 972
rect 179 970 181 972
rect 189 970 191 972
rect 199 970 201 972
rect 209 970 211 972
rect 219 970 221 972
rect 229 970 231 972
rect 239 970 241 972
rect 249 970 251 972
rect 259 970 261 972
rect 269 970 271 972
rect 279 970 281 972
rect 289 970 291 972
rect 299 970 301 972
rect 59 960 61 962
rect 69 960 71 962
rect 79 960 81 962
rect 89 960 91 962
rect 99 960 101 962
rect 109 960 111 962
rect 119 960 121 962
rect 129 960 131 962
rect 139 960 141 962
rect 149 960 151 962
rect 159 960 161 962
rect 169 960 171 962
rect 179 960 181 962
rect 189 960 191 962
rect 199 960 201 962
rect 209 960 211 962
rect 219 960 221 962
rect 229 960 231 962
rect 239 960 241 962
rect 249 960 251 962
rect 259 960 261 962
rect 269 960 271 962
rect 279 960 281 962
rect 289 960 291 962
rect 299 960 301 962
rect 59 950 61 952
rect 69 950 71 952
rect 79 950 81 952
rect 89 950 91 952
rect 99 950 101 952
rect 109 950 111 952
rect 119 950 121 952
rect 129 950 131 952
rect 139 950 141 952
rect 149 950 151 952
rect 159 950 161 952
rect 169 950 171 952
rect 179 950 181 952
rect 189 950 191 952
rect 199 950 201 952
rect 209 950 211 952
rect 219 950 221 952
rect 229 950 231 952
rect 239 950 241 952
rect 249 950 251 952
rect 259 950 261 952
rect 269 950 271 952
rect 279 950 281 952
rect 289 950 291 952
rect 299 950 301 952
rect 59 940 61 942
rect 69 940 71 942
rect 79 940 81 942
rect 89 940 91 942
rect 99 940 101 942
rect 109 940 111 942
rect 119 940 121 942
rect 129 940 131 942
rect 139 940 141 942
rect 149 940 151 942
rect 159 940 161 942
rect 169 940 171 942
rect 179 940 181 942
rect 189 940 191 942
rect 199 940 201 942
rect 209 940 211 942
rect 219 940 221 942
rect 229 940 231 942
rect 239 940 241 942
rect 249 940 251 942
rect 259 940 261 942
rect 269 940 271 942
rect 279 940 281 942
rect 289 940 291 942
rect 299 940 301 942
rect 59 930 61 932
rect 69 930 71 932
rect 79 930 81 932
rect 89 930 91 932
rect 99 930 101 932
rect 109 930 111 932
rect 119 930 121 932
rect 129 930 131 932
rect 139 930 141 932
rect 149 930 151 932
rect 159 930 161 932
rect 169 930 171 932
rect 179 930 181 932
rect 189 930 191 932
rect 199 930 201 932
rect 209 930 211 932
rect 219 930 221 932
rect 229 930 231 932
rect 239 930 241 932
rect 249 930 251 932
rect 259 930 261 932
rect 269 930 271 932
rect 279 930 281 932
rect 289 930 291 932
rect 299 930 301 932
rect 59 920 61 922
rect 69 920 71 922
rect 79 920 81 922
rect 89 920 91 922
rect 99 920 101 922
rect 109 920 111 922
rect 119 920 121 922
rect 129 920 131 922
rect 139 920 141 922
rect 149 920 151 922
rect 159 920 161 922
rect 169 920 171 922
rect 179 920 181 922
rect 189 920 191 922
rect 199 920 201 922
rect 209 920 211 922
rect 219 920 221 922
rect 229 920 231 922
rect 239 920 241 922
rect 249 920 251 922
rect 259 920 261 922
rect 269 920 271 922
rect 279 920 281 922
rect 289 920 291 922
rect 299 920 301 922
rect 59 910 61 912
rect 69 910 71 912
rect 79 910 81 912
rect 89 910 91 912
rect 99 910 101 912
rect 109 910 111 912
rect 119 910 121 912
rect 129 910 131 912
rect 139 910 141 912
rect 149 910 151 912
rect 159 910 161 912
rect 169 910 171 912
rect 179 910 181 912
rect 189 910 191 912
rect 199 910 201 912
rect 209 910 211 912
rect 219 910 221 912
rect 229 910 231 912
rect 239 910 241 912
rect 249 910 251 912
rect 259 910 261 912
rect 269 910 271 912
rect 279 910 281 912
rect 289 910 291 912
rect 299 910 301 912
rect 59 900 61 902
rect 69 900 71 902
rect 79 900 81 902
rect 89 900 91 902
rect 99 900 101 902
rect 109 900 111 902
rect 119 900 121 902
rect 129 900 131 902
rect 139 900 141 902
rect 149 900 151 902
rect 159 900 161 902
rect 169 900 171 902
rect 179 900 181 902
rect 189 900 191 902
rect 199 900 201 902
rect 209 900 211 902
rect 219 900 221 902
rect 229 900 231 902
rect 239 900 241 902
rect 249 900 251 902
rect 259 900 261 902
rect 269 900 271 902
rect 279 900 281 902
rect 289 900 291 902
rect 299 900 301 902
rect 59 890 61 892
rect 69 890 71 892
rect 79 890 81 892
rect 89 890 91 892
rect 99 890 101 892
rect 109 890 111 892
rect 119 890 121 892
rect 129 890 131 892
rect 139 890 141 892
rect 149 890 151 892
rect 159 890 161 892
rect 169 890 171 892
rect 179 890 181 892
rect 189 890 191 892
rect 199 890 201 892
rect 209 890 211 892
rect 219 890 221 892
rect 229 890 231 892
rect 239 890 241 892
rect 249 890 251 892
rect 259 890 261 892
rect 269 890 271 892
rect 279 890 281 892
rect 289 890 291 892
rect 299 890 301 892
rect 59 880 61 882
rect 69 880 71 882
rect 79 880 81 882
rect 89 880 91 882
rect 99 880 101 882
rect 109 880 111 882
rect 119 880 121 882
rect 129 880 131 882
rect 139 880 141 882
rect 149 880 151 882
rect 159 880 161 882
rect 169 880 171 882
rect 179 880 181 882
rect 189 880 191 882
rect 199 880 201 882
rect 209 880 211 882
rect 219 880 221 882
rect 229 880 231 882
rect 239 880 241 882
rect 249 880 251 882
rect 259 880 261 882
rect 269 880 271 882
rect 279 880 281 882
rect 289 880 291 882
rect 299 880 301 882
rect 59 870 61 872
rect 69 870 71 872
rect 79 870 81 872
rect 89 870 91 872
rect 99 870 101 872
rect 109 870 111 872
rect 119 870 121 872
rect 129 870 131 872
rect 139 870 141 872
rect 149 870 151 872
rect 159 870 161 872
rect 169 870 171 872
rect 179 870 181 872
rect 189 870 191 872
rect 199 870 201 872
rect 209 870 211 872
rect 219 870 221 872
rect 229 870 231 872
rect 239 870 241 872
rect 249 870 251 872
rect 259 870 261 872
rect 269 870 271 872
rect 279 870 281 872
rect 289 870 291 872
rect 299 870 301 872
rect 5 780 7 782
rect 13 780 15 782
rect 21 780 23 782
rect 29 780 31 782
rect 37 780 39 782
rect 45 780 47 782
rect 53 780 55 782
rect 61 780 63 782
rect 69 780 71 782
rect 77 780 79 782
rect 85 780 87 782
rect 93 780 95 782
rect 101 780 103 782
rect 109 780 111 782
rect 155 780 157 782
rect 163 780 165 782
rect 171 780 173 782
rect 179 780 181 782
rect 187 780 189 782
rect 195 780 197 782
rect 203 780 205 782
rect 249 780 251 782
rect 257 780 259 782
rect 265 780 267 782
rect 273 780 275 782
rect 281 780 283 782
rect 289 780 291 782
rect 297 780 299 782
rect 305 780 307 782
rect 313 780 315 782
rect 321 780 323 782
rect 329 780 331 782
rect 337 780 339 782
rect 345 780 347 782
rect 353 780 355 782
rect 5 775 7 777
rect 13 775 15 777
rect 21 775 23 777
rect 29 775 31 777
rect 37 775 39 777
rect 45 775 47 777
rect 53 775 55 777
rect 61 775 63 777
rect 69 775 71 777
rect 77 775 79 777
rect 85 775 87 777
rect 93 775 95 777
rect 101 775 103 777
rect 109 775 111 777
rect 155 775 157 777
rect 163 775 165 777
rect 171 775 173 777
rect 179 775 181 777
rect 187 775 189 777
rect 195 775 197 777
rect 203 775 205 777
rect 249 775 251 777
rect 257 775 259 777
rect 265 775 267 777
rect 273 775 275 777
rect 281 775 283 777
rect 289 775 291 777
rect 297 775 299 777
rect 305 775 307 777
rect 313 775 315 777
rect 321 775 323 777
rect 329 775 331 777
rect 337 775 339 777
rect 345 775 347 777
rect 353 775 355 777
rect 20 757 22 759
rect 25 757 27 759
rect 35 757 37 759
rect 46 757 48 759
rect 56 757 58 759
rect 66 757 68 759
rect 76 757 78 759
rect 86 757 88 759
rect 96 757 98 759
rect 106 757 108 759
rect 155 757 157 759
rect 177 757 179 759
rect 182 757 184 759
rect 203 757 205 759
rect 252 757 254 759
rect 262 757 264 759
rect 272 757 274 759
rect 282 757 284 759
rect 292 757 294 759
rect 302 757 304 759
rect 312 757 314 759
rect 322 757 324 759
rect 332 757 335 759
rect 338 757 340 759
rect 20 752 22 754
rect 25 752 27 754
rect 35 752 37 754
rect 46 752 48 754
rect 56 752 58 754
rect 66 752 68 754
rect 76 752 78 754
rect 86 752 88 754
rect 96 752 98 754
rect 106 752 108 754
rect 155 752 157 754
rect 177 752 179 754
rect 182 752 184 754
rect 203 752 205 754
rect 252 752 254 754
rect 262 752 264 754
rect 272 752 274 754
rect 282 752 284 754
rect 292 752 294 754
rect 302 752 304 754
rect 312 752 314 754
rect 322 752 324 754
rect 333 752 335 754
rect 338 752 340 754
rect 20 747 22 749
rect 25 747 27 749
rect 35 747 37 749
rect 46 747 48 749
rect 56 747 58 749
rect 66 747 68 749
rect 76 747 78 749
rect 86 747 88 749
rect 96 747 98 749
rect 106 747 108 749
rect 155 747 157 749
rect 177 747 179 749
rect 182 747 184 749
rect 203 747 205 749
rect 252 747 254 749
rect 262 747 264 749
rect 272 747 274 749
rect 282 747 284 749
rect 292 747 294 749
rect 302 747 304 749
rect 312 747 314 749
rect 322 747 324 749
rect 333 747 335 749
rect 338 747 340 749
rect 2 731 4 733
rect 7 731 9 733
rect 351 731 353 733
rect 356 731 358 733
rect 2 723 4 725
rect 7 723 9 725
rect 351 723 353 725
rect 356 723 358 725
rect 2 715 4 717
rect 7 715 9 717
rect 351 715 353 717
rect 356 715 358 717
rect 20 692 22 694
rect 25 692 27 694
rect 46 692 48 694
rect 56 692 58 694
rect 66 692 68 694
rect 76 692 78 694
rect 86 692 88 694
rect 96 692 98 694
rect 106 692 108 694
rect 155 692 157 694
rect 177 692 179 694
rect 182 692 184 694
rect 203 692 205 694
rect 252 692 254 694
rect 262 692 264 694
rect 272 692 274 694
rect 282 692 284 694
rect 292 692 294 694
rect 302 692 304 694
rect 312 692 314 694
rect 333 692 335 694
rect 338 692 340 694
rect 20 687 22 689
rect 25 687 27 689
rect 46 687 48 689
rect 56 687 58 689
rect 66 687 68 689
rect 76 687 78 689
rect 86 687 88 689
rect 96 687 98 689
rect 106 687 108 689
rect 155 687 157 689
rect 177 687 179 689
rect 182 687 184 689
rect 203 687 205 689
rect 252 687 254 689
rect 262 687 264 689
rect 272 687 274 689
rect 282 687 284 689
rect 292 687 294 689
rect 302 687 304 689
rect 312 687 314 689
rect 333 687 335 689
rect 338 687 340 689
rect 20 682 22 684
rect 25 682 27 684
rect 46 682 48 684
rect 56 682 58 684
rect 66 682 68 684
rect 76 682 78 684
rect 86 682 88 684
rect 96 682 98 684
rect 106 682 108 684
rect 155 682 157 684
rect 177 682 179 684
rect 182 682 184 684
rect 203 682 205 684
rect 252 682 254 684
rect 262 682 264 684
rect 272 682 274 684
rect 282 682 284 684
rect 292 682 294 684
rect 302 682 304 684
rect 312 682 314 684
rect 333 682 335 684
rect 338 682 340 684
rect 2 667 4 669
rect 7 667 9 669
rect 351 667 353 669
rect 356 667 358 669
rect 2 659 4 661
rect 7 659 9 661
rect 351 659 353 661
rect 356 659 358 661
rect 2 651 4 653
rect 7 651 9 653
rect 351 651 353 653
rect 356 651 358 653
rect 20 627 22 629
rect 25 627 27 629
rect 46 627 48 629
rect 56 627 58 629
rect 66 627 68 629
rect 76 627 78 629
rect 86 627 88 629
rect 96 627 98 629
rect 106 627 108 629
rect 155 627 157 629
rect 177 627 179 629
rect 182 627 184 629
rect 203 627 205 629
rect 252 627 254 629
rect 262 627 264 629
rect 272 627 274 629
rect 282 627 284 629
rect 292 627 294 629
rect 302 627 304 629
rect 312 627 314 629
rect 333 627 335 629
rect 338 627 340 629
rect 20 622 22 624
rect 25 622 27 624
rect 46 622 48 624
rect 56 622 58 624
rect 66 622 68 624
rect 76 622 78 624
rect 86 622 88 624
rect 96 622 98 624
rect 106 622 108 624
rect 155 622 157 624
rect 177 622 179 624
rect 182 622 184 624
rect 203 622 205 624
rect 252 622 254 624
rect 262 622 264 624
rect 272 622 274 624
rect 282 622 284 624
rect 292 622 294 624
rect 302 622 304 624
rect 312 622 314 624
rect 333 622 335 624
rect 338 622 340 624
rect 20 617 22 619
rect 25 617 27 619
rect 46 617 48 619
rect 56 617 58 619
rect 66 617 68 619
rect 76 617 78 619
rect 86 617 88 619
rect 96 617 98 619
rect 106 617 108 619
rect 155 617 157 619
rect 177 617 179 619
rect 182 617 184 619
rect 203 617 205 619
rect 252 617 254 619
rect 262 617 264 619
rect 272 617 274 619
rect 282 617 284 619
rect 292 617 294 619
rect 302 617 304 619
rect 312 617 314 619
rect 333 617 335 619
rect 338 617 340 619
rect 2 602 4 604
rect 7 602 9 604
rect 351 602 353 604
rect 356 602 358 604
rect 2 594 4 596
rect 7 594 9 596
rect 351 594 353 596
rect 356 594 358 596
rect 2 586 4 588
rect 7 586 9 588
rect 351 586 353 588
rect 356 586 358 588
rect 20 562 22 564
rect 25 562 27 564
rect 46 562 48 564
rect 56 562 58 564
rect 66 562 68 564
rect 76 562 78 564
rect 86 562 88 564
rect 96 562 98 564
rect 106 562 108 564
rect 155 562 157 564
rect 177 562 179 564
rect 182 562 184 564
rect 203 562 205 564
rect 252 562 254 564
rect 262 562 264 564
rect 272 562 274 564
rect 282 562 284 564
rect 292 562 294 564
rect 302 562 304 564
rect 312 562 314 564
rect 333 562 335 564
rect 338 562 340 564
rect 20 557 22 559
rect 25 557 27 559
rect 46 557 48 559
rect 56 557 58 559
rect 66 557 68 559
rect 76 557 78 559
rect 86 557 88 559
rect 96 557 98 559
rect 106 557 108 559
rect 155 557 157 559
rect 177 557 179 559
rect 182 557 184 559
rect 203 557 205 559
rect 252 557 254 559
rect 262 557 264 559
rect 272 557 274 559
rect 282 557 284 559
rect 292 557 294 559
rect 302 557 304 559
rect 312 557 314 559
rect 333 557 335 559
rect 338 557 340 559
rect 20 552 22 554
rect 25 552 27 554
rect 46 552 48 554
rect 56 552 58 554
rect 66 552 68 554
rect 76 552 78 554
rect 86 552 88 554
rect 96 552 98 554
rect 106 552 108 554
rect 155 552 157 554
rect 177 552 179 554
rect 182 552 184 554
rect 203 552 205 554
rect 252 552 254 554
rect 262 552 264 554
rect 272 552 274 554
rect 282 552 284 554
rect 292 552 294 554
rect 302 552 304 554
rect 312 552 314 554
rect 333 552 335 554
rect 338 552 340 554
rect 5 534 7 536
rect 13 534 15 536
rect 21 534 23 536
rect 45 534 47 536
rect 53 534 55 536
rect 61 534 63 536
rect 69 534 71 536
rect 77 534 79 536
rect 85 534 87 536
rect 93 534 95 536
rect 101 534 103 536
rect 109 534 111 536
rect 154 534 156 536
rect 177 534 179 536
rect 202 534 204 536
rect 249 534 251 536
rect 257 534 259 536
rect 265 534 267 536
rect 273 534 275 536
rect 281 534 283 536
rect 289 534 291 536
rect 297 534 299 536
rect 305 534 307 536
rect 313 534 315 536
rect 337 534 339 536
rect 345 534 347 536
rect 353 534 355 536
rect 5 529 7 531
rect 13 529 15 531
rect 21 529 23 531
rect 45 529 47 531
rect 53 529 55 531
rect 61 529 63 531
rect 69 529 71 531
rect 77 529 79 531
rect 85 529 87 531
rect 93 529 95 531
rect 101 529 103 531
rect 109 529 111 531
rect 154 529 156 531
rect 177 529 179 531
rect 202 529 204 531
rect 249 529 251 531
rect 257 529 259 531
rect 265 529 267 531
rect 273 529 275 531
rect 281 529 283 531
rect 289 529 291 531
rect 297 529 299 531
rect 305 529 307 531
rect 313 529 315 531
rect 337 529 339 531
rect 345 529 347 531
rect 353 529 355 531
rect 5 517 7 519
rect 13 517 15 519
rect 21 517 23 519
rect 45 517 47 519
rect 53 517 55 519
rect 61 517 63 519
rect 69 517 71 519
rect 77 517 79 519
rect 85 517 87 519
rect 93 517 95 519
rect 101 517 103 519
rect 109 517 111 519
rect 154 517 156 519
rect 177 517 179 519
rect 202 517 204 519
rect 249 517 251 519
rect 257 517 259 519
rect 265 517 267 519
rect 273 517 275 519
rect 281 517 283 519
rect 289 517 291 519
rect 297 517 299 519
rect 305 517 307 519
rect 313 517 315 519
rect 337 517 339 519
rect 345 517 347 519
rect 353 517 355 519
rect 5 512 7 514
rect 13 512 15 514
rect 21 512 23 514
rect 45 512 47 514
rect 53 512 55 514
rect 61 512 63 514
rect 69 512 71 514
rect 77 512 79 514
rect 85 512 87 514
rect 93 512 95 514
rect 101 512 103 514
rect 109 512 111 514
rect 154 512 156 514
rect 177 512 179 514
rect 202 512 204 514
rect 249 512 251 514
rect 257 512 259 514
rect 265 512 267 514
rect 273 512 275 514
rect 281 512 283 514
rect 289 512 291 514
rect 297 512 299 514
rect 305 512 307 514
rect 313 512 315 514
rect 337 512 339 514
rect 345 512 347 514
rect 353 512 355 514
rect 33 503 35 505
rect 38 503 40 505
rect 169 503 171 505
rect 174 503 176 505
rect 179 503 181 505
rect 184 503 186 505
rect 189 503 191 505
rect 320 503 322 505
rect 325 503 327 505
rect 33 498 35 500
rect 38 498 40 500
rect 169 498 171 500
rect 174 498 176 500
rect 179 498 181 500
rect 184 498 186 500
rect 189 498 191 500
rect 320 498 322 500
rect 325 498 327 500
rect 5 489 7 491
rect 13 489 15 491
rect 21 489 23 491
rect 29 489 31 491
rect 37 489 39 491
rect 45 489 47 491
rect 53 489 55 491
rect 61 489 63 491
rect 69 489 71 491
rect 77 489 79 491
rect 85 489 87 491
rect 93 489 95 491
rect 101 489 103 491
rect 109 489 111 491
rect 154 489 156 491
rect 177 489 179 491
rect 202 489 204 491
rect 249 489 251 491
rect 257 489 259 491
rect 265 489 267 491
rect 273 489 275 491
rect 281 489 283 491
rect 289 489 291 491
rect 297 489 299 491
rect 305 489 307 491
rect 313 489 315 491
rect 321 489 323 491
rect 329 489 331 491
rect 337 489 339 491
rect 345 489 347 491
rect 353 489 355 491
rect 5 484 7 486
rect 13 484 15 486
rect 21 484 23 486
rect 29 484 31 486
rect 37 484 39 486
rect 45 484 47 486
rect 53 484 55 486
rect 61 484 63 486
rect 69 484 71 486
rect 77 484 79 486
rect 85 484 87 486
rect 93 484 95 486
rect 101 484 103 486
rect 109 484 111 486
rect 154 484 156 486
rect 177 484 179 486
rect 202 484 204 486
rect 249 484 251 486
rect 257 484 259 486
rect 265 484 267 486
rect 273 484 275 486
rect 281 484 283 486
rect 289 484 291 486
rect 297 484 299 486
rect 305 484 307 486
rect 313 484 315 486
rect 321 484 323 486
rect 329 484 331 486
rect 337 484 339 486
rect 345 484 347 486
rect 353 484 355 486
rect 5 472 7 474
rect 13 472 15 474
rect 21 472 23 474
rect 29 472 31 474
rect 37 472 39 474
rect 45 472 47 474
rect 53 472 55 474
rect 61 472 63 474
rect 69 472 71 474
rect 77 472 79 474
rect 85 472 87 474
rect 93 472 95 474
rect 101 472 103 474
rect 109 472 111 474
rect 154 472 156 474
rect 177 472 179 474
rect 202 472 204 474
rect 249 472 251 474
rect 257 472 259 474
rect 265 472 267 474
rect 273 472 275 474
rect 281 472 283 474
rect 289 472 291 474
rect 297 472 299 474
rect 305 472 307 474
rect 313 472 315 474
rect 321 472 323 474
rect 329 472 331 474
rect 337 472 339 474
rect 345 472 347 474
rect 353 472 355 474
rect 5 467 7 469
rect 13 467 15 469
rect 21 467 23 469
rect 29 467 31 469
rect 37 467 39 469
rect 45 467 47 469
rect 53 467 55 469
rect 61 467 63 469
rect 69 467 71 469
rect 77 467 79 469
rect 85 467 87 469
rect 93 467 95 469
rect 101 467 103 469
rect 109 467 111 469
rect 154 467 156 469
rect 177 467 179 469
rect 202 467 204 469
rect 249 467 251 469
rect 257 467 259 469
rect 265 467 267 469
rect 273 467 275 469
rect 281 467 283 469
rect 289 467 291 469
rect 297 467 299 469
rect 305 467 307 469
rect 313 467 315 469
rect 321 467 323 469
rect 329 467 331 469
rect 337 467 339 469
rect 345 467 347 469
rect 353 467 355 469
rect 20 449 22 451
rect 25 449 27 451
rect 46 449 48 451
rect 56 449 58 451
rect 66 449 68 451
rect 76 449 78 451
rect 86 449 88 451
rect 96 449 98 451
rect 106 449 108 451
rect 149 449 151 451
rect 177 449 179 451
rect 182 449 184 451
rect 209 449 211 451
rect 252 449 254 451
rect 262 449 264 451
rect 272 449 274 451
rect 282 449 284 451
rect 292 449 294 451
rect 302 449 304 451
rect 312 449 314 451
rect 333 449 335 451
rect 338 449 340 451
rect 20 444 22 446
rect 25 444 27 446
rect 46 444 48 446
rect 56 444 58 446
rect 66 444 68 446
rect 76 444 78 446
rect 86 444 88 446
rect 96 444 98 446
rect 106 444 108 446
rect 149 444 151 446
rect 177 444 179 446
rect 182 444 184 446
rect 209 444 211 446
rect 252 444 254 446
rect 262 444 264 446
rect 272 444 274 446
rect 282 444 284 446
rect 292 444 294 446
rect 302 444 304 446
rect 312 444 314 446
rect 333 444 335 446
rect 338 444 340 446
rect 20 439 22 441
rect 25 439 27 441
rect 46 439 48 441
rect 56 439 58 441
rect 66 439 68 441
rect 76 439 78 441
rect 86 439 88 441
rect 96 439 98 441
rect 106 439 108 441
rect 149 439 151 441
rect 177 439 179 441
rect 182 439 184 441
rect 209 439 211 441
rect 252 439 254 441
rect 262 439 264 441
rect 272 439 274 441
rect 282 439 284 441
rect 292 439 294 441
rect 302 439 304 441
rect 312 439 314 441
rect 333 439 335 441
rect 338 439 340 441
rect 2 423 4 425
rect 7 423 9 425
rect 351 423 353 425
rect 356 423 358 425
rect 2 415 4 417
rect 7 415 9 417
rect 351 415 353 417
rect 356 415 358 417
rect 2 407 4 409
rect 7 407 9 409
rect 351 407 353 409
rect 356 407 358 409
rect 20 384 22 386
rect 25 384 27 386
rect 46 384 48 386
rect 56 384 58 386
rect 66 384 68 386
rect 76 384 78 386
rect 86 384 88 386
rect 96 384 98 386
rect 106 384 108 386
rect 149 384 151 386
rect 177 384 179 386
rect 182 384 184 386
rect 209 384 211 386
rect 252 384 254 386
rect 262 384 264 386
rect 272 384 274 386
rect 282 384 284 386
rect 292 384 294 386
rect 302 384 304 386
rect 312 384 314 386
rect 333 384 335 386
rect 338 384 340 386
rect 20 379 22 381
rect 25 379 27 381
rect 46 379 48 381
rect 56 379 58 381
rect 66 379 68 381
rect 76 379 78 381
rect 86 379 88 381
rect 96 379 98 381
rect 106 379 108 381
rect 149 379 151 381
rect 177 379 179 381
rect 182 379 184 381
rect 209 379 211 381
rect 252 379 254 381
rect 262 379 264 381
rect 272 379 274 381
rect 282 379 284 381
rect 292 379 294 381
rect 302 379 304 381
rect 312 379 314 381
rect 333 379 335 381
rect 338 379 340 381
rect 20 374 22 376
rect 25 374 27 376
rect 46 374 48 376
rect 56 374 58 376
rect 66 374 68 376
rect 76 374 78 376
rect 86 374 88 376
rect 96 374 98 376
rect 106 374 108 376
rect 149 374 151 376
rect 177 374 179 376
rect 182 374 184 376
rect 209 374 211 376
rect 252 374 254 376
rect 262 374 264 376
rect 272 374 274 376
rect 282 374 284 376
rect 292 374 294 376
rect 302 374 304 376
rect 312 374 314 376
rect 333 374 335 376
rect 338 374 340 376
rect 2 359 4 361
rect 7 359 9 361
rect 351 359 353 361
rect 356 359 358 361
rect 2 351 4 353
rect 7 351 9 353
rect 351 351 353 353
rect 356 351 358 353
rect 2 343 4 345
rect 7 343 9 345
rect 351 343 353 345
rect 356 343 358 345
rect 20 319 22 321
rect 25 319 27 321
rect 46 319 48 321
rect 56 319 58 321
rect 66 319 68 321
rect 76 319 78 321
rect 86 319 88 321
rect 96 319 98 321
rect 106 319 108 321
rect 149 319 151 321
rect 177 319 179 321
rect 182 319 184 321
rect 209 319 211 321
rect 252 319 254 321
rect 262 319 264 321
rect 272 319 274 321
rect 282 319 284 321
rect 292 319 294 321
rect 302 319 304 321
rect 312 319 314 321
rect 333 319 335 321
rect 338 319 340 321
rect 20 314 22 316
rect 25 314 27 316
rect 46 314 48 316
rect 56 314 58 316
rect 66 314 68 316
rect 76 314 78 316
rect 86 314 88 316
rect 96 314 98 316
rect 106 314 108 316
rect 149 314 151 316
rect 177 314 179 316
rect 182 314 184 316
rect 209 314 211 316
rect 252 314 254 316
rect 262 314 264 316
rect 272 314 274 316
rect 282 314 284 316
rect 292 314 294 316
rect 302 314 304 316
rect 312 314 314 316
rect 333 314 335 316
rect 338 314 340 316
rect 20 309 22 311
rect 25 309 27 311
rect 46 309 48 311
rect 56 309 58 311
rect 66 309 68 311
rect 76 309 78 311
rect 86 309 88 311
rect 96 309 98 311
rect 106 309 108 311
rect 149 309 151 311
rect 177 309 179 311
rect 182 309 184 311
rect 209 309 211 311
rect 252 309 254 311
rect 262 309 264 311
rect 272 309 274 311
rect 282 309 284 311
rect 292 309 294 311
rect 302 309 304 311
rect 312 309 314 311
rect 333 309 335 311
rect 338 309 340 311
rect 2 294 4 296
rect 7 294 9 296
rect 351 294 353 296
rect 356 294 358 296
rect 2 286 4 288
rect 7 286 9 288
rect 351 286 353 288
rect 356 286 358 288
rect 2 278 4 280
rect 7 278 9 280
rect 351 278 353 280
rect 356 278 358 280
rect 20 254 22 256
rect 25 254 27 256
rect 46 254 48 256
rect 56 254 58 256
rect 66 254 68 256
rect 76 254 78 256
rect 86 254 88 256
rect 96 254 98 256
rect 106 254 108 256
rect 149 254 151 256
rect 177 254 179 256
rect 182 254 184 256
rect 209 254 211 256
rect 252 254 254 256
rect 262 254 264 256
rect 272 254 274 256
rect 282 254 284 256
rect 292 254 294 256
rect 302 254 304 256
rect 312 254 314 256
rect 333 254 335 256
rect 338 254 340 256
rect 20 249 22 251
rect 25 249 27 251
rect 46 249 48 251
rect 56 249 58 251
rect 66 249 68 251
rect 76 249 78 251
rect 86 249 88 251
rect 96 249 98 251
rect 106 249 108 251
rect 149 249 151 251
rect 177 249 179 251
rect 182 249 184 251
rect 209 249 211 251
rect 252 249 254 251
rect 262 249 264 251
rect 272 249 274 251
rect 282 249 284 251
rect 292 249 294 251
rect 302 249 304 251
rect 312 249 314 251
rect 333 249 335 251
rect 338 249 340 251
rect 20 244 22 246
rect 25 244 27 246
rect 46 244 48 246
rect 56 244 58 246
rect 66 244 68 246
rect 76 244 78 246
rect 86 244 88 246
rect 96 244 98 246
rect 106 244 108 246
rect 149 244 151 246
rect 177 244 179 246
rect 182 244 184 246
rect 209 244 211 246
rect 252 244 254 246
rect 262 244 264 246
rect 272 244 274 246
rect 282 244 284 246
rect 292 244 294 246
rect 302 244 304 246
rect 312 244 314 246
rect 333 244 335 246
rect 338 244 340 246
rect 5 226 7 228
rect 13 226 15 228
rect 21 226 23 228
rect 45 226 47 228
rect 53 226 55 228
rect 61 226 63 228
rect 69 226 71 228
rect 77 226 79 228
rect 85 226 87 228
rect 93 226 95 228
rect 101 226 103 228
rect 109 226 111 228
rect 149 226 151 228
rect 181 226 183 228
rect 209 226 211 228
rect 249 226 251 228
rect 257 226 259 228
rect 265 226 267 228
rect 273 226 275 228
rect 281 226 283 228
rect 289 226 291 228
rect 297 226 299 228
rect 305 226 307 228
rect 313 226 315 228
rect 337 226 339 228
rect 345 226 347 228
rect 353 226 355 228
rect 5 221 7 223
rect 13 221 15 223
rect 21 221 23 223
rect 45 221 47 223
rect 53 221 55 223
rect 61 221 63 223
rect 69 221 71 223
rect 77 221 79 223
rect 85 221 87 223
rect 93 221 95 223
rect 101 221 103 223
rect 109 221 111 223
rect 149 221 151 223
rect 181 221 183 223
rect 209 221 211 223
rect 249 221 251 223
rect 257 221 259 223
rect 265 221 267 223
rect 273 221 275 223
rect 281 221 283 223
rect 289 221 291 223
rect 297 221 299 223
rect 305 221 307 223
rect 313 221 315 223
rect 337 221 339 223
rect 345 221 347 223
rect 353 221 355 223
rect 5 209 7 211
rect 13 209 15 211
rect 21 209 23 211
rect 45 209 47 211
rect 53 209 55 211
rect 61 209 63 211
rect 69 209 71 211
rect 77 209 79 211
rect 85 209 87 211
rect 93 209 95 211
rect 101 209 103 211
rect 109 209 111 211
rect 149 209 151 211
rect 181 209 183 211
rect 209 209 211 211
rect 249 209 251 211
rect 257 209 259 211
rect 265 209 267 211
rect 273 209 275 211
rect 281 209 283 211
rect 289 209 291 211
rect 297 209 299 211
rect 305 209 307 211
rect 313 209 315 211
rect 337 209 339 211
rect 345 209 347 211
rect 353 209 355 211
rect 5 204 7 206
rect 13 204 15 206
rect 21 204 23 206
rect 45 204 47 206
rect 53 204 55 206
rect 61 204 63 206
rect 69 204 71 206
rect 77 204 79 206
rect 85 204 87 206
rect 93 204 95 206
rect 101 204 103 206
rect 109 204 111 206
rect 149 204 151 206
rect 181 204 183 206
rect 209 204 211 206
rect 249 204 251 206
rect 257 204 259 206
rect 265 204 267 206
rect 273 204 275 206
rect 281 204 283 206
rect 289 204 291 206
rect 297 204 299 206
rect 305 204 307 206
rect 313 204 315 206
rect 337 204 339 206
rect 345 204 347 206
rect 353 204 355 206
rect 33 195 35 197
rect 38 195 40 197
rect 157 195 159 197
rect 162 195 164 197
rect 196 195 198 197
rect 201 195 203 197
rect 320 195 322 197
rect 325 195 327 197
rect 33 190 35 192
rect 38 190 40 192
rect 157 190 159 192
rect 162 190 164 192
rect 196 190 198 192
rect 201 190 203 192
rect 320 190 322 192
rect 325 190 327 192
rect 169 181 171 183
rect 174 181 176 183
rect 179 181 181 183
rect 184 181 186 183
rect 189 181 191 183
rect 320 181 322 183
rect 325 181 327 183
rect 169 176 171 178
rect 174 176 176 178
rect 179 176 181 178
rect 184 176 186 178
rect 189 176 191 178
rect 320 176 322 178
rect 325 176 327 178
rect 3 96 5 98
rect 45 96 47 98
rect 53 96 55 98
rect 61 96 63 98
rect 69 96 71 98
rect 77 96 79 98
rect 85 96 87 98
rect 93 96 95 98
rect 101 96 103 98
rect 109 96 111 98
rect 117 96 119 98
rect 125 96 127 98
rect 133 96 135 98
rect 141 96 143 98
rect 149 96 151 98
rect 157 96 159 98
rect 165 96 167 98
rect 193 96 195 98
rect 201 96 203 98
rect 209 96 211 98
rect 217 96 219 98
rect 225 96 227 98
rect 233 96 235 98
rect 241 96 243 98
rect 249 96 251 98
rect 257 96 259 98
rect 265 96 267 98
rect 273 96 275 98
rect 281 96 283 98
rect 289 96 291 98
rect 297 96 299 98
rect 305 96 307 98
rect 313 96 315 98
rect 355 96 357 98
rect 3 91 5 93
rect 45 91 47 93
rect 53 91 55 93
rect 61 91 63 93
rect 69 91 71 93
rect 77 91 79 93
rect 85 91 87 93
rect 93 91 95 93
rect 101 91 103 93
rect 109 91 111 93
rect 117 91 119 93
rect 125 91 127 93
rect 133 91 135 93
rect 141 91 143 93
rect 149 91 151 93
rect 157 91 159 93
rect 165 91 167 93
rect 193 91 195 93
rect 201 91 203 93
rect 209 91 211 93
rect 217 91 219 93
rect 225 91 227 93
rect 233 91 235 93
rect 241 91 243 93
rect 249 91 251 93
rect 257 91 259 93
rect 265 91 267 93
rect 273 91 275 93
rect 281 91 283 93
rect 289 91 291 93
rect 297 91 299 93
rect 305 91 307 93
rect 313 91 315 93
rect 355 91 357 93
rect 3 81 5 83
rect 127 81 129 83
rect 301 81 303 83
rect 355 81 357 83
rect 81 66 83 68
rect 105 52 107 54
rect 119 52 121 54
rect 239 52 241 54
rect 253 52 255 54
rect 112 45 114 47
rect 246 45 248 47
rect 277 38 279 40
rect 3 2 5 4
rect 72 2 74 4
rect 284 2 286 4
rect 348 2 350 4
<< metal3 >>
rect 51 1116 309 1120
rect 51 866 55 1116
rect 305 866 309 1116
rect 51 862 309 866
<< gv2 >>
rect 64 1105 66 1107
rect 74 1105 76 1107
rect 84 1105 86 1107
rect 94 1105 96 1107
rect 104 1105 106 1107
rect 114 1105 116 1107
rect 124 1105 126 1107
rect 134 1105 136 1107
rect 144 1105 146 1107
rect 154 1105 156 1107
rect 164 1105 166 1107
rect 174 1105 176 1107
rect 184 1105 186 1107
rect 194 1105 196 1107
rect 204 1105 206 1107
rect 214 1105 216 1107
rect 224 1105 226 1107
rect 234 1105 236 1107
rect 244 1105 246 1107
rect 254 1105 256 1107
rect 264 1105 266 1107
rect 274 1105 276 1107
rect 284 1105 286 1107
rect 294 1105 296 1107
rect 64 1095 66 1097
rect 74 1095 76 1097
rect 84 1095 86 1097
rect 94 1095 96 1097
rect 104 1095 106 1097
rect 114 1095 116 1097
rect 124 1095 126 1097
rect 134 1095 136 1097
rect 144 1095 146 1097
rect 154 1095 156 1097
rect 164 1095 166 1097
rect 174 1095 176 1097
rect 184 1095 186 1097
rect 194 1095 196 1097
rect 204 1095 206 1097
rect 214 1095 216 1097
rect 224 1095 226 1097
rect 234 1095 236 1097
rect 244 1095 246 1097
rect 254 1095 256 1097
rect 264 1095 266 1097
rect 274 1095 276 1097
rect 284 1095 286 1097
rect 294 1095 296 1097
rect 64 1085 66 1087
rect 74 1085 76 1087
rect 84 1085 86 1087
rect 94 1085 96 1087
rect 104 1085 106 1087
rect 114 1085 116 1087
rect 124 1085 126 1087
rect 134 1085 136 1087
rect 144 1085 146 1087
rect 154 1085 156 1087
rect 164 1085 166 1087
rect 174 1085 176 1087
rect 184 1085 186 1087
rect 194 1085 196 1087
rect 204 1085 206 1087
rect 214 1085 216 1087
rect 224 1085 226 1087
rect 234 1085 236 1087
rect 244 1085 246 1087
rect 254 1085 256 1087
rect 264 1085 266 1087
rect 274 1085 276 1087
rect 284 1085 286 1087
rect 294 1085 296 1087
rect 64 1075 66 1077
rect 74 1075 76 1077
rect 84 1075 86 1077
rect 94 1075 96 1077
rect 104 1075 106 1077
rect 114 1075 116 1077
rect 124 1075 126 1077
rect 134 1075 136 1077
rect 144 1075 146 1077
rect 154 1075 156 1077
rect 164 1075 166 1077
rect 174 1075 176 1077
rect 184 1075 186 1077
rect 194 1075 196 1077
rect 204 1075 206 1077
rect 214 1075 216 1077
rect 224 1075 226 1077
rect 234 1075 236 1077
rect 244 1075 246 1077
rect 254 1075 256 1077
rect 264 1075 266 1077
rect 274 1075 276 1077
rect 284 1075 286 1077
rect 294 1075 296 1077
rect 64 1065 66 1067
rect 74 1065 76 1067
rect 84 1065 86 1067
rect 94 1065 96 1067
rect 104 1065 106 1067
rect 114 1065 116 1067
rect 124 1065 126 1067
rect 134 1065 136 1067
rect 144 1065 146 1067
rect 154 1065 156 1067
rect 164 1065 166 1067
rect 174 1065 176 1067
rect 184 1065 186 1067
rect 194 1065 196 1067
rect 204 1065 206 1067
rect 214 1065 216 1067
rect 224 1065 226 1067
rect 234 1065 236 1067
rect 244 1065 246 1067
rect 254 1065 256 1067
rect 264 1065 266 1067
rect 274 1065 276 1067
rect 284 1065 286 1067
rect 294 1065 296 1067
rect 64 1055 66 1057
rect 74 1055 76 1057
rect 84 1055 86 1057
rect 94 1055 96 1057
rect 104 1055 106 1057
rect 114 1055 116 1057
rect 124 1055 126 1057
rect 134 1055 136 1057
rect 144 1055 146 1057
rect 154 1055 156 1057
rect 164 1055 166 1057
rect 174 1055 176 1057
rect 184 1055 186 1057
rect 194 1055 196 1057
rect 204 1055 206 1057
rect 214 1055 216 1057
rect 224 1055 226 1057
rect 234 1055 236 1057
rect 244 1055 246 1057
rect 254 1055 256 1057
rect 264 1055 266 1057
rect 274 1055 276 1057
rect 284 1055 286 1057
rect 294 1055 296 1057
rect 64 1045 66 1047
rect 74 1045 76 1047
rect 84 1045 86 1047
rect 94 1045 96 1047
rect 104 1045 106 1047
rect 114 1045 116 1047
rect 124 1045 126 1047
rect 134 1045 136 1047
rect 144 1045 146 1047
rect 154 1045 156 1047
rect 164 1045 166 1047
rect 174 1045 176 1047
rect 184 1045 186 1047
rect 194 1045 196 1047
rect 204 1045 206 1047
rect 214 1045 216 1047
rect 224 1045 226 1047
rect 234 1045 236 1047
rect 244 1045 246 1047
rect 254 1045 256 1047
rect 264 1045 266 1047
rect 274 1045 276 1047
rect 284 1045 286 1047
rect 294 1045 296 1047
rect 64 1035 66 1037
rect 74 1035 76 1037
rect 84 1035 86 1037
rect 94 1035 96 1037
rect 104 1035 106 1037
rect 114 1035 116 1037
rect 124 1035 126 1037
rect 134 1035 136 1037
rect 144 1035 146 1037
rect 154 1035 156 1037
rect 164 1035 166 1037
rect 174 1035 176 1037
rect 184 1035 186 1037
rect 194 1035 196 1037
rect 204 1035 206 1037
rect 214 1035 216 1037
rect 224 1035 226 1037
rect 234 1035 236 1037
rect 244 1035 246 1037
rect 254 1035 256 1037
rect 264 1035 266 1037
rect 274 1035 276 1037
rect 284 1035 286 1037
rect 294 1035 296 1037
rect 64 1025 66 1027
rect 74 1025 76 1027
rect 84 1025 86 1027
rect 94 1025 96 1027
rect 104 1025 106 1027
rect 114 1025 116 1027
rect 124 1025 126 1027
rect 134 1025 136 1027
rect 144 1025 146 1027
rect 154 1025 156 1027
rect 164 1025 166 1027
rect 174 1025 176 1027
rect 184 1025 186 1027
rect 194 1025 196 1027
rect 204 1025 206 1027
rect 214 1025 216 1027
rect 224 1025 226 1027
rect 234 1025 236 1027
rect 244 1025 246 1027
rect 254 1025 256 1027
rect 264 1025 266 1027
rect 274 1025 276 1027
rect 284 1025 286 1027
rect 294 1025 296 1027
rect 64 1015 66 1017
rect 74 1015 76 1017
rect 84 1015 86 1017
rect 94 1015 96 1017
rect 104 1015 106 1017
rect 114 1015 116 1017
rect 124 1015 126 1017
rect 134 1015 136 1017
rect 144 1015 146 1017
rect 154 1015 156 1017
rect 164 1015 166 1017
rect 174 1015 176 1017
rect 184 1015 186 1017
rect 194 1015 196 1017
rect 204 1015 206 1017
rect 214 1015 216 1017
rect 224 1015 226 1017
rect 234 1015 236 1017
rect 244 1015 246 1017
rect 254 1015 256 1017
rect 264 1015 266 1017
rect 274 1015 276 1017
rect 284 1015 286 1017
rect 294 1015 296 1017
rect 64 1005 66 1007
rect 74 1005 76 1007
rect 84 1005 86 1007
rect 94 1005 96 1007
rect 104 1005 106 1007
rect 114 1005 116 1007
rect 124 1005 126 1007
rect 134 1005 136 1007
rect 144 1005 146 1007
rect 154 1005 156 1007
rect 164 1005 166 1007
rect 174 1005 176 1007
rect 184 1005 186 1007
rect 194 1005 196 1007
rect 204 1005 206 1007
rect 214 1005 216 1007
rect 224 1005 226 1007
rect 234 1005 236 1007
rect 244 1005 246 1007
rect 254 1005 256 1007
rect 264 1005 266 1007
rect 274 1005 276 1007
rect 284 1005 286 1007
rect 294 1005 296 1007
rect 64 995 66 997
rect 74 995 76 997
rect 84 995 86 997
rect 94 995 96 997
rect 104 995 106 997
rect 114 995 116 997
rect 124 995 126 997
rect 134 995 136 997
rect 144 995 146 997
rect 154 995 156 997
rect 164 995 166 997
rect 174 995 176 997
rect 184 995 186 997
rect 194 995 196 997
rect 204 995 206 997
rect 214 995 216 997
rect 224 995 226 997
rect 234 995 236 997
rect 244 995 246 997
rect 254 995 256 997
rect 264 995 266 997
rect 274 995 276 997
rect 284 995 286 997
rect 294 995 296 997
rect 64 985 66 987
rect 74 985 76 987
rect 84 985 86 987
rect 94 985 96 987
rect 104 985 106 987
rect 114 985 116 987
rect 124 985 126 987
rect 134 985 136 987
rect 144 985 146 987
rect 154 985 156 987
rect 164 985 166 987
rect 174 985 176 987
rect 184 985 186 987
rect 194 985 196 987
rect 204 985 206 987
rect 214 985 216 987
rect 224 985 226 987
rect 234 985 236 987
rect 244 985 246 987
rect 254 985 256 987
rect 264 985 266 987
rect 274 985 276 987
rect 284 985 286 987
rect 294 985 296 987
rect 64 975 66 977
rect 74 975 76 977
rect 84 975 86 977
rect 94 975 96 977
rect 104 975 106 977
rect 114 975 116 977
rect 124 975 126 977
rect 134 975 136 977
rect 144 975 146 977
rect 154 975 156 977
rect 164 975 166 977
rect 174 975 176 977
rect 184 975 186 977
rect 194 975 196 977
rect 204 975 206 977
rect 214 975 216 977
rect 224 975 226 977
rect 234 975 236 977
rect 244 975 246 977
rect 254 975 256 977
rect 264 975 266 977
rect 274 975 276 977
rect 284 975 286 977
rect 294 975 296 977
rect 64 965 66 967
rect 74 965 76 967
rect 84 965 86 967
rect 94 965 96 967
rect 104 965 106 967
rect 114 965 116 967
rect 124 965 126 967
rect 134 965 136 967
rect 144 965 146 967
rect 154 965 156 967
rect 164 965 166 967
rect 174 965 176 967
rect 184 965 186 967
rect 194 965 196 967
rect 204 965 206 967
rect 214 965 216 967
rect 224 965 226 967
rect 234 965 236 967
rect 244 965 246 967
rect 254 965 256 967
rect 264 965 266 967
rect 274 965 276 967
rect 284 965 286 967
rect 294 965 296 967
rect 64 955 66 957
rect 74 955 76 957
rect 84 955 86 957
rect 94 955 96 957
rect 104 955 106 957
rect 114 955 116 957
rect 124 955 126 957
rect 134 955 136 957
rect 144 955 146 957
rect 154 955 156 957
rect 164 955 166 957
rect 174 955 176 957
rect 184 955 186 957
rect 194 955 196 957
rect 204 955 206 957
rect 214 955 216 957
rect 224 955 226 957
rect 234 955 236 957
rect 244 955 246 957
rect 254 955 256 957
rect 264 955 266 957
rect 274 955 276 957
rect 284 955 286 957
rect 294 955 296 957
rect 64 945 66 947
rect 74 945 76 947
rect 84 945 86 947
rect 94 945 96 947
rect 104 945 106 947
rect 114 945 116 947
rect 124 945 126 947
rect 134 945 136 947
rect 144 945 146 947
rect 154 945 156 947
rect 164 945 166 947
rect 174 945 176 947
rect 184 945 186 947
rect 194 945 196 947
rect 204 945 206 947
rect 214 945 216 947
rect 224 945 226 947
rect 234 945 236 947
rect 244 945 246 947
rect 254 945 256 947
rect 264 945 266 947
rect 274 945 276 947
rect 284 945 286 947
rect 294 945 296 947
rect 64 935 66 937
rect 74 935 76 937
rect 84 935 86 937
rect 94 935 96 937
rect 104 935 106 937
rect 114 935 116 937
rect 124 935 126 937
rect 134 935 136 937
rect 144 935 146 937
rect 154 935 156 937
rect 164 935 166 937
rect 174 935 176 937
rect 184 935 186 937
rect 194 935 196 937
rect 204 935 206 937
rect 214 935 216 937
rect 224 935 226 937
rect 234 935 236 937
rect 244 935 246 937
rect 254 935 256 937
rect 264 935 266 937
rect 274 935 276 937
rect 284 935 286 937
rect 294 935 296 937
rect 64 925 66 927
rect 74 925 76 927
rect 84 925 86 927
rect 94 925 96 927
rect 104 925 106 927
rect 114 925 116 927
rect 124 925 126 927
rect 134 925 136 927
rect 144 925 146 927
rect 154 925 156 927
rect 164 925 166 927
rect 174 925 176 927
rect 184 925 186 927
rect 194 925 196 927
rect 204 925 206 927
rect 214 925 216 927
rect 224 925 226 927
rect 234 925 236 927
rect 244 925 246 927
rect 254 925 256 927
rect 264 925 266 927
rect 274 925 276 927
rect 284 925 286 927
rect 294 925 296 927
rect 64 915 66 917
rect 74 915 76 917
rect 84 915 86 917
rect 94 915 96 917
rect 104 915 106 917
rect 114 915 116 917
rect 124 915 126 917
rect 134 915 136 917
rect 144 915 146 917
rect 154 915 156 917
rect 164 915 166 917
rect 174 915 176 917
rect 184 915 186 917
rect 194 915 196 917
rect 204 915 206 917
rect 214 915 216 917
rect 224 915 226 917
rect 234 915 236 917
rect 244 915 246 917
rect 254 915 256 917
rect 264 915 266 917
rect 274 915 276 917
rect 284 915 286 917
rect 294 915 296 917
rect 64 905 66 907
rect 74 905 76 907
rect 84 905 86 907
rect 94 905 96 907
rect 104 905 106 907
rect 114 905 116 907
rect 124 905 126 907
rect 134 905 136 907
rect 144 905 146 907
rect 154 905 156 907
rect 164 905 166 907
rect 174 905 176 907
rect 184 905 186 907
rect 194 905 196 907
rect 204 905 206 907
rect 214 905 216 907
rect 224 905 226 907
rect 234 905 236 907
rect 244 905 246 907
rect 254 905 256 907
rect 264 905 266 907
rect 274 905 276 907
rect 284 905 286 907
rect 294 905 296 907
rect 64 895 66 897
rect 74 895 76 897
rect 84 895 86 897
rect 94 895 96 897
rect 104 895 106 897
rect 114 895 116 897
rect 124 895 126 897
rect 134 895 136 897
rect 144 895 146 897
rect 154 895 156 897
rect 164 895 166 897
rect 174 895 176 897
rect 184 895 186 897
rect 194 895 196 897
rect 204 895 206 897
rect 214 895 216 897
rect 224 895 226 897
rect 234 895 236 897
rect 244 895 246 897
rect 254 895 256 897
rect 264 895 266 897
rect 274 895 276 897
rect 284 895 286 897
rect 294 895 296 897
rect 64 885 66 887
rect 74 885 76 887
rect 84 885 86 887
rect 94 885 96 887
rect 104 885 106 887
rect 114 885 116 887
rect 124 885 126 887
rect 134 885 136 887
rect 144 885 146 887
rect 154 885 156 887
rect 164 885 166 887
rect 174 885 176 887
rect 184 885 186 887
rect 194 885 196 887
rect 204 885 206 887
rect 214 885 216 887
rect 224 885 226 887
rect 234 885 236 887
rect 244 885 246 887
rect 254 885 256 887
rect 264 885 266 887
rect 274 885 276 887
rect 284 885 286 887
rect 294 885 296 887
rect 64 875 66 877
rect 74 875 76 877
rect 84 875 86 877
rect 94 875 96 877
rect 104 875 106 877
rect 114 875 116 877
rect 124 875 126 877
rect 134 875 136 877
rect 144 875 146 877
rect 154 875 156 877
rect 164 875 166 877
rect 174 875 176 877
rect 184 875 186 877
rect 194 875 196 877
rect 204 875 206 877
rect 214 875 216 877
rect 224 875 226 877
rect 234 875 236 877
rect 244 875 246 877
rect 254 875 256 877
rect 264 875 266 877
rect 274 875 276 877
rect 284 875 286 877
rect 294 875 296 877
<< pad >>
rect 55 866 305 1116
<< pseudo_rnwell >>
rect 80 136 81 160
rect 279 136 280 160
<< rnwell >>
rect 81 136 279 160
use inv_e  inv_e_0
timestamp 1592016665
transform 1 0 23 0 -1 82
box -4 0 44 81
use nor2_b  nor2_b_0
timestamp 1591571333
transform -1 0 125 0 -1 82
box -3 0 28 81
use nand2_c  nand2_c_0
timestamp 1592098687
transform 1 0 62 0 -1 82
box -4 0 44 81
use subc_2  subc_2_0
timestamp 1592016765
transform 1 0 -3 0 -1 82
box -1 0 15 81
use nand2_b  nand2_b_1
timestamp 1592278238
transform 1 0 235 0 -1 82
box -4 0 28 81
use nor2_c  nor2_c_0
timestamp 1592096983
transform 1 0 258 0 -1 82
box -3 0 43 81
use inv_e  inv_e_1
timestamp 1592016665
transform 1 0 297 0 -1 82
box -4 0 44 81
use subc_2  subc_2_1
timestamp 1592016765
transform 1 0 349 0 -1 82
box -1 0 15 81
<< labels >>
rlabel metal1 s 145 800 145 800 2 pad
port 1 ne
rlabel nwell s -2 220 -2 220 2 vdd
rlabel metal2 s 340 208 340 208 2 vss
rlabel metal2 s 340 532 340 532 2 vss
port 8 ne
rlabel metal2 s 340 488 340 488 2 vss
rlabel metal2 s 336 447 336 447 2 vss
rlabel metal2 s 340 470 340 470 2 vdd
rlabel metal2 s 340 515 340 515 2 vdd
rlabel metal2 s 336 555 336 555 2 vdd
port 7 ne
rlabel metal2 48 191 48 191 2 pd
rlabel rnwell s 168 146 168 146 2 r0_body
rlabel metal2 s -13 15 -13 15 2 vss
rlabel metal2 s 166 75 166 75 4 ntri
port 6 ne
rlabel metal2 s 207 68 207 68 4 tri
port 5 ne
rlabel metal2 s 207 61 207 61 4 adly
rlabel metal2 s 208 54 208 54 4 a
rlabel metal1 s 79 4 79 4 4 vdd
rlabel metal1 s 75 83 75 83 4 vss
rlabel metal2 57 68 57 68 4 npd
rlabel metal2 109 46 109 46 4 apd
rlabel metal2 s 312 94 312 94 2 vss
rlabel metal2 256 47 256 47 4 anpu
rlabel metal2 289 40 289 40 4 pu
rlabel metal1 s 178 93 178 93 2 xpad
port 2 ne
rlabel metal2 323 179 323 179 2 npu
<< end >>
