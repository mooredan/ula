magic
tech amic5n
timestamp 1608317706
<< poly2 >>
rect 930 1200 1080 1350
rect 4020 1200 4200 1350
