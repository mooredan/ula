`celldefine
module xor2_a (z, a, b);
  output z;
  input  a;
  input  b;

  xor G1 (z, a, b);
endmodule
`endcelldefine
