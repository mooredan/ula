magic
tech amic5n
timestamp 1624413463
<< nwell >>
rect -130 550 1780 1495
<< ntransistor >>
rect 225 95 285 400
rect 465 95 525 400
rect 1045 125 1105 400
rect 1235 125 1295 400
rect 1425 125 1485 400
<< ptransistor >>
rect 225 705 285 1345
rect 465 705 525 1345
rect 1045 705 1105 1290
rect 1235 705 1295 1290
rect 1425 705 1485 1290
<< nselect >>
rect 760 765 925 1290
rect -10 350 1660 430
rect -10 125 760 350
rect 925 125 1660 350
rect -10 0 1660 125
<< pselect >>
rect -10 1290 1660 1440
rect -10 765 760 1290
rect 925 765 1660 1290
rect -10 670 1660 765
rect 760 125 925 350
<< ndiffusion >>
rect 105 370 225 400
rect 105 320 135 370
rect 185 320 225 370
rect 105 175 225 320
rect 105 125 135 175
rect 185 125 225 175
rect 105 95 225 125
rect 285 95 465 400
rect 525 345 645 400
rect 925 370 1045 400
rect 525 295 565 345
rect 615 295 645 345
rect 525 185 645 295
rect 525 135 565 185
rect 615 135 645 185
rect 525 95 645 135
rect 925 320 955 370
rect 1005 320 1045 370
rect 925 205 1045 320
rect 925 155 955 205
rect 1005 155 1045 205
rect 925 125 1045 155
rect 1105 370 1235 400
rect 1105 320 1145 370
rect 1195 320 1235 370
rect 1105 205 1235 320
rect 1105 155 1145 205
rect 1195 155 1235 205
rect 1105 125 1235 155
rect 1295 345 1425 400
rect 1295 295 1335 345
rect 1385 295 1425 345
rect 1295 205 1425 295
rect 1295 155 1335 205
rect 1385 155 1425 205
rect 1295 125 1425 155
rect 1485 370 1605 400
rect 1485 320 1525 370
rect 1575 320 1605 370
rect 1485 205 1605 320
rect 1485 155 1525 205
rect 1575 155 1605 205
rect 1485 125 1605 155
<< pdiffusion >>
rect 105 1315 225 1345
rect 105 1265 135 1315
rect 185 1265 225 1315
rect 105 1215 225 1265
rect 105 1165 135 1215
rect 185 1165 225 1215
rect 105 1115 225 1165
rect 105 1065 135 1115
rect 185 1065 225 1115
rect 105 1015 225 1065
rect 105 965 135 1015
rect 185 965 225 1015
rect 105 915 225 965
rect 105 865 135 915
rect 185 865 225 915
rect 105 705 225 865
rect 285 1315 465 1345
rect 285 1265 350 1315
rect 400 1265 465 1315
rect 285 1185 465 1265
rect 285 1135 350 1185
rect 400 1135 465 1185
rect 285 1085 465 1135
rect 285 1035 350 1085
rect 400 1035 465 1085
rect 285 985 465 1035
rect 285 935 350 985
rect 400 935 465 985
rect 285 885 465 935
rect 285 835 350 885
rect 400 835 465 885
rect 285 785 465 835
rect 285 735 350 785
rect 400 735 465 785
rect 285 705 465 735
rect 525 1315 645 1345
rect 525 1265 565 1315
rect 615 1265 645 1315
rect 525 1215 645 1265
rect 525 1165 565 1215
rect 615 1165 645 1215
rect 525 1115 645 1165
rect 525 1065 565 1115
rect 615 1065 645 1115
rect 525 1015 645 1065
rect 525 965 565 1015
rect 615 965 645 1015
rect 525 915 645 965
rect 525 865 565 915
rect 615 865 645 915
rect 525 815 645 865
rect 525 765 565 815
rect 615 765 645 815
rect 925 1260 1045 1290
rect 925 1210 955 1260
rect 1005 1210 1045 1260
rect 925 1115 1045 1210
rect 925 1065 955 1115
rect 1005 1065 1045 1115
rect 925 1015 1045 1065
rect 925 965 955 1015
rect 1005 965 1045 1015
rect 925 915 1045 965
rect 925 865 955 915
rect 1005 865 1045 915
rect 925 815 1045 865
rect 925 765 955 815
rect 1005 765 1045 815
rect 525 705 645 765
rect 925 705 1045 765
rect 1105 1260 1235 1290
rect 1105 1210 1145 1260
rect 1195 1210 1235 1260
rect 1105 1080 1235 1210
rect 1105 1030 1145 1080
rect 1195 1030 1235 1080
rect 1105 980 1235 1030
rect 1105 930 1145 980
rect 1195 930 1235 980
rect 1105 825 1235 930
rect 1105 775 1145 825
rect 1195 775 1235 825
rect 1105 705 1235 775
rect 1295 1260 1425 1290
rect 1295 1210 1335 1260
rect 1385 1210 1425 1260
rect 1295 1115 1425 1210
rect 1295 1065 1335 1115
rect 1385 1065 1425 1115
rect 1295 975 1425 1065
rect 1295 925 1335 975
rect 1385 925 1425 975
rect 1295 705 1425 925
rect 1485 1260 1605 1290
rect 1485 1210 1525 1260
rect 1575 1210 1605 1260
rect 1485 1085 1605 1210
rect 1485 1035 1525 1085
rect 1575 1035 1605 1085
rect 1485 985 1605 1035
rect 1485 935 1525 985
rect 1575 935 1605 985
rect 1485 885 1605 935
rect 1485 835 1525 885
rect 1575 835 1605 885
rect 1485 785 1605 835
rect 1485 735 1525 785
rect 1575 735 1605 785
rect 1485 705 1605 735
<< psubstratepdiff >>
rect 810 320 925 350
rect 810 270 840 320
rect 890 270 925 320
rect 810 205 925 270
rect 810 155 840 205
rect 890 155 925 205
rect 810 125 925 155
<< nsubstratendiff >>
rect 810 1260 925 1290
rect 810 1210 845 1260
rect 895 1210 925 1260
rect 810 1160 925 1210
rect 810 1110 840 1160
rect 890 1110 925 1160
rect 810 1060 925 1110
rect 810 1010 840 1060
rect 890 1010 925 1060
rect 810 960 925 1010
rect 810 910 840 960
rect 890 910 925 960
rect 810 855 925 910
rect 810 805 840 855
rect 890 805 925 855
rect 810 765 925 805
<< nsubstratencontact >>
rect 845 1210 895 1260
rect 840 1110 890 1160
rect 840 1010 890 1060
rect 840 910 890 960
rect 840 805 890 855
<< psubstratepcontact >>
rect 840 270 890 320
rect 840 155 890 205
<< ndcontact >>
rect 135 320 185 370
rect 135 125 185 175
rect 565 295 615 345
rect 565 135 615 185
rect 955 320 1005 370
rect 955 155 1005 205
rect 1145 320 1195 370
rect 1145 155 1195 205
rect 1335 295 1385 345
rect 1335 155 1385 205
rect 1525 320 1575 370
rect 1525 155 1575 205
<< pdcontact >>
rect 135 1265 185 1315
rect 135 1165 185 1215
rect 135 1065 185 1115
rect 135 965 185 1015
rect 135 865 185 915
rect 350 1265 400 1315
rect 350 1135 400 1185
rect 350 1035 400 1085
rect 350 935 400 985
rect 350 835 400 885
rect 350 735 400 785
rect 565 1265 615 1315
rect 565 1165 615 1215
rect 565 1065 615 1115
rect 565 965 615 1015
rect 565 865 615 915
rect 565 765 615 815
rect 955 1210 1005 1260
rect 955 1065 1005 1115
rect 955 965 1005 1015
rect 955 865 1005 915
rect 955 765 1005 815
rect 1145 1210 1195 1260
rect 1145 1030 1195 1080
rect 1145 930 1195 980
rect 1145 775 1195 825
rect 1335 1210 1385 1260
rect 1335 1065 1385 1115
rect 1335 925 1385 975
rect 1525 1210 1575 1260
rect 1525 1035 1575 1085
rect 1525 935 1575 985
rect 1525 835 1575 885
rect 1525 735 1575 785
<< polysilicon >>
rect 225 1345 285 1410
rect 465 1345 525 1410
rect 1045 1290 1105 1355
rect 1235 1290 1295 1355
rect 1425 1290 1485 1355
rect 225 685 285 705
rect 115 665 285 685
rect 115 615 135 665
rect 185 615 285 665
rect 115 595 285 615
rect 225 400 285 595
rect 465 525 525 705
rect 1045 685 1105 705
rect 1235 685 1295 705
rect 1425 685 1485 705
rect 935 665 1485 685
rect 935 615 955 665
rect 1005 615 1055 665
rect 1105 615 1155 665
rect 1205 615 1255 665
rect 1305 615 1355 665
rect 1405 615 1485 665
rect 935 595 1485 615
rect 465 505 635 525
rect 465 455 565 505
rect 615 455 635 505
rect 465 435 635 455
rect 465 400 525 435
rect 1045 400 1105 595
rect 1235 400 1295 595
rect 1425 400 1485 595
rect 225 30 285 95
rect 465 30 525 95
rect 1045 60 1105 125
rect 1235 60 1295 125
rect 1425 60 1485 125
<< polycontact >>
rect 135 615 185 665
rect 955 615 1005 665
rect 1055 615 1105 665
rect 1155 615 1205 665
rect 1255 615 1305 665
rect 1355 615 1405 665
rect 565 455 615 505
<< metal1 >>
rect 0 1395 1650 1485
rect 115 1315 205 1395
rect 115 1265 135 1315
rect 185 1265 205 1315
rect 115 1215 205 1265
rect 115 1165 135 1215
rect 185 1165 205 1215
rect 115 1115 205 1165
rect 115 1065 135 1115
rect 185 1065 205 1115
rect 115 1015 205 1065
rect 115 965 135 1015
rect 185 965 205 1015
rect 115 915 205 965
rect 115 865 135 915
rect 185 865 205 915
rect 115 760 205 865
rect 330 1315 420 1335
rect 330 1265 350 1315
rect 400 1265 420 1315
rect 330 1185 420 1265
rect 330 1135 350 1185
rect 400 1135 420 1185
rect 330 1085 420 1135
rect 330 1035 350 1085
rect 400 1035 420 1085
rect 330 985 420 1035
rect 330 935 350 985
rect 400 935 420 985
rect 330 885 420 935
rect 330 835 350 885
rect 400 835 420 885
rect 330 785 420 835
rect 330 735 350 785
rect 400 735 420 785
rect 545 1315 635 1395
rect 545 1265 565 1315
rect 615 1265 635 1315
rect 545 1215 635 1265
rect 545 1165 565 1215
rect 615 1165 635 1215
rect 545 1115 635 1165
rect 545 1065 565 1115
rect 615 1065 635 1115
rect 545 1015 635 1065
rect 545 965 565 1015
rect 615 965 635 1015
rect 545 915 635 965
rect 545 865 565 915
rect 615 865 635 915
rect 545 815 635 865
rect 545 765 565 815
rect 615 765 635 815
rect 545 745 635 765
rect 820 1260 1025 1395
rect 820 1210 845 1260
rect 895 1210 955 1260
rect 1005 1210 1025 1260
rect 820 1160 1025 1210
rect 820 1110 840 1160
rect 890 1115 1025 1160
rect 890 1110 955 1115
rect 820 1065 955 1110
rect 1005 1065 1025 1115
rect 820 1060 1025 1065
rect 820 1010 840 1060
rect 890 1015 1025 1060
rect 890 1010 955 1015
rect 820 965 955 1010
rect 1005 965 1025 1015
rect 820 960 1025 965
rect 820 910 840 960
rect 890 915 1025 960
rect 890 910 955 915
rect 820 865 955 910
rect 1005 865 1025 915
rect 820 855 1025 865
rect 820 805 840 855
rect 890 815 1025 855
rect 890 805 955 815
rect 820 765 955 805
rect 1005 765 1025 815
rect 820 760 1025 765
rect 930 745 1025 760
rect 1125 1260 1215 1280
rect 1125 1210 1145 1260
rect 1195 1210 1215 1260
rect 1125 1080 1215 1210
rect 1125 1030 1145 1080
rect 1195 1030 1215 1080
rect 1125 980 1215 1030
rect 1125 930 1145 980
rect 1195 930 1215 980
rect 1125 845 1215 930
rect 1315 1260 1405 1395
rect 1315 1210 1335 1260
rect 1385 1210 1405 1260
rect 1315 1115 1405 1210
rect 1315 1065 1335 1115
rect 1385 1065 1405 1115
rect 1315 975 1405 1065
rect 1315 925 1335 975
rect 1385 925 1405 975
rect 1315 905 1405 925
rect 1505 1260 1595 1280
rect 1505 1210 1525 1260
rect 1575 1210 1595 1260
rect 1505 1085 1595 1210
rect 1505 1035 1525 1085
rect 1575 1035 1595 1085
rect 1505 985 1595 1035
rect 1505 935 1525 985
rect 1575 935 1595 985
rect 1505 885 1595 935
rect 1505 845 1525 885
rect 1125 835 1525 845
rect 1575 835 1595 885
rect 1125 825 1595 835
rect 1125 775 1145 825
rect 1195 785 1595 825
rect 1195 775 1525 785
rect 1125 755 1525 775
rect 330 685 420 735
rect 1505 735 1525 755
rect 1575 735 1595 785
rect 115 665 205 685
rect 115 615 135 665
rect 185 615 205 665
rect 115 595 205 615
rect 330 665 1425 685
rect 330 615 955 665
rect 1005 615 1055 665
rect 1105 615 1155 665
rect 1205 615 1255 665
rect 1305 615 1355 665
rect 1405 615 1425 665
rect 330 595 1425 615
rect 115 370 205 390
rect 115 320 135 370
rect 185 320 205 370
rect 115 175 205 320
rect 330 365 420 595
rect 1505 525 1595 735
rect 545 505 720 525
rect 545 455 565 505
rect 615 455 720 505
rect 545 435 720 455
rect 1125 435 1595 525
rect 935 370 1025 390
rect 330 345 635 365
rect 330 295 565 345
rect 615 295 635 345
rect 935 340 955 370
rect 330 275 635 295
rect 115 125 135 175
rect 185 125 205 175
rect 115 45 205 125
rect 545 185 635 275
rect 545 135 565 185
rect 615 135 635 185
rect 545 105 635 135
rect 820 320 955 340
rect 1005 320 1025 370
rect 820 270 840 320
rect 890 270 1025 320
rect 820 205 1025 270
rect 820 155 840 205
rect 890 155 955 205
rect 1005 155 1025 205
rect 820 45 1025 155
rect 1125 370 1215 435
rect 1125 320 1145 370
rect 1195 320 1215 370
rect 1505 370 1595 435
rect 1125 205 1215 320
rect 1125 155 1145 205
rect 1195 155 1215 205
rect 1125 135 1215 155
rect 1315 345 1405 365
rect 1315 295 1335 345
rect 1385 295 1405 345
rect 1315 205 1405 295
rect 1315 155 1335 205
rect 1385 155 1405 205
rect 1315 45 1405 155
rect 1505 320 1525 370
rect 1575 320 1595 370
rect 1505 205 1595 320
rect 1505 155 1525 205
rect 1575 155 1595 205
rect 1505 135 1595 155
rect 0 -45 1650 45
<< labels >>
flabel metal1 s 616 445 616 445 2 FreeSans 400 0 0 0 b
port 2 ne
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel nwell 5 585 5 585 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 1155 470 1155 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 135 605 135 605 2 FreeSans 400 0 0 0 a
port 1 ne
<< properties >>
string FIXED_BBOX 0 0 1650 1440
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
