magic
tech scmos
timestamp 1591463877
<< error_p >>
rect 0 16 2 17
rect 0 15 1 16
rect 0 7 2 9
rect 0 4 2 6
<< nwell >>
rect -9 -5 26 26
<< ptransistor >>
rect 5 2 7 20
<< pdiffusion >>
rect -2 2 5 20
rect 7 2 14 20
<< polysilicon >>
rect 5 20 7 37
rect 5 -11 7 2
<< genericcontact >>
rect 0 14 2 16
rect 0 4 2 6
<< metal1 >>
rect -1 12 3 18
rect -7 1 3 12
rect -1 -10 3 1
<< metal2 >>
rect -19 0 5 20
<< gv1 >>
rect 0 15 2 17
rect 0 7 2 9
rect -2 4 0 6
<< end >>
