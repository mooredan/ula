magic
tech scmos
timestamp 1570494029
<< error_p >>
rect 4 8 10 10
rect 4 6 6 8
rect 8 6 10 8
rect 4 4 10 6
rect -1 2 3 3
rect -1 0 0 2
rect 2 0 3 2
rect -1 -1 3 0
<< gv1 >>
rect 0 0 2 2
<< gv2 >>
rect 6 6 8 8
<< properties >>
string path 27.000 27.000 36.000 27.000 36.000 36.000 27.000 36.000 27.000 27.000 
<< end >>
