magic
tech amic5n
timestamp 1624309315
<< nwell >>
rect -130 550 880 1495
<< ntransistor >>
rect 160 125 220 400
rect 350 125 410 400
rect 540 125 600 400
<< ptransistor >>
rect 160 705 220 1290
rect 350 705 410 1290
rect 540 705 600 1290
<< nselect >>
rect -10 0 760 430
<< pselect >>
rect -10 670 760 1440
<< ndiffusion >>
rect 40 370 160 400
rect 40 320 70 370
rect 120 320 160 370
rect 40 205 160 320
rect 40 155 70 205
rect 120 155 160 205
rect 40 125 160 155
rect 220 370 350 400
rect 220 320 260 370
rect 310 320 350 370
rect 220 205 350 320
rect 220 155 260 205
rect 310 155 350 205
rect 220 125 350 155
rect 410 345 540 400
rect 410 295 450 345
rect 500 295 540 345
rect 410 205 540 295
rect 410 155 450 205
rect 500 155 540 205
rect 410 125 540 155
rect 600 370 720 400
rect 600 320 640 370
rect 690 320 720 370
rect 600 205 720 320
rect 600 155 640 205
rect 690 155 720 205
rect 600 125 720 155
<< pdiffusion >>
rect 40 1260 160 1290
rect 40 1210 70 1260
rect 120 1210 160 1260
rect 40 1115 160 1210
rect 40 1065 70 1115
rect 120 1065 160 1115
rect 40 1015 160 1065
rect 40 965 70 1015
rect 120 965 160 1015
rect 40 915 160 965
rect 40 865 70 915
rect 120 865 160 915
rect 40 815 160 865
rect 40 765 70 815
rect 120 765 160 815
rect 40 705 160 765
rect 220 1260 350 1290
rect 220 1210 260 1260
rect 310 1210 350 1260
rect 220 1080 350 1210
rect 220 1030 260 1080
rect 310 1030 350 1080
rect 220 980 350 1030
rect 220 930 260 980
rect 310 930 350 980
rect 220 825 350 930
rect 220 775 260 825
rect 310 775 350 825
rect 220 705 350 775
rect 410 1260 540 1290
rect 410 1210 450 1260
rect 500 1210 540 1260
rect 410 1115 540 1210
rect 410 1065 450 1115
rect 500 1065 540 1115
rect 410 975 540 1065
rect 410 925 450 975
rect 500 925 540 975
rect 410 705 540 925
rect 600 1260 720 1290
rect 600 1210 640 1260
rect 690 1210 720 1260
rect 600 1085 720 1210
rect 600 1035 640 1085
rect 690 1035 720 1085
rect 600 985 720 1035
rect 600 935 640 985
rect 690 935 720 985
rect 600 885 720 935
rect 600 835 640 885
rect 690 835 720 885
rect 600 785 720 835
rect 600 735 640 785
rect 690 735 720 785
rect 600 705 720 735
<< ndcontact >>
rect 70 320 120 370
rect 70 155 120 205
rect 260 320 310 370
rect 260 155 310 205
rect 450 295 500 345
rect 450 155 500 205
rect 640 320 690 370
rect 640 155 690 205
<< pdcontact >>
rect 70 1210 120 1260
rect 70 1065 120 1115
rect 70 965 120 1015
rect 70 865 120 915
rect 70 765 120 815
rect 260 1210 310 1260
rect 260 1030 310 1080
rect 260 930 310 980
rect 260 775 310 825
rect 450 1210 500 1260
rect 450 1065 500 1115
rect 450 925 500 975
rect 640 1210 690 1260
rect 640 1035 690 1085
rect 640 935 690 985
rect 640 835 690 885
rect 640 735 690 785
<< polysilicon >>
rect 160 1290 220 1355
rect 350 1290 410 1355
rect 540 1290 600 1355
rect 160 685 220 705
rect 350 685 410 705
rect 540 685 600 705
rect 50 665 600 685
rect 50 615 70 665
rect 120 615 170 665
rect 220 615 270 665
rect 320 615 370 665
rect 420 615 470 665
rect 520 615 600 665
rect 50 595 600 615
rect 160 400 220 595
rect 350 400 410 595
rect 540 400 600 595
rect 160 60 220 125
rect 350 60 410 125
rect 540 60 600 125
<< polycontact >>
rect 70 615 120 665
rect 170 615 220 665
rect 270 615 320 665
rect 370 615 420 665
rect 470 615 520 665
<< metal1 >>
rect 0 1395 750 1485
rect 50 1260 140 1395
rect 50 1210 70 1260
rect 120 1210 140 1260
rect 50 1115 140 1210
rect 50 1065 70 1115
rect 120 1065 140 1115
rect 50 1015 140 1065
rect 50 965 70 1015
rect 120 965 140 1015
rect 50 915 140 965
rect 50 865 70 915
rect 120 865 140 915
rect 50 815 140 865
rect 50 765 70 815
rect 120 765 140 815
rect 50 745 140 765
rect 240 1260 330 1280
rect 240 1210 260 1260
rect 310 1210 330 1260
rect 240 1080 330 1210
rect 240 1030 260 1080
rect 310 1030 330 1080
rect 240 980 330 1030
rect 240 930 260 980
rect 310 930 330 980
rect 240 845 330 930
rect 430 1260 520 1395
rect 430 1210 450 1260
rect 500 1210 520 1260
rect 430 1115 520 1210
rect 430 1065 450 1115
rect 500 1065 520 1115
rect 430 975 520 1065
rect 430 925 450 975
rect 500 925 520 975
rect 430 905 520 925
rect 620 1260 710 1280
rect 620 1210 640 1260
rect 690 1210 710 1260
rect 620 1085 710 1210
rect 620 1035 640 1085
rect 690 1035 710 1085
rect 620 985 710 1035
rect 620 935 640 985
rect 690 935 710 985
rect 620 885 710 935
rect 620 845 640 885
rect 240 835 640 845
rect 690 835 710 885
rect 240 825 710 835
rect 240 775 260 825
rect 310 785 710 825
rect 310 775 640 785
rect 240 755 640 775
rect 620 735 640 755
rect 690 735 710 785
rect 50 665 540 685
rect 50 615 70 665
rect 120 615 170 665
rect 220 615 270 665
rect 320 615 370 665
rect 420 615 470 665
rect 520 615 540 665
rect 50 595 540 615
rect 620 525 710 735
rect 240 435 710 525
rect 50 370 140 390
rect 50 320 70 370
rect 120 320 140 370
rect 50 205 140 320
rect 50 155 70 205
rect 120 155 140 205
rect 50 45 140 155
rect 240 370 330 435
rect 240 320 260 370
rect 310 320 330 370
rect 620 370 710 435
rect 240 205 330 320
rect 240 155 260 205
rect 310 155 330 205
rect 240 135 330 155
rect 430 345 520 365
rect 430 295 450 345
rect 500 295 520 345
rect 430 205 520 295
rect 430 155 450 205
rect 500 155 520 205
rect 430 45 520 155
rect 620 320 640 370
rect 690 320 710 370
rect 620 205 710 320
rect 620 155 640 205
rect 690 155 710 205
rect 620 135 710 155
rect 0 -45 750 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 3 ne
flabel metal1 s 20 1430 20 1430 2 FreeSans 400 0 0 0 vdd
port 2 ne
flabel metal1 s 270 470 270 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 70 605 70 605 2 FreeSans 400 0 0 0 a
port 1 ne
flabel nwell 35 555 35 555 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
<< end >>
