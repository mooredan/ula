magic
tech scmos
magscale 1 2
timestamp 1589157096
<< nwell >>
rect 30 1208 572 1304
rect 28 950 572 1208
rect 28 850 570 950
rect 284 848 570 850
rect -12 507 606 677
rect -6 498 606 507
rect -6 22 22 498
rect 572 22 606 498
rect -6 -6 606 22
<< ntransistor >>
rect 76 432 276 438
rect 76 342 276 348
rect 76 300 276 306
rect 76 212 276 218
rect 76 170 276 176
rect 76 82 276 88
rect 324 432 524 438
rect 324 342 524 348
rect 324 300 524 306
rect 324 212 524 218
rect 324 170 524 176
rect 324 82 524 88
<< ptransistor >>
rect 76 1248 276 1254
rect 76 1160 276 1166
rect 76 1118 276 1124
rect 76 1032 276 1038
rect 76 990 276 996
rect 76 902 276 908
rect 324 1248 524 1254
rect 324 1160 524 1166
rect 324 1118 524 1124
rect 324 1032 524 1038
rect 324 990 524 996
rect 324 902 524 908
<< ndiffusion >>
rect 76 438 276 456
rect 76 348 276 432
rect 76 306 276 342
rect 76 218 276 300
rect 76 176 276 212
rect 76 88 276 170
rect 76 64 276 82
rect 324 438 524 456
rect 324 348 524 432
rect 324 306 524 342
rect 324 218 524 300
rect 324 176 524 212
rect 324 88 524 170
rect 324 64 524 82
<< pdiffusion >>
rect 72 1260 280 1272
rect 76 1258 280 1260
rect 320 1260 528 1272
rect 320 1258 524 1260
rect 76 1254 276 1258
rect 76 1166 276 1248
rect 76 1124 276 1160
rect 76 1038 276 1118
rect 76 996 276 1032
rect 76 908 276 990
rect 76 884 276 902
rect 324 1254 524 1258
rect 324 1166 524 1248
rect 324 1124 524 1160
rect 324 1038 524 1118
rect 324 996 524 1032
rect 324 908 524 990
rect 324 884 524 902
<< psubstratepdiff >>
rect 0 1314 600 1340
rect 0 840 22 1314
rect 578 840 600 1314
rect 0 820 600 840
rect 0 696 12 820
rect 588 696 600 820
rect 0 684 600 696
rect 28 460 562 492
rect 28 60 60 460
rect 76 456 276 460
rect 76 60 276 64
rect 286 60 314 460
rect 324 456 524 460
rect 324 60 524 64
rect 540 60 562 460
rect 28 28 562 60
<< nsubstratendiff >>
rect 38 1272 562 1296
rect 38 1260 72 1272
rect 38 880 60 1260
rect 280 1258 320 1272
rect 528 1260 562 1272
rect 76 880 276 884
rect 284 880 316 1258
rect 324 880 524 884
rect 540 880 562 1260
rect 38 860 562 880
rect 0 652 600 664
rect 0 522 12 652
rect 588 530 600 652
rect 72 522 86 530
rect 112 522 600 530
rect 0 504 600 522
rect 0 16 16 504
rect 578 16 600 504
rect 0 0 600 16
<< polysilicon >>
rect 62 1248 76 1254
rect 276 1248 282 1254
rect 62 1166 74 1248
rect 278 1166 282 1248
rect 62 1160 76 1166
rect 276 1160 282 1166
rect 62 1124 74 1160
rect 278 1124 282 1160
rect 62 1118 76 1124
rect 276 1118 282 1124
rect 62 1038 74 1118
rect 278 1038 282 1118
rect 62 1032 76 1038
rect 276 1032 282 1038
rect 62 996 74 1032
rect 278 996 282 1032
rect 62 990 76 996
rect 276 990 282 996
rect 62 908 74 990
rect 278 908 282 990
rect 62 902 76 908
rect 276 902 282 908
rect 318 1248 324 1254
rect 524 1248 538 1254
rect 318 1166 322 1248
rect 526 1166 538 1248
rect 318 1160 324 1166
rect 524 1160 538 1166
rect 318 1124 322 1160
rect 526 1124 538 1160
rect 318 1118 324 1124
rect 524 1118 538 1124
rect 318 1038 322 1118
rect 526 1038 538 1118
rect 318 1032 324 1038
rect 524 1032 538 1038
rect 318 996 322 1032
rect 526 996 538 1032
rect 318 990 324 996
rect 524 990 538 996
rect 318 908 322 990
rect 526 908 538 990
rect 318 902 324 908
rect 524 902 538 908
rect 62 432 76 438
rect 276 432 284 438
rect 62 348 74 432
rect 278 348 284 432
rect 62 342 76 348
rect 276 342 284 348
rect 62 306 74 342
rect 278 306 284 342
rect 62 300 76 306
rect 276 300 284 306
rect 62 218 74 300
rect 278 218 284 300
rect 62 212 76 218
rect 276 212 284 218
rect 62 176 74 212
rect 278 176 284 212
rect 62 170 76 176
rect 276 170 284 176
rect 62 88 74 170
rect 278 88 284 170
rect 62 82 76 88
rect 276 82 284 88
rect 316 432 324 438
rect 524 432 538 438
rect 316 348 322 432
rect 526 348 538 432
rect 316 342 324 348
rect 524 342 538 348
rect 316 306 322 342
rect 526 306 538 342
rect 316 300 324 306
rect 524 300 538 306
rect 316 218 322 300
rect 526 218 538 300
rect 316 212 324 218
rect 524 212 538 218
rect 316 176 322 212
rect 526 176 538 212
rect 316 170 324 176
rect 524 170 538 176
rect 316 88 322 170
rect 526 88 538 170
rect 316 82 324 88
rect 524 82 538 88
<< genericcontact >>
rect 4 1328 8 1332
rect 16 1328 20 1332
rect 26 1328 30 1332
rect 36 1328 40 1332
rect 46 1328 50 1332
rect 56 1328 60 1332
rect 66 1328 70 1332
rect 76 1328 80 1332
rect 86 1328 90 1332
rect 96 1328 100 1332
rect 106 1328 110 1332
rect 116 1328 120 1332
rect 126 1328 130 1332
rect 136 1328 140 1332
rect 146 1328 150 1332
rect 156 1328 160 1332
rect 166 1328 170 1332
rect 176 1328 180 1332
rect 186 1328 190 1332
rect 196 1328 200 1332
rect 206 1328 210 1332
rect 216 1328 220 1332
rect 226 1328 230 1332
rect 370 1328 374 1332
rect 380 1328 384 1332
rect 390 1328 394 1332
rect 400 1328 404 1332
rect 410 1328 414 1332
rect 420 1328 424 1332
rect 430 1328 434 1332
rect 440 1328 444 1332
rect 450 1328 454 1332
rect 460 1328 464 1332
rect 470 1328 474 1332
rect 480 1328 484 1332
rect 490 1328 494 1332
rect 500 1328 504 1332
rect 510 1328 514 1332
rect 520 1328 524 1332
rect 530 1328 534 1332
rect 540 1328 544 1332
rect 550 1328 554 1332
rect 560 1328 564 1332
rect 570 1328 574 1332
rect 582 1326 586 1330
rect 592 1326 596 1330
rect 4 1318 8 1322
rect 16 1318 20 1322
rect 26 1318 30 1322
rect 36 1318 40 1322
rect 46 1318 50 1322
rect 56 1318 60 1322
rect 66 1318 70 1322
rect 76 1318 80 1322
rect 86 1318 90 1322
rect 96 1318 100 1322
rect 106 1318 110 1322
rect 116 1318 120 1322
rect 126 1318 130 1322
rect 136 1318 140 1322
rect 146 1318 150 1322
rect 156 1318 160 1322
rect 166 1318 170 1322
rect 176 1318 180 1322
rect 186 1318 190 1322
rect 196 1318 200 1322
rect 206 1318 210 1322
rect 216 1318 220 1322
rect 226 1318 230 1322
rect 370 1318 374 1322
rect 380 1318 384 1322
rect 390 1318 394 1322
rect 400 1318 404 1322
rect 410 1318 414 1322
rect 420 1318 424 1322
rect 430 1318 434 1322
rect 440 1318 444 1322
rect 450 1318 454 1322
rect 460 1318 464 1322
rect 470 1318 474 1322
rect 480 1318 484 1322
rect 490 1318 494 1322
rect 500 1318 504 1322
rect 510 1318 514 1322
rect 520 1318 524 1322
rect 530 1318 534 1322
rect 540 1318 544 1322
rect 550 1318 554 1322
rect 560 1318 564 1322
rect 570 1318 574 1322
rect 582 1316 586 1320
rect 592 1316 596 1320
rect 4 1308 8 1312
rect 14 1308 18 1312
rect 582 1306 586 1310
rect 592 1306 596 1310
rect 4 1298 8 1302
rect 14 1298 18 1302
rect 582 1296 586 1300
rect 592 1296 596 1300
rect 4 1288 8 1292
rect 14 1288 18 1292
rect 298 1288 302 1292
rect 92 1284 96 1288
rect 102 1284 106 1288
rect 114 1284 118 1288
rect 134 1284 138 1288
rect 144 1284 148 1288
rect 164 1284 168 1288
rect 174 1284 178 1288
rect 194 1284 198 1288
rect 204 1284 208 1288
rect 224 1284 228 1288
rect 368 1284 372 1288
rect 388 1284 392 1288
rect 398 1284 402 1288
rect 418 1284 422 1288
rect 428 1284 432 1288
rect 448 1284 452 1288
rect 458 1284 462 1288
rect 478 1284 482 1288
rect 490 1284 494 1288
rect 500 1284 504 1288
rect 582 1286 586 1290
rect 592 1286 596 1290
rect 4 1278 8 1282
rect 14 1278 18 1282
rect 42 1274 46 1278
rect 52 1274 56 1278
rect 92 1274 96 1278
rect 102 1274 106 1278
rect 114 1274 118 1278
rect 134 1274 138 1278
rect 144 1274 148 1278
rect 164 1274 168 1278
rect 174 1274 178 1278
rect 194 1274 198 1278
rect 204 1274 208 1278
rect 224 1274 228 1278
rect 368 1274 372 1278
rect 388 1274 392 1278
rect 398 1274 402 1278
rect 418 1274 422 1278
rect 428 1274 432 1278
rect 448 1274 452 1278
rect 458 1274 462 1278
rect 478 1274 482 1278
rect 490 1274 494 1278
rect 500 1274 504 1278
rect 544 1274 548 1278
rect 554 1274 558 1278
rect 582 1276 586 1280
rect 592 1276 596 1280
rect 4 1268 8 1272
rect 14 1268 18 1272
rect 298 1268 302 1272
rect 42 1264 46 1268
rect 52 1264 56 1268
rect 92 1264 96 1268
rect 102 1264 106 1268
rect 114 1264 118 1268
rect 134 1264 138 1268
rect 144 1264 148 1268
rect 164 1264 168 1268
rect 174 1264 178 1268
rect 194 1264 198 1268
rect 204 1264 208 1268
rect 224 1264 228 1268
rect 368 1264 372 1268
rect 388 1264 392 1268
rect 398 1264 402 1268
rect 418 1264 422 1268
rect 428 1264 432 1268
rect 448 1264 452 1268
rect 458 1264 462 1268
rect 478 1264 482 1268
rect 490 1264 494 1268
rect 500 1264 504 1268
rect 544 1264 548 1268
rect 554 1264 558 1268
rect 582 1266 586 1270
rect 592 1266 596 1270
rect 4 1258 8 1262
rect 14 1258 18 1262
rect 298 1258 302 1262
rect 42 1254 46 1258
rect 52 1254 56 1258
rect 544 1254 548 1258
rect 554 1254 558 1258
rect 582 1256 586 1260
rect 592 1256 596 1260
rect 4 1248 8 1252
rect 14 1248 18 1252
rect 298 1248 302 1252
rect 582 1246 586 1250
rect 592 1246 596 1250
rect 4 1238 8 1242
rect 14 1238 18 1242
rect 42 1234 46 1238
rect 52 1234 56 1238
rect 544 1234 548 1238
rect 554 1234 558 1238
rect 582 1236 586 1240
rect 592 1236 596 1240
rect 4 1228 8 1232
rect 14 1228 18 1232
rect 298 1228 302 1232
rect 42 1224 46 1228
rect 52 1224 56 1228
rect 66 1222 70 1226
rect 544 1224 548 1228
rect 554 1224 558 1228
rect 582 1226 586 1230
rect 592 1226 596 1230
rect 4 1218 8 1222
rect 14 1218 18 1222
rect 298 1218 302 1222
rect 530 1219 534 1223
rect 42 1214 46 1218
rect 52 1214 56 1218
rect 66 1212 70 1216
rect 544 1214 548 1218
rect 554 1214 558 1218
rect 582 1216 586 1220
rect 592 1216 596 1220
rect 4 1208 8 1212
rect 14 1208 18 1212
rect 114 1210 118 1214
rect 124 1210 128 1214
rect 134 1210 138 1214
rect 144 1210 148 1214
rect 154 1210 158 1214
rect 164 1210 168 1214
rect 174 1210 178 1214
rect 184 1210 188 1214
rect 194 1210 198 1214
rect 204 1210 208 1214
rect 214 1210 218 1214
rect 224 1210 228 1214
rect 234 1210 238 1214
rect 298 1208 302 1212
rect 362 1210 366 1214
rect 372 1210 376 1214
rect 382 1210 386 1214
rect 392 1210 396 1214
rect 402 1210 406 1214
rect 412 1210 416 1214
rect 422 1210 426 1214
rect 432 1210 436 1214
rect 442 1210 446 1214
rect 452 1210 456 1214
rect 462 1210 466 1214
rect 472 1210 476 1214
rect 482 1210 486 1214
rect 530 1209 534 1213
rect 582 1206 586 1210
rect 592 1206 596 1210
rect 66 1202 70 1206
rect 4 1198 8 1202
rect 14 1198 18 1202
rect 114 1200 118 1204
rect 124 1200 128 1204
rect 134 1200 138 1204
rect 144 1200 148 1204
rect 154 1200 158 1204
rect 164 1200 168 1204
rect 174 1200 178 1204
rect 184 1200 188 1204
rect 194 1200 198 1204
rect 204 1200 208 1204
rect 214 1200 218 1204
rect 224 1200 228 1204
rect 234 1200 238 1204
rect 362 1200 366 1204
rect 372 1200 376 1204
rect 382 1200 386 1204
rect 392 1200 396 1204
rect 402 1200 406 1204
rect 412 1200 416 1204
rect 422 1200 426 1204
rect 432 1200 436 1204
rect 442 1200 446 1204
rect 452 1200 456 1204
rect 462 1200 466 1204
rect 472 1200 476 1204
rect 482 1200 486 1204
rect 530 1199 534 1203
rect 42 1194 46 1198
rect 52 1194 56 1198
rect 66 1192 70 1196
rect 544 1194 548 1198
rect 554 1194 558 1198
rect 582 1196 586 1200
rect 592 1196 596 1200
rect 4 1188 8 1192
rect 14 1188 18 1192
rect 298 1188 302 1192
rect 530 1189 534 1193
rect 42 1184 46 1188
rect 52 1184 56 1188
rect 544 1184 548 1188
rect 554 1184 558 1188
rect 582 1186 586 1190
rect 592 1186 596 1190
rect 4 1178 8 1182
rect 14 1178 18 1182
rect 298 1178 302 1182
rect 42 1174 46 1178
rect 52 1174 56 1178
rect 544 1174 548 1178
rect 554 1174 558 1178
rect 582 1176 586 1180
rect 592 1176 596 1180
rect 4 1168 8 1172
rect 14 1168 18 1172
rect 298 1168 302 1172
rect 582 1166 586 1170
rect 592 1166 596 1170
rect 4 1158 8 1162
rect 14 1158 18 1162
rect 42 1154 46 1158
rect 52 1154 56 1158
rect 544 1154 548 1158
rect 554 1154 558 1158
rect 582 1156 586 1160
rect 592 1156 596 1160
rect 4 1148 8 1152
rect 14 1148 18 1152
rect 42 1144 46 1148
rect 52 1144 56 1148
rect 125 1146 129 1150
rect 135 1146 139 1150
rect 155 1146 159 1150
rect 165 1146 169 1150
rect 185 1146 189 1150
rect 195 1146 199 1150
rect 215 1146 219 1150
rect 225 1146 229 1150
rect 298 1148 302 1152
rect 370 1146 374 1150
rect 380 1146 384 1150
rect 400 1146 404 1150
rect 410 1146 414 1150
rect 430 1146 434 1150
rect 440 1146 444 1150
rect 460 1146 464 1150
rect 470 1146 474 1150
rect 544 1144 548 1148
rect 554 1144 558 1148
rect 582 1146 586 1150
rect 592 1146 596 1150
rect 4 1138 8 1142
rect 14 1138 18 1142
rect 298 1138 302 1142
rect 42 1134 46 1138
rect 52 1134 56 1138
rect 125 1134 129 1138
rect 135 1134 139 1138
rect 155 1134 159 1138
rect 165 1134 169 1138
rect 185 1134 189 1138
rect 195 1134 199 1138
rect 215 1134 219 1138
rect 225 1134 229 1138
rect 370 1134 374 1138
rect 380 1134 384 1138
rect 400 1134 404 1138
rect 410 1134 414 1138
rect 430 1134 434 1138
rect 440 1134 444 1138
rect 460 1134 464 1138
rect 470 1134 474 1138
rect 544 1134 548 1138
rect 554 1134 558 1138
rect 582 1136 586 1140
rect 592 1136 596 1140
rect 4 1128 8 1132
rect 14 1128 18 1132
rect 298 1128 302 1132
rect 582 1126 586 1130
rect 592 1126 596 1130
rect 4 1118 8 1122
rect 14 1118 18 1122
rect 42 1114 46 1118
rect 52 1114 56 1118
rect 544 1114 548 1118
rect 554 1114 558 1118
rect 582 1116 586 1120
rect 592 1116 596 1120
rect 4 1108 8 1112
rect 14 1108 18 1112
rect 298 1108 302 1112
rect 42 1104 46 1108
rect 52 1104 56 1108
rect 544 1104 548 1108
rect 554 1104 558 1108
rect 582 1106 586 1110
rect 592 1106 596 1110
rect 4 1098 8 1102
rect 14 1098 18 1102
rect 298 1098 302 1102
rect 42 1094 46 1098
rect 52 1094 56 1098
rect 66 1092 70 1096
rect 530 1092 534 1096
rect 544 1094 548 1098
rect 554 1094 558 1098
rect 582 1096 586 1100
rect 592 1096 596 1100
rect 4 1088 8 1092
rect 14 1088 18 1092
rect 298 1088 302 1092
rect 582 1086 586 1090
rect 592 1086 596 1090
rect 66 1082 70 1086
rect 4 1078 8 1082
rect 14 1078 18 1082
rect 114 1081 118 1085
rect 124 1081 128 1085
rect 134 1081 138 1085
rect 144 1081 148 1085
rect 154 1081 158 1085
rect 164 1081 168 1085
rect 174 1081 178 1085
rect 184 1081 188 1085
rect 194 1081 198 1085
rect 204 1081 208 1085
rect 214 1081 218 1085
rect 224 1081 228 1085
rect 234 1081 238 1085
rect 362 1081 366 1085
rect 372 1081 376 1085
rect 382 1081 386 1085
rect 392 1081 396 1085
rect 402 1081 406 1085
rect 412 1081 416 1085
rect 422 1081 426 1085
rect 432 1081 436 1085
rect 442 1081 446 1085
rect 452 1081 456 1085
rect 462 1081 466 1085
rect 472 1081 476 1085
rect 482 1081 486 1085
rect 530 1082 534 1086
rect 42 1074 46 1078
rect 52 1074 56 1078
rect 66 1072 70 1076
rect 4 1068 8 1072
rect 14 1068 18 1072
rect 114 1071 118 1075
rect 124 1071 128 1075
rect 134 1071 138 1075
rect 144 1071 148 1075
rect 154 1071 158 1075
rect 164 1071 168 1075
rect 174 1071 178 1075
rect 184 1071 188 1075
rect 194 1071 198 1075
rect 204 1071 208 1075
rect 214 1071 218 1075
rect 224 1071 228 1075
rect 234 1071 238 1075
rect 298 1068 302 1072
rect 362 1071 366 1075
rect 372 1071 376 1075
rect 382 1071 386 1075
rect 392 1071 396 1075
rect 402 1071 406 1075
rect 412 1071 416 1075
rect 422 1071 426 1075
rect 432 1071 436 1075
rect 442 1071 446 1075
rect 452 1071 456 1075
rect 462 1071 466 1075
rect 472 1071 476 1075
rect 482 1071 486 1075
rect 530 1072 534 1076
rect 544 1074 548 1078
rect 554 1074 558 1078
rect 582 1076 586 1080
rect 592 1076 596 1080
rect 42 1064 46 1068
rect 52 1064 56 1068
rect 66 1062 70 1066
rect 530 1062 534 1066
rect 544 1064 548 1068
rect 554 1064 558 1068
rect 582 1066 586 1070
rect 592 1066 596 1070
rect 4 1058 8 1062
rect 14 1058 18 1062
rect 298 1058 302 1062
rect 42 1054 46 1058
rect 52 1054 56 1058
rect 544 1054 548 1058
rect 554 1054 558 1058
rect 582 1056 586 1060
rect 592 1056 596 1060
rect 4 1048 8 1052
rect 14 1048 18 1052
rect 298 1048 302 1052
rect 582 1046 586 1050
rect 592 1046 596 1050
rect 4 1038 8 1042
rect 14 1038 18 1042
rect 42 1034 46 1038
rect 52 1034 56 1038
rect 544 1034 548 1038
rect 554 1034 558 1038
rect 582 1036 586 1040
rect 592 1036 596 1040
rect 4 1028 8 1032
rect 14 1028 18 1032
rect 298 1028 302 1032
rect 42 1024 46 1028
rect 52 1024 56 1028
rect 544 1024 548 1028
rect 554 1024 558 1028
rect 582 1026 586 1030
rect 592 1026 596 1030
rect 4 1018 8 1022
rect 14 1018 18 1022
rect 124 1018 128 1022
rect 134 1018 138 1022
rect 154 1018 158 1022
rect 164 1018 168 1022
rect 184 1018 188 1022
rect 194 1018 198 1022
rect 214 1018 218 1022
rect 224 1018 228 1022
rect 298 1018 302 1022
rect 369 1018 373 1022
rect 379 1018 383 1022
rect 399 1018 403 1022
rect 409 1018 413 1022
rect 429 1018 433 1022
rect 439 1018 443 1022
rect 459 1018 463 1022
rect 469 1018 473 1022
rect 42 1014 46 1018
rect 52 1014 56 1018
rect 544 1014 548 1018
rect 554 1014 558 1018
rect 582 1016 586 1020
rect 592 1016 596 1020
rect 4 1008 8 1012
rect 14 1008 18 1012
rect 124 1006 128 1010
rect 134 1006 138 1010
rect 154 1006 158 1010
rect 164 1006 168 1010
rect 184 1006 188 1010
rect 194 1006 198 1010
rect 214 1006 218 1010
rect 224 1006 228 1010
rect 298 1008 302 1012
rect 369 1006 373 1010
rect 379 1006 383 1010
rect 399 1006 403 1010
rect 409 1006 413 1010
rect 429 1006 433 1010
rect 439 1006 443 1010
rect 459 1006 463 1010
rect 469 1006 473 1010
rect 582 1006 586 1010
rect 592 1006 596 1010
rect 4 998 8 1002
rect 14 998 18 1002
rect 42 994 46 998
rect 52 994 56 998
rect 544 994 548 998
rect 554 994 558 998
rect 582 996 586 1000
rect 592 996 596 1000
rect 4 988 8 992
rect 14 988 18 992
rect 298 988 302 992
rect 42 984 46 988
rect 52 984 56 988
rect 544 984 548 988
rect 554 984 558 988
rect 582 986 586 990
rect 592 986 596 990
rect 4 978 8 982
rect 14 978 18 982
rect 298 978 302 982
rect 42 974 46 978
rect 52 974 56 978
rect 544 974 548 978
rect 554 974 558 978
rect 582 976 586 980
rect 592 976 596 980
rect 4 968 8 972
rect 14 968 18 972
rect 298 968 302 972
rect 582 966 586 970
rect 592 966 596 970
rect 530 962 534 966
rect 4 958 8 962
rect 14 958 18 962
rect 42 954 46 958
rect 52 954 56 958
rect 66 956 70 960
rect 114 952 118 956
rect 124 952 128 956
rect 134 952 138 956
rect 144 952 148 956
rect 154 952 158 956
rect 164 952 168 956
rect 174 952 178 956
rect 184 952 188 956
rect 194 952 198 956
rect 204 952 208 956
rect 214 952 218 956
rect 224 952 228 956
rect 234 952 238 956
rect 362 952 366 956
rect 372 952 376 956
rect 382 952 386 956
rect 392 952 396 956
rect 402 952 406 956
rect 412 952 416 956
rect 422 952 426 956
rect 432 952 436 956
rect 442 952 446 956
rect 452 952 456 956
rect 462 952 466 956
rect 472 952 476 956
rect 482 952 486 956
rect 530 952 534 956
rect 544 954 548 958
rect 554 954 558 958
rect 582 956 586 960
rect 592 956 596 960
rect 4 948 8 952
rect 14 948 18 952
rect 42 944 46 948
rect 52 944 56 948
rect 66 946 70 950
rect 298 948 302 952
rect 114 942 118 946
rect 124 942 128 946
rect 134 942 138 946
rect 144 942 148 946
rect 154 942 158 946
rect 164 942 168 946
rect 174 942 178 946
rect 184 942 188 946
rect 194 942 198 946
rect 204 942 208 946
rect 214 942 218 946
rect 224 942 228 946
rect 234 942 238 946
rect 362 942 366 946
rect 372 942 376 946
rect 382 942 386 946
rect 392 942 396 946
rect 402 942 406 946
rect 412 942 416 946
rect 422 942 426 946
rect 432 942 436 946
rect 442 942 446 946
rect 452 942 456 946
rect 462 942 466 946
rect 472 942 476 946
rect 482 942 486 946
rect 530 942 534 946
rect 544 944 548 948
rect 554 944 558 948
rect 582 946 586 950
rect 592 946 596 950
rect 4 938 8 942
rect 14 938 18 942
rect 42 934 46 938
rect 52 934 56 938
rect 66 936 70 940
rect 298 938 302 942
rect 530 932 534 936
rect 544 934 548 938
rect 554 934 558 938
rect 582 936 586 940
rect 592 936 596 940
rect 4 928 8 932
rect 14 928 18 932
rect 66 926 70 930
rect 298 928 302 932
rect 582 926 586 930
rect 592 926 596 930
rect 530 922 534 926
rect 4 918 8 922
rect 14 918 18 922
rect 42 914 46 918
rect 52 914 56 918
rect 66 916 70 920
rect 530 912 534 916
rect 544 914 548 918
rect 554 914 558 918
rect 582 916 586 920
rect 592 916 596 920
rect 4 908 8 912
rect 14 908 18 912
rect 42 904 46 908
rect 52 904 56 908
rect 66 906 70 910
rect 298 908 302 912
rect 544 904 548 908
rect 554 904 558 908
rect 582 906 586 910
rect 592 906 596 910
rect 4 898 8 902
rect 14 898 18 902
rect 298 898 302 902
rect 42 894 46 898
rect 52 894 56 898
rect 544 894 548 898
rect 554 894 558 898
rect 582 896 586 900
rect 592 896 596 900
rect 4 888 8 892
rect 14 888 18 892
rect 125 888 129 892
rect 135 888 139 892
rect 155 888 159 892
rect 165 888 169 892
rect 185 888 189 892
rect 195 888 199 892
rect 215 888 219 892
rect 225 888 229 892
rect 298 888 302 892
rect 371 888 375 892
rect 381 888 385 892
rect 401 888 405 892
rect 411 888 415 892
rect 431 888 435 892
rect 441 888 445 892
rect 461 888 465 892
rect 471 888 475 892
rect 582 886 586 890
rect 592 886 596 890
rect 4 878 8 882
rect 14 878 18 882
rect 42 874 46 878
rect 52 874 56 878
rect 105 876 109 880
rect 125 876 129 880
rect 135 876 139 880
rect 155 876 159 880
rect 165 876 169 880
rect 185 876 189 880
rect 195 876 199 880
rect 215 876 219 880
rect 225 876 229 880
rect 371 876 375 880
rect 381 876 385 880
rect 401 876 405 880
rect 411 876 415 880
rect 431 876 435 880
rect 441 876 445 880
rect 461 876 465 880
rect 471 876 475 880
rect 491 876 495 880
rect 544 874 548 878
rect 554 874 558 878
rect 582 876 586 880
rect 592 876 596 880
rect 4 868 8 872
rect 14 868 18 872
rect 298 868 302 872
rect 42 864 46 868
rect 52 864 56 868
rect 95 864 99 868
rect 105 864 109 868
rect 115 864 119 868
rect 125 864 129 868
rect 135 864 139 868
rect 145 864 149 868
rect 155 864 159 868
rect 165 864 169 868
rect 175 864 179 868
rect 185 864 189 868
rect 195 864 199 868
rect 205 864 209 868
rect 215 864 219 868
rect 225 864 229 868
rect 371 864 375 868
rect 381 864 385 868
rect 391 864 395 868
rect 401 864 405 868
rect 411 864 415 868
rect 421 864 425 868
rect 431 864 435 868
rect 441 864 445 868
rect 451 864 455 868
rect 461 864 465 868
rect 471 864 475 868
rect 481 864 485 868
rect 491 864 495 868
rect 501 864 505 868
rect 544 864 548 868
rect 554 864 558 868
rect 582 866 586 870
rect 592 866 596 870
rect 4 858 8 862
rect 14 858 18 862
rect 582 856 586 860
rect 592 856 596 860
rect 4 848 8 852
rect 14 848 18 852
rect 582 846 586 850
rect 592 846 596 850
rect 4 838 8 842
rect 14 838 18 842
rect 32 833 36 837
rect 42 833 46 837
rect 52 833 56 837
rect 80 833 84 837
rect 90 833 94 837
rect 100 833 104 837
rect 110 833 114 837
rect 120 833 124 837
rect 130 833 134 837
rect 140 833 144 837
rect 150 833 154 837
rect 160 833 164 837
rect 170 833 174 837
rect 180 833 184 837
rect 190 833 194 837
rect 200 833 204 837
rect 210 833 214 837
rect 220 833 224 837
rect 298 833 302 837
rect 370 833 374 837
rect 380 833 384 837
rect 390 833 394 837
rect 400 833 404 837
rect 410 833 414 837
rect 420 833 424 837
rect 430 833 434 837
rect 440 833 444 837
rect 450 833 454 837
rect 460 833 464 837
rect 470 833 474 837
rect 480 833 484 837
rect 490 833 494 837
rect 500 833 504 837
rect 510 833 514 837
rect 550 833 554 837
rect 560 833 564 837
rect 570 833 574 837
rect 582 836 586 840
rect 592 836 596 840
rect 4 828 8 832
rect 14 828 18 832
rect 32 823 36 827
rect 42 823 46 827
rect 52 823 56 827
rect 80 823 84 827
rect 90 823 94 827
rect 100 823 104 827
rect 110 823 114 827
rect 120 823 124 827
rect 130 823 134 827
rect 140 823 144 827
rect 150 823 154 827
rect 160 823 164 827
rect 170 823 174 827
rect 180 823 184 827
rect 190 823 194 827
rect 200 823 204 827
rect 210 823 214 827
rect 220 823 224 827
rect 298 823 302 827
rect 370 823 374 827
rect 380 823 384 827
rect 390 823 394 827
rect 400 823 404 827
rect 410 823 414 827
rect 420 823 424 827
rect 430 823 434 827
rect 440 823 444 827
rect 450 823 454 827
rect 460 823 464 827
rect 470 823 474 827
rect 480 823 484 827
rect 490 823 494 827
rect 500 823 504 827
rect 510 823 514 827
rect 550 823 554 827
rect 560 823 564 827
rect 570 823 574 827
rect 582 826 586 830
rect 592 826 596 830
rect 4 808 8 812
rect 592 807 596 811
rect 4 798 8 802
rect 4 788 8 792
rect 592 787 596 791
rect 4 778 8 782
rect 4 768 8 772
rect 592 767 596 771
rect 4 758 8 762
rect 4 748 8 752
rect 592 747 596 751
rect 4 738 8 742
rect 4 728 8 732
rect 592 727 596 731
rect 4 718 8 722
rect 4 708 8 712
rect 592 707 596 711
rect 4 698 8 702
rect 4 688 8 692
rect 36 688 40 692
rect 92 687 96 691
rect 130 687 134 691
rect 140 687 144 691
rect 150 687 154 691
rect 160 687 164 691
rect 200 689 204 693
rect 218 689 222 693
rect 390 687 394 691
rect 400 687 404 691
rect 410 687 414 691
rect 420 687 424 691
rect 448 688 452 692
rect 486 687 490 691
rect 496 687 500 691
rect 516 687 520 691
rect 544 686 548 690
rect 582 687 586 691
rect 592 687 596 691
rect 4 656 8 660
rect 36 657 40 661
rect 92 657 96 661
rect 130 657 134 661
rect 150 657 154 661
rect 160 657 164 661
rect 198 657 202 661
rect 220 657 224 661
rect 390 657 394 661
rect 400 657 404 661
rect 420 657 424 661
rect 448 657 452 661
rect 486 657 490 661
rect 496 657 500 661
rect 516 657 520 661
rect 544 657 548 661
rect 582 658 586 662
rect 592 658 596 662
rect 4 646 8 650
rect 592 648 596 652
rect 4 626 8 630
rect 592 628 596 632
rect 4 606 8 610
rect 592 608 596 612
rect 4 586 8 590
rect 592 588 596 592
rect 4 566 8 570
rect 592 568 596 572
rect 4 546 8 550
rect 592 548 596 552
rect 4 526 8 530
rect 592 528 596 532
rect 120 520 124 524
rect 130 520 134 524
rect 140 520 144 524
rect 150 520 154 524
rect 160 520 164 524
rect 170 520 174 524
rect 180 520 184 524
rect 190 520 194 524
rect 200 520 204 524
rect 210 520 214 524
rect 220 520 224 524
rect 388 523 392 527
rect 484 523 488 527
rect 6 506 10 510
rect 110 508 114 512
rect 120 508 124 512
rect 130 508 134 512
rect 140 508 144 512
rect 150 508 154 512
rect 160 508 164 512
rect 170 508 174 512
rect 180 508 184 512
rect 190 508 194 512
rect 200 508 204 512
rect 210 508 214 512
rect 220 510 224 514
rect 391 510 395 514
rect 401 510 405 514
rect 411 510 415 514
rect 421 510 425 514
rect 431 510 435 514
rect 441 510 445 514
rect 451 510 455 514
rect 482 513 486 517
rect 492 513 496 517
rect 502 513 506 517
rect 552 515 556 519
rect 562 515 566 519
rect 572 515 576 519
rect 582 515 586 519
rect 592 506 596 510
rect 6 496 10 500
rect 582 496 586 500
rect 592 496 596 500
rect 6 486 10 490
rect 582 486 586 490
rect 592 486 596 490
rect 6 476 10 480
rect 36 478 40 482
rect 46 478 50 482
rect 108 480 112 484
rect 118 480 122 484
rect 128 480 132 484
rect 138 480 142 484
rect 148 480 152 484
rect 158 480 162 484
rect 168 480 172 484
rect 178 480 182 484
rect 188 480 192 484
rect 198 480 202 484
rect 208 480 212 484
rect 218 480 222 484
rect 228 480 232 484
rect 366 480 370 484
rect 376 480 380 484
rect 386 480 390 484
rect 396 480 400 484
rect 406 480 410 484
rect 416 480 420 484
rect 426 480 430 484
rect 436 480 440 484
rect 446 480 450 484
rect 456 480 460 484
rect 466 480 470 484
rect 476 480 480 484
rect 486 480 490 484
rect 544 478 548 482
rect 554 478 558 482
rect 582 476 586 480
rect 592 476 596 480
rect 6 466 10 470
rect 36 468 40 472
rect 46 468 50 472
rect 108 470 112 474
rect 118 470 122 474
rect 128 470 132 474
rect 138 470 142 474
rect 148 470 152 474
rect 158 470 162 474
rect 168 470 172 474
rect 178 470 182 474
rect 188 470 192 474
rect 198 470 202 474
rect 208 470 212 474
rect 218 470 222 474
rect 228 470 232 474
rect 298 472 302 476
rect 366 470 370 474
rect 376 470 380 474
rect 386 470 390 474
rect 396 470 400 474
rect 406 470 410 474
rect 416 470 420 474
rect 426 470 430 474
rect 436 470 440 474
rect 446 470 450 474
rect 456 470 460 474
rect 466 470 470 474
rect 476 470 480 474
rect 486 470 490 474
rect 544 468 548 472
rect 554 468 558 472
rect 582 466 586 470
rect 592 466 596 470
rect 6 456 10 460
rect 36 458 40 462
rect 46 458 50 462
rect 110 460 114 464
rect 120 460 124 464
rect 140 460 144 464
rect 150 460 154 464
rect 170 460 174 464
rect 180 460 184 464
rect 200 460 204 464
rect 210 460 214 464
rect 230 460 234 464
rect 298 462 302 466
rect 366 460 370 464
rect 376 460 380 464
rect 396 460 400 464
rect 406 460 410 464
rect 426 460 430 464
rect 436 460 440 464
rect 456 460 460 464
rect 466 460 470 464
rect 486 460 490 464
rect 544 455 548 459
rect 554 455 558 459
rect 582 456 586 460
rect 592 456 596 460
rect 6 446 10 450
rect 110 448 114 452
rect 120 448 124 452
rect 140 448 144 452
rect 150 448 154 452
rect 170 448 174 452
rect 180 448 184 452
rect 200 448 204 452
rect 210 448 214 452
rect 230 448 234 452
rect 366 448 370 452
rect 376 448 380 452
rect 396 448 400 452
rect 406 448 410 452
rect 426 448 430 452
rect 436 448 440 452
rect 456 448 460 452
rect 466 448 470 452
rect 486 448 490 452
rect 582 446 586 450
rect 592 446 596 450
rect 298 442 302 446
rect 6 436 10 440
rect 36 438 40 442
rect 46 438 50 442
rect 298 432 302 436
rect 544 435 548 439
rect 554 435 558 439
rect 582 436 586 440
rect 592 436 596 440
rect 6 426 10 430
rect 36 428 40 432
rect 46 428 50 432
rect 66 428 70 432
rect 530 428 534 432
rect 544 425 548 429
rect 554 425 558 429
rect 582 426 586 430
rect 592 426 596 430
rect 6 416 10 420
rect 36 418 40 422
rect 46 418 50 422
rect 66 418 70 422
rect 530 418 534 422
rect 298 412 302 416
rect 544 415 548 419
rect 554 415 558 419
rect 582 416 586 420
rect 592 416 596 420
rect 6 406 10 410
rect 66 408 70 412
rect 530 408 534 412
rect 582 406 586 410
rect 592 406 596 410
rect 298 402 302 406
rect 6 396 10 400
rect 36 398 40 402
rect 46 398 50 402
rect 66 398 70 402
rect 530 398 534 402
rect 114 394 118 398
rect 124 394 128 398
rect 134 394 138 398
rect 144 394 148 398
rect 154 394 158 398
rect 164 394 168 398
rect 174 394 178 398
rect 184 394 188 398
rect 194 394 198 398
rect 204 394 208 398
rect 214 394 218 398
rect 224 394 228 398
rect 234 394 238 398
rect 362 394 366 398
rect 372 394 376 398
rect 382 394 386 398
rect 392 394 396 398
rect 402 394 406 398
rect 412 394 416 398
rect 422 394 426 398
rect 432 394 436 398
rect 442 394 446 398
rect 452 394 456 398
rect 462 394 466 398
rect 472 394 476 398
rect 482 394 486 398
rect 544 395 548 399
rect 554 395 558 399
rect 582 396 586 400
rect 592 396 596 400
rect 6 386 10 390
rect 36 388 40 392
rect 46 388 50 392
rect 66 388 70 392
rect 530 388 534 392
rect 114 382 118 386
rect 124 382 128 386
rect 134 382 138 386
rect 144 382 148 386
rect 154 382 158 386
rect 164 382 168 386
rect 174 382 178 386
rect 184 382 188 386
rect 194 382 198 386
rect 204 382 208 386
rect 214 382 218 386
rect 224 382 228 386
rect 234 382 238 386
rect 298 382 302 386
rect 362 382 366 386
rect 372 382 376 386
rect 382 382 386 386
rect 392 382 396 386
rect 402 382 406 386
rect 412 382 416 386
rect 422 382 426 386
rect 432 382 436 386
rect 442 382 446 386
rect 452 382 456 386
rect 462 382 466 386
rect 472 382 476 386
rect 482 382 486 386
rect 544 385 548 389
rect 554 385 558 389
rect 582 386 586 390
rect 592 386 596 390
rect 6 376 10 380
rect 36 378 40 382
rect 46 378 50 382
rect 66 378 70 382
rect 530 378 534 382
rect 298 372 302 376
rect 544 375 548 379
rect 554 375 558 379
rect 582 376 586 380
rect 592 376 596 380
rect 6 366 10 370
rect 66 368 70 372
rect 530 368 534 372
rect 582 366 586 370
rect 592 366 596 370
rect 6 356 10 360
rect 36 358 40 362
rect 46 358 50 362
rect 66 358 70 362
rect 530 358 534 362
rect 298 352 302 356
rect 544 355 548 359
rect 554 355 558 359
rect 582 356 586 360
rect 592 356 596 360
rect 6 346 10 350
rect 36 348 40 352
rect 46 348 50 352
rect 66 348 70 352
rect 530 348 534 352
rect 298 342 302 346
rect 544 345 548 349
rect 554 345 558 349
rect 582 346 586 350
rect 592 346 596 350
rect 6 336 10 340
rect 36 338 40 342
rect 46 338 50 342
rect 66 338 70 342
rect 530 338 534 342
rect 544 335 548 339
rect 554 335 558 339
rect 582 336 586 340
rect 592 336 596 340
rect 6 326 10 330
rect 66 328 70 332
rect 112 328 116 332
rect 122 328 126 332
rect 142 328 146 332
rect 152 328 156 332
rect 172 328 176 332
rect 182 328 186 332
rect 202 328 206 332
rect 212 328 216 332
rect 232 328 236 332
rect 365 329 369 333
rect 375 329 379 333
rect 395 329 399 333
rect 405 329 409 333
rect 425 329 429 333
rect 435 329 439 333
rect 455 329 459 333
rect 465 329 469 333
rect 485 329 489 333
rect 530 328 534 332
rect 582 326 586 330
rect 592 326 596 330
rect 298 322 302 326
rect 6 316 10 320
rect 36 318 40 322
rect 46 318 50 322
rect 66 318 70 322
rect 112 316 116 320
rect 122 316 126 320
rect 142 316 146 320
rect 152 316 156 320
rect 172 316 176 320
rect 182 316 186 320
rect 202 316 206 320
rect 212 316 216 320
rect 232 316 236 320
rect 365 317 369 321
rect 375 317 379 321
rect 395 317 399 321
rect 405 317 409 321
rect 425 317 429 321
rect 435 317 439 321
rect 455 317 459 321
rect 465 317 469 321
rect 485 317 489 321
rect 530 318 534 322
rect 298 312 302 316
rect 544 315 548 319
rect 554 315 558 319
rect 582 316 586 320
rect 592 316 596 320
rect 6 306 10 310
rect 36 308 40 312
rect 46 308 50 312
rect 66 308 70 312
rect 530 308 534 312
rect 544 305 548 309
rect 554 305 558 309
rect 582 306 586 310
rect 592 306 596 310
rect 6 296 10 300
rect 36 298 40 302
rect 46 298 50 302
rect 66 298 70 302
rect 530 298 534 302
rect 544 295 548 299
rect 554 295 558 299
rect 582 296 586 300
rect 592 296 596 300
rect 6 286 10 290
rect 66 288 70 292
rect 530 288 534 292
rect 582 286 586 290
rect 592 286 596 290
rect 298 282 302 286
rect 6 276 10 280
rect 36 278 40 282
rect 46 278 50 282
rect 66 278 70 282
rect 530 278 534 282
rect 544 275 548 279
rect 554 275 558 279
rect 582 276 586 280
rect 592 276 596 280
rect 6 266 10 270
rect 36 268 40 272
rect 46 268 50 272
rect 66 268 70 272
rect 530 268 534 272
rect 114 262 118 266
rect 124 262 128 266
rect 134 262 138 266
rect 144 262 148 266
rect 154 262 158 266
rect 164 262 168 266
rect 174 262 178 266
rect 184 262 188 266
rect 194 262 198 266
rect 204 262 208 266
rect 214 262 218 266
rect 224 262 228 266
rect 234 262 238 266
rect 298 262 302 266
rect 362 262 366 266
rect 372 262 376 266
rect 382 262 386 266
rect 392 262 396 266
rect 402 262 406 266
rect 412 262 416 266
rect 422 262 426 266
rect 432 262 436 266
rect 442 262 446 266
rect 452 262 456 266
rect 462 262 466 266
rect 472 262 476 266
rect 482 262 486 266
rect 544 265 548 269
rect 554 265 558 269
rect 582 266 586 270
rect 592 266 596 270
rect 6 256 10 260
rect 36 258 40 262
rect 46 258 50 262
rect 66 258 70 262
rect 530 258 534 262
rect 114 252 118 256
rect 124 252 128 256
rect 134 252 138 256
rect 144 252 148 256
rect 154 252 158 256
rect 164 252 168 256
rect 174 252 178 256
rect 184 252 188 256
rect 194 252 198 256
rect 204 252 208 256
rect 214 252 218 256
rect 224 252 228 256
rect 234 252 238 256
rect 298 252 302 256
rect 362 252 366 256
rect 372 252 376 256
rect 382 252 386 256
rect 392 252 396 256
rect 402 252 406 256
rect 412 252 416 256
rect 422 252 426 256
rect 432 252 436 256
rect 442 252 446 256
rect 452 252 456 256
rect 462 252 466 256
rect 472 252 476 256
rect 482 252 486 256
rect 544 255 548 259
rect 554 255 558 259
rect 582 256 586 260
rect 592 256 596 260
rect 6 246 10 250
rect 66 248 70 252
rect 530 248 534 252
rect 582 246 586 250
rect 592 246 596 250
rect 6 236 10 240
rect 36 238 40 242
rect 46 238 50 242
rect 66 238 70 242
rect 530 238 534 242
rect 298 232 302 236
rect 544 235 548 239
rect 554 235 558 239
rect 582 236 586 240
rect 592 236 596 240
rect 6 226 10 230
rect 36 228 40 232
rect 46 228 50 232
rect 66 228 70 232
rect 530 228 534 232
rect 298 222 302 226
rect 544 225 548 229
rect 554 225 558 229
rect 582 226 586 230
rect 592 226 596 230
rect 6 216 10 220
rect 36 218 40 222
rect 46 218 50 222
rect 66 218 70 222
rect 530 218 534 222
rect 544 215 548 219
rect 554 215 558 219
rect 582 216 586 220
rect 592 216 596 220
rect 6 206 10 210
rect 66 208 70 212
rect 530 208 534 212
rect 582 206 586 210
rect 592 206 596 210
rect 298 202 302 206
rect 6 196 10 200
rect 36 198 40 202
rect 46 198 50 202
rect 66 198 70 202
rect 111 198 115 202
rect 121 198 125 202
rect 141 198 145 202
rect 151 198 155 202
rect 171 198 175 202
rect 181 198 185 202
rect 201 198 205 202
rect 211 198 215 202
rect 231 198 235 202
rect 366 198 370 202
rect 376 198 380 202
rect 396 198 400 202
rect 406 198 410 202
rect 426 198 430 202
rect 436 198 440 202
rect 456 198 460 202
rect 466 198 470 202
rect 486 198 490 202
rect 530 198 534 202
rect 298 192 302 196
rect 544 195 548 199
rect 554 195 558 199
rect 582 196 586 200
rect 592 196 596 200
rect 6 186 10 190
rect 36 188 40 192
rect 46 188 50 192
rect 66 188 70 192
rect 111 186 115 190
rect 121 186 125 190
rect 141 186 145 190
rect 151 186 155 190
rect 171 186 175 190
rect 181 186 185 190
rect 201 186 205 190
rect 211 186 215 190
rect 231 186 235 190
rect 366 186 370 190
rect 376 186 380 190
rect 396 186 400 190
rect 406 186 410 190
rect 426 186 430 190
rect 436 186 440 190
rect 456 186 460 190
rect 466 186 470 190
rect 486 186 490 190
rect 530 188 534 192
rect 544 185 548 189
rect 554 185 558 189
rect 582 186 586 190
rect 592 186 596 190
rect 6 176 10 180
rect 36 178 40 182
rect 46 178 50 182
rect 66 178 70 182
rect 530 178 534 182
rect 298 172 302 176
rect 544 175 548 179
rect 554 175 558 179
rect 582 176 586 180
rect 592 176 596 180
rect 6 166 10 170
rect 66 168 70 172
rect 530 168 534 172
rect 582 166 586 170
rect 592 166 596 170
rect 6 156 10 160
rect 36 158 40 162
rect 46 158 50 162
rect 66 158 70 162
rect 530 158 534 162
rect 544 155 548 159
rect 554 155 558 159
rect 582 156 586 160
rect 592 156 596 160
rect 6 146 10 150
rect 36 148 40 152
rect 46 148 50 152
rect 66 148 70 152
rect 530 148 534 152
rect 298 142 302 146
rect 544 145 548 149
rect 554 145 558 149
rect 582 146 586 150
rect 592 146 596 150
rect 6 136 10 140
rect 36 138 40 142
rect 46 138 50 142
rect 66 138 70 142
rect 530 138 534 142
rect 114 132 118 136
rect 124 132 128 136
rect 134 132 138 136
rect 144 132 148 136
rect 154 132 158 136
rect 164 132 168 136
rect 174 132 178 136
rect 184 132 188 136
rect 194 132 198 136
rect 204 132 208 136
rect 214 132 218 136
rect 224 132 228 136
rect 234 132 238 136
rect 298 132 302 136
rect 362 132 366 136
rect 372 132 376 136
rect 382 132 386 136
rect 392 132 396 136
rect 402 132 406 136
rect 412 132 416 136
rect 422 132 426 136
rect 432 132 436 136
rect 442 132 446 136
rect 452 132 456 136
rect 462 132 466 136
rect 472 132 476 136
rect 482 132 486 136
rect 544 135 548 139
rect 554 135 558 139
rect 582 136 586 140
rect 592 136 596 140
rect 6 126 10 130
rect 66 128 70 132
rect 530 128 534 132
rect 582 126 586 130
rect 592 126 596 130
rect 114 122 118 126
rect 124 122 128 126
rect 134 122 138 126
rect 144 122 148 126
rect 154 122 158 126
rect 164 122 168 126
rect 174 122 178 126
rect 184 122 188 126
rect 194 122 198 126
rect 204 122 208 126
rect 214 122 218 126
rect 224 122 228 126
rect 234 122 238 126
rect 362 122 366 126
rect 372 122 376 126
rect 382 122 386 126
rect 392 122 396 126
rect 402 122 406 126
rect 412 122 416 126
rect 422 122 426 126
rect 432 122 436 126
rect 442 122 446 126
rect 452 122 456 126
rect 462 122 466 126
rect 472 122 476 126
rect 482 122 486 126
rect 6 116 10 120
rect 36 118 40 122
rect 46 118 50 122
rect 66 118 70 122
rect 530 118 534 122
rect 298 112 302 116
rect 544 115 548 119
rect 554 115 558 119
rect 582 116 586 120
rect 592 116 596 120
rect 6 106 10 110
rect 36 108 40 112
rect 46 108 50 112
rect 66 108 70 112
rect 530 108 534 112
rect 544 105 548 109
rect 554 105 558 109
rect 582 106 586 110
rect 592 106 596 110
rect 6 96 10 100
rect 36 98 40 102
rect 46 98 50 102
rect 66 98 70 102
rect 530 98 534 102
rect 544 95 548 99
rect 554 95 558 99
rect 582 96 586 100
rect 592 96 596 100
rect 6 86 10 90
rect 66 88 70 92
rect 530 88 534 92
rect 582 86 586 90
rect 592 86 596 90
rect 6 76 10 80
rect 36 78 40 82
rect 46 78 50 82
rect 544 75 548 79
rect 554 75 558 79
rect 582 76 586 80
rect 592 76 596 80
rect 6 66 10 70
rect 36 68 40 72
rect 46 68 50 72
rect 80 69 84 73
rect 109 68 113 72
rect 120 68 124 72
rect 130 68 134 72
rect 140 68 144 72
rect 150 68 154 72
rect 160 68 164 72
rect 170 68 174 72
rect 180 68 184 72
rect 190 68 194 72
rect 200 68 204 72
rect 210 68 214 72
rect 220 68 224 72
rect 230 68 234 72
rect 366 68 370 72
rect 376 68 380 72
rect 386 68 390 72
rect 396 68 400 72
rect 406 68 410 72
rect 416 68 420 72
rect 426 68 430 72
rect 436 68 440 72
rect 446 68 450 72
rect 456 68 460 72
rect 466 68 470 72
rect 476 68 480 72
rect 486 68 490 72
rect 544 65 548 69
rect 554 65 558 69
rect 582 66 586 70
rect 592 66 596 70
rect 6 56 10 60
rect 80 58 84 62
rect 109 58 113 62
rect 130 56 134 60
rect 150 56 154 60
rect 170 56 174 60
rect 190 56 194 60
rect 210 56 214 60
rect 230 56 234 60
rect 366 56 370 60
rect 386 56 390 60
rect 406 56 410 60
rect 426 56 430 60
rect 446 56 450 60
rect 466 56 470 60
rect 486 58 490 62
rect 582 56 586 60
rect 592 56 596 60
rect 36 52 40 56
rect 50 52 54 56
rect 60 52 64 56
rect 70 52 74 56
rect 528 52 532 56
rect 538 52 542 56
rect 554 52 558 56
rect 6 46 10 50
rect 109 48 113 52
rect 130 46 134 50
rect 150 46 154 50
rect 170 46 174 50
rect 190 46 194 50
rect 210 46 214 50
rect 230 46 234 50
rect 366 46 370 50
rect 386 46 390 50
rect 406 46 410 50
rect 426 46 430 50
rect 446 46 450 50
rect 466 46 470 50
rect 486 48 490 52
rect 582 46 586 50
rect 592 46 596 50
rect 6 36 10 40
rect 80 38 84 42
rect 109 38 113 42
rect 130 36 134 40
rect 150 36 154 40
rect 170 36 174 40
rect 190 36 194 40
rect 210 36 214 40
rect 230 36 234 40
rect 366 36 370 40
rect 386 36 390 40
rect 406 36 410 40
rect 426 36 430 40
rect 446 36 450 40
rect 466 36 470 40
rect 486 38 490 42
rect 50 32 54 36
rect 60 32 64 36
rect 70 32 74 36
rect 528 34 532 38
rect 582 36 586 40
rect 592 36 596 40
rect 554 32 558 36
rect 6 26 10 30
rect 582 26 586 30
rect 592 26 596 30
rect 6 16 10 20
rect 582 16 586 20
rect 592 16 596 20
rect 6 6 10 10
rect 16 4 20 8
rect 26 4 30 8
rect 36 4 40 8
rect 48 4 52 8
rect 58 6 62 10
rect 68 6 72 10
rect 78 4 82 8
rect 88 4 92 8
rect 98 4 102 8
rect 108 4 112 8
rect 118 6 122 10
rect 128 6 132 10
rect 138 6 142 10
rect 148 6 152 10
rect 158 6 162 10
rect 168 6 172 10
rect 178 6 182 10
rect 188 6 192 10
rect 198 6 202 10
rect 208 6 212 10
rect 218 6 222 10
rect 228 6 232 10
rect 238 6 242 10
rect 248 6 252 10
rect 258 6 262 10
rect 268 6 272 10
rect 278 6 282 10
rect 288 6 292 10
rect 298 6 302 10
rect 308 6 312 10
rect 318 6 322 10
rect 328 6 332 10
rect 340 6 344 10
rect 350 6 354 10
rect 360 6 364 10
rect 370 6 374 10
rect 380 6 384 10
rect 390 6 394 10
rect 400 6 404 10
rect 410 6 414 10
rect 420 6 424 10
rect 430 6 434 10
rect 440 6 444 10
rect 450 6 454 10
rect 460 6 464 10
rect 470 6 474 10
rect 480 4 484 8
rect 490 4 494 8
rect 500 4 504 8
rect 510 4 514 8
rect 520 4 524 8
rect 530 4 534 8
rect 540 6 544 10
rect 550 6 554 10
rect 560 6 564 10
rect 570 6 574 10
rect 580 6 584 10
rect 592 6 596 10
<< metal1 >>
rect 124 1400 476 1480
rect 204 1380 396 1400
rect 224 1360 376 1380
rect 0 1316 232 1338
rect 0 850 20 1316
rect 28 1234 234 1310
rect 240 1308 360 1360
rect 368 1316 600 1338
rect 28 860 58 1234
rect 64 872 72 1228
rect 78 1184 104 1234
rect 240 1224 286 1308
rect 112 1191 286 1224
rect 78 1104 234 1184
rect 78 1054 104 1104
rect 240 1096 286 1191
rect 111 1061 286 1096
rect 78 976 234 1054
rect 78 924 104 976
rect 240 966 286 1061
rect 111 933 286 966
rect 78 878 232 924
rect 64 860 82 872
rect 88 860 232 878
rect 0 808 58 850
rect 0 708 22 808
rect 0 696 12 708
rect 0 684 44 696
rect 0 652 44 664
rect 0 640 12 652
rect 0 544 22 640
rect 0 16 16 544
rect 34 75 58 486
rect 64 86 72 860
rect 78 820 231 850
rect 78 808 216 820
rect 240 814 286 933
rect 294 860 306 1296
rect 314 1224 360 1308
rect 366 1232 572 1310
rect 314 1191 489 1224
rect 314 1096 360 1191
rect 497 1181 522 1232
rect 366 1104 522 1181
rect 314 1061 489 1096
rect 314 966 360 1061
rect 497 1054 522 1104
rect 366 976 522 1054
rect 314 933 489 966
rect 296 820 304 850
rect 314 814 360 933
rect 497 924 522 976
rect 368 878 522 924
rect 368 860 512 878
rect 528 872 536 1226
rect 518 860 536 872
rect 542 860 572 1232
rect 368 820 520 850
rect 222 786 380 814
rect 240 776 380 786
rect 80 684 230 696
rect 80 652 230 664
rect 240 578 286 776
rect 300 770 380 776
rect 246 532 286 578
rect 316 532 380 770
rect 388 684 522 696
rect 388 672 426 684
rect 388 652 522 664
rect 78 508 228 526
rect 78 506 216 508
rect 78 494 214 506
rect 78 360 100 494
rect 246 492 380 532
rect 386 520 394 536
rect 482 520 490 536
rect 386 494 460 520
rect 480 508 508 520
rect 246 488 352 492
rect 106 420 240 486
rect 246 410 286 488
rect 112 372 286 410
rect 106 360 240 364
rect 78 286 240 360
rect 78 234 106 286
rect 246 278 286 372
rect 112 242 286 278
rect 78 166 240 234
rect 106 158 240 166
rect 246 148 286 242
rect 106 112 286 148
rect 34 32 86 75
rect 106 36 238 104
rect 46 28 80 32
rect 114 28 238 36
rect 246 98 286 112
rect 294 108 306 481
rect 314 411 352 488
rect 359 419 494 486
rect 314 371 494 411
rect 314 278 352 371
rect 360 286 494 365
rect 314 241 494 278
rect 314 148 352 241
rect 360 158 494 234
rect 314 112 494 148
rect 314 98 352 112
rect 246 25 352 98
rect 360 32 494 104
rect 528 86 536 860
rect 580 850 600 1316
rect 544 820 600 850
rect 586 784 600 820
rect 576 776 600 784
rect 578 710 600 776
rect 580 696 600 710
rect 542 684 600 696
rect 542 652 550 664
rect 580 640 600 664
rect 578 522 600 640
rect 546 494 600 522
rect 542 75 572 486
rect 526 32 572 75
rect 360 28 482 32
rect 538 28 572 32
rect 578 16 600 494
rect 0 0 600 16
<< metal2 >>
rect 0 1190 600 1340
rect 0 1180 104 1190
rect 284 1180 316 1190
rect 497 1180 600 1190
rect 0 1040 600 1180
rect 0 1030 104 1040
rect 284 1030 316 1040
rect 500 1030 600 1040
rect 0 880 600 1030
rect 0 878 58 880
rect 90 874 510 880
rect 542 878 600 880
rect 64 866 82 872
rect 518 866 536 872
rect 64 860 536 866
rect 72 858 536 860
rect 20 844 576 850
rect 0 777 600 844
rect 0 767 68 777
rect 123 767 163 777
rect 238 767 280 777
rect 381 767 421 777
rect 500 767 600 777
rect 0 686 600 767
rect 273 683 426 686
rect 484 685 522 686
rect 388 673 426 683
rect 16 662 36 663
rect 62 662 180 663
rect 206 662 230 663
rect 16 652 230 662
rect 273 659 426 665
rect 484 659 522 663
rect 273 652 522 659
rect 0 582 600 652
rect 0 572 36 582
rect 92 572 136 582
rect 188 572 232 582
rect 336 572 379 582
rect 447 572 490 582
rect 561 572 600 582
rect 0 492 600 572
rect 64 474 536 484
rect 64 466 72 474
rect 528 466 536 474
rect 0 456 70 460
rect 108 456 492 466
rect 542 456 600 460
rect 0 310 600 456
rect 0 300 100 310
rect 286 300 314 310
rect 500 300 600 310
rect 0 160 600 300
rect 0 150 100 160
rect 286 150 314 160
rect 500 150 600 160
rect 0 47 600 150
rect 0 38 246 47
rect 0 0 14 38
rect 48 0 80 38
rect 114 0 246 38
rect 256 0 344 39
rect 352 35 600 47
rect 352 0 480 35
rect 540 0 600 35
<< gv1 >>
rect 30 1302 34 1306
rect 40 1302 44 1306
rect 50 1302 54 1306
rect 60 1302 64 1306
rect 70 1302 74 1306
rect 80 1302 84 1306
rect 90 1302 94 1306
rect 100 1302 104 1306
rect 110 1302 114 1306
rect 120 1302 124 1306
rect 130 1302 134 1306
rect 140 1302 144 1306
rect 150 1302 154 1306
rect 160 1302 164 1306
rect 170 1302 174 1306
rect 180 1302 184 1306
rect 190 1302 194 1306
rect 200 1302 204 1306
rect 210 1302 214 1306
rect 220 1302 224 1306
rect 376 1304 380 1308
rect 386 1304 390 1308
rect 396 1304 400 1308
rect 406 1304 410 1308
rect 416 1304 420 1308
rect 426 1304 430 1308
rect 436 1304 440 1308
rect 446 1304 450 1308
rect 456 1304 460 1308
rect 466 1304 470 1308
rect 476 1304 480 1308
rect 486 1304 490 1308
rect 496 1304 500 1308
rect 506 1304 510 1308
rect 516 1304 520 1308
rect 546 1304 550 1308
rect 556 1304 560 1308
rect 566 1304 570 1308
rect 30 1292 34 1296
rect 566 1294 570 1298
rect 30 1282 34 1286
rect 42 1284 46 1288
rect 52 1284 56 1288
rect 62 1284 66 1288
rect 72 1284 76 1288
rect 82 1284 86 1288
rect 124 1284 128 1288
rect 154 1284 158 1288
rect 184 1284 188 1288
rect 214 1284 218 1288
rect 378 1284 382 1288
rect 408 1284 412 1288
rect 438 1284 442 1288
rect 468 1284 472 1288
rect 510 1284 514 1288
rect 544 1284 548 1288
rect 554 1284 558 1288
rect 566 1284 570 1288
rect 298 1278 302 1282
rect 30 1272 34 1276
rect 62 1274 66 1278
rect 72 1274 76 1278
rect 82 1274 86 1278
rect 124 1274 128 1278
rect 154 1274 158 1278
rect 184 1274 188 1278
rect 214 1274 218 1278
rect 378 1274 382 1278
rect 408 1274 412 1278
rect 438 1274 442 1278
rect 468 1274 472 1278
rect 510 1274 514 1278
rect 566 1274 570 1278
rect 30 1262 34 1266
rect 62 1264 66 1268
rect 72 1264 76 1268
rect 82 1264 86 1268
rect 124 1264 128 1268
rect 154 1264 158 1268
rect 184 1264 188 1268
rect 214 1264 218 1268
rect 378 1264 382 1268
rect 408 1264 412 1268
rect 438 1264 442 1268
rect 468 1264 472 1268
rect 510 1264 514 1268
rect 566 1264 570 1268
rect 30 1252 34 1256
rect 566 1254 570 1258
rect 30 1242 34 1246
rect 42 1244 46 1248
rect 52 1244 56 1248
rect 66 1245 70 1249
rect 544 1244 548 1248
rect 554 1244 558 1248
rect 566 1244 570 1248
rect 86 1238 90 1242
rect 96 1238 100 1242
rect 106 1238 110 1242
rect 116 1238 120 1242
rect 126 1238 130 1242
rect 136 1238 140 1242
rect 146 1238 150 1242
rect 156 1238 160 1242
rect 166 1238 170 1242
rect 176 1238 180 1242
rect 186 1238 190 1242
rect 196 1238 200 1242
rect 206 1238 210 1242
rect 216 1238 220 1242
rect 226 1238 230 1242
rect 298 1238 302 1242
rect 370 1238 374 1242
rect 380 1238 384 1242
rect 390 1238 394 1242
rect 400 1238 404 1242
rect 410 1238 414 1242
rect 420 1238 424 1242
rect 430 1238 434 1242
rect 440 1238 444 1242
rect 450 1238 454 1242
rect 460 1238 464 1242
rect 470 1238 474 1242
rect 480 1238 484 1242
rect 490 1238 494 1242
rect 500 1238 504 1242
rect 510 1238 514 1242
rect 30 1232 34 1236
rect 566 1234 570 1238
rect 84 1227 88 1231
rect 94 1227 98 1231
rect 30 1222 34 1226
rect 500 1223 504 1227
rect 510 1223 514 1227
rect 566 1224 570 1228
rect 84 1217 88 1221
rect 94 1217 98 1221
rect 30 1212 34 1216
rect 500 1213 504 1217
rect 510 1213 514 1217
rect 566 1214 570 1218
rect 30 1202 34 1206
rect 42 1204 46 1208
rect 52 1204 56 1208
rect 84 1207 88 1211
rect 94 1207 98 1211
rect 500 1203 504 1207
rect 510 1203 514 1207
rect 544 1204 548 1208
rect 554 1204 558 1208
rect 566 1204 570 1208
rect 84 1197 88 1201
rect 94 1197 98 1201
rect 298 1198 302 1202
rect 30 1192 34 1196
rect 500 1193 504 1197
rect 510 1193 514 1197
rect 566 1194 570 1198
rect 84 1187 88 1191
rect 94 1187 98 1191
rect 30 1182 34 1186
rect 500 1183 504 1187
rect 510 1183 514 1187
rect 566 1184 570 1188
rect 30 1172 34 1176
rect 86 1174 90 1178
rect 96 1174 100 1178
rect 106 1174 110 1178
rect 116 1174 120 1178
rect 126 1174 130 1178
rect 136 1174 140 1178
rect 146 1174 150 1178
rect 156 1174 160 1178
rect 166 1174 170 1178
rect 176 1174 180 1178
rect 186 1174 190 1178
rect 196 1174 200 1178
rect 206 1174 210 1178
rect 216 1174 220 1178
rect 226 1174 230 1178
rect 370 1172 374 1176
rect 380 1172 384 1176
rect 390 1172 394 1176
rect 400 1172 404 1176
rect 410 1172 414 1176
rect 420 1172 424 1176
rect 430 1172 434 1176
rect 440 1172 444 1176
rect 450 1172 454 1176
rect 460 1172 464 1176
rect 470 1172 474 1176
rect 480 1172 484 1176
rect 490 1172 494 1176
rect 500 1172 504 1176
rect 510 1172 514 1176
rect 566 1174 570 1178
rect 30 1162 34 1166
rect 42 1164 46 1168
rect 52 1164 56 1168
rect 544 1164 548 1168
rect 554 1164 558 1168
rect 566 1164 570 1168
rect 298 1158 302 1162
rect 30 1152 34 1156
rect 566 1154 570 1158
rect 85 1146 89 1150
rect 95 1146 99 1150
rect 105 1146 109 1150
rect 115 1146 119 1150
rect 145 1146 149 1150
rect 175 1146 179 1150
rect 205 1146 209 1150
rect 390 1146 394 1150
rect 420 1146 424 1150
rect 450 1146 454 1150
rect 480 1146 484 1150
rect 490 1146 494 1150
rect 500 1146 504 1150
rect 510 1146 514 1150
rect 30 1142 34 1146
rect 566 1144 570 1148
rect 30 1132 34 1136
rect 85 1134 89 1138
rect 95 1134 99 1138
rect 105 1134 109 1138
rect 115 1134 119 1138
rect 145 1134 149 1138
rect 175 1134 179 1138
rect 205 1134 209 1138
rect 390 1134 394 1138
rect 420 1134 424 1138
rect 450 1134 454 1138
rect 480 1134 484 1138
rect 490 1134 494 1138
rect 500 1134 504 1138
rect 510 1134 514 1138
rect 566 1134 570 1138
rect 30 1122 34 1126
rect 42 1124 46 1128
rect 52 1124 56 1128
rect 544 1124 548 1128
rect 554 1124 558 1128
rect 566 1124 570 1128
rect 298 1118 302 1122
rect 30 1112 34 1116
rect 566 1114 570 1118
rect 86 1107 90 1111
rect 96 1107 100 1111
rect 106 1107 110 1111
rect 116 1107 120 1111
rect 126 1107 130 1111
rect 136 1107 140 1111
rect 146 1107 150 1111
rect 156 1107 160 1111
rect 166 1107 170 1111
rect 176 1107 180 1111
rect 186 1107 190 1111
rect 196 1107 200 1111
rect 206 1107 210 1111
rect 216 1107 220 1111
rect 226 1107 230 1111
rect 370 1108 374 1112
rect 380 1108 384 1112
rect 390 1108 394 1112
rect 400 1108 404 1112
rect 410 1108 414 1112
rect 420 1108 424 1112
rect 430 1108 434 1112
rect 440 1108 444 1112
rect 450 1108 454 1112
rect 460 1108 464 1112
rect 470 1108 474 1112
rect 480 1108 484 1112
rect 490 1108 494 1112
rect 500 1108 504 1112
rect 510 1108 514 1112
rect 30 1102 34 1106
rect 566 1104 570 1108
rect 86 1097 90 1101
rect 96 1097 100 1101
rect 500 1097 504 1101
rect 510 1097 514 1101
rect 30 1092 34 1096
rect 566 1094 570 1098
rect 30 1082 34 1086
rect 42 1084 46 1088
rect 52 1084 56 1088
rect 86 1087 90 1091
rect 96 1087 100 1091
rect 500 1087 504 1091
rect 510 1087 514 1091
rect 544 1084 548 1088
rect 554 1084 558 1088
rect 566 1084 570 1088
rect 86 1077 90 1081
rect 96 1077 100 1081
rect 298 1078 302 1082
rect 500 1077 504 1081
rect 510 1077 514 1081
rect 30 1072 34 1076
rect 566 1074 570 1078
rect 86 1067 90 1071
rect 96 1067 100 1071
rect 500 1067 504 1071
rect 510 1067 514 1071
rect 30 1062 34 1066
rect 566 1064 570 1068
rect 86 1057 90 1061
rect 96 1057 100 1061
rect 500 1057 504 1061
rect 510 1057 514 1061
rect 30 1052 34 1056
rect 566 1054 570 1058
rect 30 1042 34 1046
rect 42 1044 46 1048
rect 52 1044 56 1048
rect 86 1046 90 1050
rect 96 1046 100 1050
rect 106 1046 110 1050
rect 116 1046 120 1050
rect 126 1046 130 1050
rect 136 1046 140 1050
rect 146 1046 150 1050
rect 156 1046 160 1050
rect 166 1046 170 1050
rect 176 1046 180 1050
rect 186 1046 190 1050
rect 196 1046 200 1050
rect 206 1046 210 1050
rect 216 1046 220 1050
rect 226 1046 230 1050
rect 370 1046 374 1050
rect 380 1046 384 1050
rect 390 1046 394 1050
rect 400 1046 404 1050
rect 410 1046 414 1050
rect 420 1046 424 1050
rect 430 1046 434 1050
rect 440 1046 444 1050
rect 450 1046 454 1050
rect 460 1046 464 1050
rect 470 1046 474 1050
rect 480 1046 484 1050
rect 490 1046 494 1050
rect 500 1046 504 1050
rect 510 1046 514 1050
rect 544 1044 548 1048
rect 554 1044 558 1048
rect 566 1044 570 1048
rect 298 1038 302 1042
rect 30 1032 34 1036
rect 566 1034 570 1038
rect 30 1022 34 1026
rect 566 1024 570 1028
rect 84 1018 88 1022
rect 94 1018 98 1022
rect 104 1018 108 1022
rect 114 1018 118 1022
rect 144 1018 148 1022
rect 174 1018 178 1022
rect 204 1018 208 1022
rect 389 1018 393 1022
rect 419 1018 423 1022
rect 449 1018 453 1022
rect 479 1018 483 1022
rect 489 1018 493 1022
rect 499 1018 503 1022
rect 509 1018 513 1022
rect 30 1012 34 1016
rect 566 1014 570 1018
rect 30 1002 34 1006
rect 42 1004 46 1008
rect 52 1004 56 1008
rect 84 1006 88 1010
rect 94 1006 98 1010
rect 104 1006 108 1010
rect 114 1006 118 1010
rect 144 1006 148 1010
rect 174 1006 178 1010
rect 204 1006 208 1010
rect 389 1006 393 1010
rect 419 1006 423 1010
rect 449 1006 453 1010
rect 479 1006 483 1010
rect 489 1006 493 1010
rect 499 1006 503 1010
rect 509 1006 513 1010
rect 544 1004 548 1008
rect 554 1004 558 1008
rect 566 1004 570 1008
rect 298 998 302 1002
rect 30 992 34 996
rect 566 994 570 998
rect 30 982 34 986
rect 566 984 570 988
rect 86 980 90 984
rect 96 980 100 984
rect 106 980 110 984
rect 116 980 120 984
rect 126 980 130 984
rect 136 980 140 984
rect 146 980 150 984
rect 156 980 160 984
rect 166 980 170 984
rect 176 980 180 984
rect 186 980 190 984
rect 196 980 200 984
rect 206 980 210 984
rect 216 980 220 984
rect 226 980 230 984
rect 370 980 374 984
rect 380 980 384 984
rect 390 980 394 984
rect 400 980 404 984
rect 410 980 414 984
rect 420 980 424 984
rect 430 980 434 984
rect 440 980 444 984
rect 450 980 454 984
rect 460 980 464 984
rect 470 980 474 984
rect 480 980 484 984
rect 490 980 494 984
rect 500 980 504 984
rect 510 980 514 984
rect 30 972 34 976
rect 566 974 570 978
rect 86 969 90 973
rect 96 969 100 973
rect 502 968 506 972
rect 512 968 516 972
rect 30 962 34 966
rect 42 964 46 968
rect 52 964 56 968
rect 544 964 548 968
rect 554 964 558 968
rect 566 964 570 968
rect 86 959 90 963
rect 96 959 100 963
rect 298 958 302 962
rect 502 958 506 962
rect 512 958 516 962
rect 30 952 34 956
rect 566 954 570 958
rect 86 949 90 953
rect 96 949 100 953
rect 502 948 506 952
rect 512 948 516 952
rect 30 942 34 946
rect 566 944 570 948
rect 86 939 90 943
rect 96 939 100 943
rect 502 938 506 942
rect 512 938 516 942
rect 30 932 34 936
rect 566 934 570 938
rect 86 929 90 933
rect 96 929 100 933
rect 502 928 506 932
rect 512 928 516 932
rect 30 922 34 926
rect 42 924 46 928
rect 52 924 56 928
rect 544 924 548 928
rect 554 924 558 928
rect 566 924 570 928
rect 84 916 88 920
rect 94 916 98 920
rect 104 916 108 920
rect 114 916 118 920
rect 124 916 128 920
rect 134 916 138 920
rect 144 916 148 920
rect 154 916 158 920
rect 164 916 168 920
rect 174 916 178 920
rect 184 916 188 920
rect 194 916 198 920
rect 204 916 208 920
rect 214 916 218 920
rect 224 916 228 920
rect 298 918 302 922
rect 372 916 376 920
rect 382 916 386 920
rect 392 916 396 920
rect 402 916 406 920
rect 412 916 416 920
rect 422 916 426 920
rect 432 916 436 920
rect 442 916 446 920
rect 452 916 456 920
rect 462 916 466 920
rect 472 916 476 920
rect 482 916 486 920
rect 492 916 496 920
rect 502 916 506 920
rect 512 916 516 920
rect 30 912 34 916
rect 566 914 570 918
rect 30 902 34 906
rect 566 904 570 908
rect 30 892 34 896
rect 566 894 570 898
rect 82 888 86 892
rect 93 888 97 892
rect 104 888 108 892
rect 115 888 119 892
rect 145 888 149 892
rect 175 888 179 892
rect 205 888 209 892
rect 391 888 395 892
rect 421 888 425 892
rect 451 888 455 892
rect 481 888 485 892
rect 492 888 496 892
rect 503 888 507 892
rect 514 888 518 892
rect 30 882 34 886
rect 42 884 46 888
rect 52 884 56 888
rect 544 884 548 888
rect 554 884 558 888
rect 566 884 570 888
rect 95 876 99 880
rect 115 876 119 880
rect 145 876 149 880
rect 175 876 179 880
rect 205 876 209 880
rect 298 878 302 882
rect 391 876 395 880
rect 421 876 425 880
rect 451 876 455 880
rect 481 876 485 880
rect 501 876 505 880
rect 66 864 70 868
rect 76 864 80 868
rect 520 864 524 868
rect 530 864 534 868
rect 32 844 36 848
rect 42 844 46 848
rect 52 844 56 848
rect 80 844 84 848
rect 90 844 94 848
rect 100 844 104 848
rect 110 844 114 848
rect 120 844 124 848
rect 130 844 134 848
rect 140 844 144 848
rect 150 844 154 848
rect 160 844 164 848
rect 170 844 174 848
rect 180 844 184 848
rect 190 844 194 848
rect 200 844 204 848
rect 210 844 214 848
rect 220 844 224 848
rect 298 844 302 848
rect 370 844 374 848
rect 380 844 384 848
rect 390 844 394 848
rect 400 844 404 848
rect 410 844 414 848
rect 420 844 424 848
rect 430 844 434 848
rect 440 844 444 848
rect 450 844 454 848
rect 460 844 464 848
rect 470 844 474 848
rect 480 844 484 848
rect 490 844 494 848
rect 500 844 504 848
rect 510 844 514 848
rect 550 844 554 848
rect 560 844 564 848
rect 570 844 574 848
rect 592 817 596 821
rect 16 812 20 816
rect 28 812 32 816
rect 38 812 42 816
rect 48 812 52 816
rect 80 812 84 816
rect 90 812 94 816
rect 100 812 104 816
rect 110 812 114 816
rect 120 812 124 816
rect 130 812 134 816
rect 140 812 144 816
rect 150 812 154 816
rect 160 812 164 816
rect 170 812 174 816
rect 180 812 184 816
rect 190 812 194 816
rect 200 812 204 816
rect 210 812 214 816
rect 16 802 20 806
rect 592 797 596 801
rect 16 792 20 796
rect 16 780 20 784
rect 578 778 582 782
rect 592 777 596 781
rect 16 770 20 774
rect 16 760 20 764
rect 592 757 596 761
rect 16 750 20 754
rect 580 745 584 749
rect 16 740 20 744
rect 592 737 596 741
rect 16 730 20 734
rect 580 725 584 729
rect 16 720 20 724
rect 592 717 596 721
rect 16 710 20 714
rect 582 699 586 703
rect 592 697 596 701
rect 208 689 212 693
rect 506 687 510 691
rect 390 675 394 679
rect 400 675 404 679
rect 410 675 414 679
rect 420 675 424 679
rect 140 657 144 661
rect 210 657 214 661
rect 410 657 414 661
rect 506 657 510 661
rect 4 636 8 640
rect 592 638 596 642
rect 16 630 20 634
rect 16 620 20 624
rect 4 616 8 620
rect 580 617 584 621
rect 592 618 596 622
rect 16 610 20 614
rect 16 600 20 604
rect 4 596 8 600
rect 580 597 584 601
rect 592 598 596 602
rect 16 590 20 594
rect 16 580 20 584
rect 4 576 8 580
rect 580 577 584 581
rect 592 578 596 582
rect 16 570 20 574
rect 16 560 20 564
rect 4 556 8 560
rect 580 557 584 561
rect 592 558 596 562
rect 16 550 20 554
rect 4 536 8 540
rect 582 535 586 539
rect 592 538 596 542
rect 4 516 8 520
rect 592 518 596 522
rect 108 496 112 500
rect 118 496 122 500
rect 128 496 132 500
rect 138 496 142 500
rect 148 496 152 500
rect 158 496 162 500
rect 168 496 172 500
rect 178 496 182 500
rect 188 496 192 500
rect 198 496 202 500
rect 208 496 212 500
rect 391 496 395 500
rect 401 496 405 500
rect 411 496 415 500
rect 421 496 425 500
rect 431 496 435 500
rect 441 496 445 500
rect 451 496 455 500
rect 549 496 553 500
rect 559 496 563 500
rect 569 496 573 500
rect 66 478 70 482
rect 530 478 534 482
rect 66 468 70 472
rect 530 468 534 472
rect 130 460 134 464
rect 160 460 164 464
rect 190 460 194 464
rect 220 460 224 464
rect 386 460 390 464
rect 416 460 420 464
rect 446 460 450 464
rect 476 460 480 464
rect 298 452 302 456
rect 566 453 570 457
rect 36 448 40 452
rect 46 448 50 452
rect 130 448 134 452
rect 160 448 164 452
rect 190 448 194 452
rect 220 448 224 452
rect 386 448 390 452
rect 416 448 420 452
rect 446 448 450 452
rect 476 448 480 452
rect 544 445 548 449
rect 554 445 558 449
rect 566 443 570 447
rect 566 433 570 437
rect 110 423 114 427
rect 120 423 124 427
rect 130 423 134 427
rect 140 423 144 427
rect 150 423 154 427
rect 160 423 164 427
rect 170 423 174 427
rect 180 423 184 427
rect 190 423 194 427
rect 200 423 204 427
rect 210 423 214 427
rect 220 423 224 427
rect 230 423 234 427
rect 298 422 302 426
rect 366 423 370 427
rect 376 423 380 427
rect 386 423 390 427
rect 396 423 400 427
rect 406 423 410 427
rect 416 423 420 427
rect 426 423 430 427
rect 436 423 440 427
rect 446 423 450 427
rect 456 423 460 427
rect 466 423 470 427
rect 476 423 480 427
rect 486 423 490 427
rect 566 423 570 427
rect 566 413 570 417
rect 36 408 40 412
rect 46 408 50 412
rect 544 405 548 409
rect 554 405 558 409
rect 566 403 570 407
rect 298 392 302 396
rect 566 393 570 397
rect 566 383 570 387
rect 566 373 570 377
rect 36 368 40 372
rect 46 368 50 372
rect 298 362 302 366
rect 544 365 548 369
rect 554 365 558 369
rect 566 363 570 367
rect 114 356 118 360
rect 124 356 128 360
rect 134 356 138 360
rect 144 356 148 360
rect 154 356 158 360
rect 164 356 168 360
rect 174 356 178 360
rect 184 356 188 360
rect 194 356 198 360
rect 204 356 208 360
rect 214 356 218 360
rect 224 356 228 360
rect 234 356 238 360
rect 366 356 370 360
rect 376 356 380 360
rect 386 356 390 360
rect 396 356 400 360
rect 406 356 410 360
rect 416 356 420 360
rect 426 356 430 360
rect 436 356 440 360
rect 446 356 450 360
rect 456 356 460 360
rect 466 356 470 360
rect 476 356 480 360
rect 486 356 490 360
rect 566 353 570 357
rect 566 343 570 347
rect 298 332 302 336
rect 566 333 570 337
rect 36 328 40 332
rect 46 328 50 332
rect 132 328 136 332
rect 162 328 166 332
rect 192 328 196 332
rect 222 328 226 332
rect 385 329 389 333
rect 415 329 419 333
rect 445 329 449 333
rect 475 329 479 333
rect 544 325 548 329
rect 554 325 558 329
rect 566 323 570 327
rect 132 316 136 320
rect 162 316 166 320
rect 192 316 196 320
rect 222 316 226 320
rect 385 317 389 321
rect 415 317 419 321
rect 445 317 449 321
rect 475 317 479 321
rect 566 313 570 317
rect 298 302 302 306
rect 566 303 570 307
rect 36 288 40 292
rect 46 288 50 292
rect 112 290 116 294
rect 122 290 126 294
rect 132 290 136 294
rect 142 290 146 294
rect 152 290 156 294
rect 162 290 166 294
rect 172 290 176 294
rect 182 290 186 294
rect 192 290 196 294
rect 202 290 206 294
rect 212 290 216 294
rect 222 290 226 294
rect 232 290 236 294
rect 365 290 369 294
rect 375 290 379 294
rect 385 290 389 294
rect 395 290 399 294
rect 405 290 409 294
rect 415 290 419 294
rect 425 290 429 294
rect 435 290 439 294
rect 445 290 449 294
rect 455 290 459 294
rect 465 290 469 294
rect 475 290 479 294
rect 485 290 489 294
rect 566 293 570 297
rect 544 285 548 289
rect 554 285 558 289
rect 566 283 570 287
rect 298 272 302 276
rect 566 273 570 277
rect 566 263 570 267
rect 566 253 570 257
rect 36 248 40 252
rect 46 248 50 252
rect 298 242 302 246
rect 544 245 548 249
rect 554 245 558 249
rect 566 243 570 247
rect 566 233 570 237
rect 112 226 116 230
rect 122 226 126 230
rect 132 226 136 230
rect 142 226 146 230
rect 152 226 156 230
rect 162 226 166 230
rect 172 226 176 230
rect 182 226 186 230
rect 192 226 196 230
rect 202 226 206 230
rect 212 226 216 230
rect 222 226 226 230
rect 232 226 236 230
rect 366 225 370 229
rect 376 225 380 229
rect 386 225 390 229
rect 396 225 400 229
rect 406 225 410 229
rect 416 225 420 229
rect 426 225 430 229
rect 436 225 440 229
rect 446 225 450 229
rect 456 225 460 229
rect 466 225 470 229
rect 476 225 480 229
rect 486 225 490 229
rect 566 223 570 227
rect 298 212 302 216
rect 566 213 570 217
rect 36 208 40 212
rect 46 208 50 212
rect 544 205 548 209
rect 554 205 558 209
rect 566 203 570 207
rect 131 198 135 202
rect 161 198 165 202
rect 191 198 195 202
rect 221 198 225 202
rect 386 198 390 202
rect 416 198 420 202
rect 446 198 450 202
rect 476 198 480 202
rect 566 193 570 197
rect 131 186 135 190
rect 161 186 165 190
rect 191 186 195 190
rect 221 186 225 190
rect 386 186 390 190
rect 416 186 420 190
rect 446 186 450 190
rect 476 186 480 190
rect 298 182 302 186
rect 566 183 570 187
rect 566 173 570 177
rect 36 168 40 172
rect 46 168 50 172
rect 112 162 116 166
rect 122 162 126 166
rect 132 162 136 166
rect 142 162 146 166
rect 152 162 156 166
rect 162 162 166 166
rect 172 162 176 166
rect 182 162 186 166
rect 192 162 196 166
rect 202 162 206 166
rect 212 162 216 166
rect 222 162 226 166
rect 232 162 236 166
rect 366 162 370 166
rect 376 162 380 166
rect 386 162 390 166
rect 396 162 400 166
rect 406 162 410 166
rect 416 162 420 166
rect 426 162 430 166
rect 436 162 440 166
rect 446 162 450 166
rect 456 162 460 166
rect 466 162 470 166
rect 476 162 480 166
rect 486 162 490 166
rect 544 165 548 169
rect 554 165 558 169
rect 566 163 570 167
rect 298 152 302 156
rect 566 153 570 157
rect 566 143 570 147
rect 566 133 570 137
rect 36 128 40 132
rect 46 128 50 132
rect 298 122 302 126
rect 544 125 548 129
rect 554 125 558 129
rect 566 123 570 127
rect 566 113 570 117
rect 566 103 570 107
rect 110 96 114 100
rect 120 96 124 100
rect 130 96 134 100
rect 140 96 144 100
rect 150 96 154 100
rect 160 96 164 100
rect 170 96 174 100
rect 180 96 184 100
rect 190 96 194 100
rect 200 96 204 100
rect 210 96 214 100
rect 220 96 224 100
rect 230 96 234 100
rect 366 97 370 101
rect 376 97 380 101
rect 386 97 390 101
rect 396 97 400 101
rect 406 97 410 101
rect 416 97 420 101
rect 426 97 430 101
rect 436 97 440 101
rect 446 97 450 101
rect 456 97 460 101
rect 466 97 470 101
rect 476 97 480 101
rect 486 97 490 101
rect 566 93 570 97
rect 36 88 40 92
rect 46 88 50 92
rect 544 85 548 89
rect 554 85 558 89
rect 566 83 570 87
rect 566 73 570 77
rect 66 66 70 70
rect 530 67 534 71
rect 566 63 570 67
rect 120 56 124 60
rect 140 56 144 60
rect 160 56 164 60
rect 180 56 184 60
rect 200 56 204 60
rect 220 56 224 60
rect 376 56 380 60
rect 396 56 400 60
rect 416 56 420 60
rect 436 56 440 60
rect 456 56 460 60
rect 476 58 480 62
rect 566 53 570 57
rect 80 48 84 52
rect 120 46 124 50
rect 140 46 144 50
rect 160 46 164 50
rect 180 46 184 50
rect 200 46 204 50
rect 220 46 224 50
rect 376 46 380 50
rect 396 46 400 50
rect 416 46 420 50
rect 436 46 440 50
rect 456 46 460 50
rect 476 48 480 52
rect 36 42 40 46
rect 50 42 54 46
rect 60 42 64 46
rect 70 42 74 46
rect 538 42 542 46
rect 554 42 558 46
rect 566 43 570 47
rect 120 36 124 40
rect 140 36 144 40
rect 160 36 164 40
rect 180 36 184 40
rect 200 36 204 40
rect 220 36 224 40
rect 376 36 380 40
rect 396 36 400 40
rect 416 36 420 40
rect 436 36 440 40
rect 456 36 460 40
rect 476 38 480 42
rect 258 32 262 36
rect 268 32 272 36
rect 278 32 282 36
rect 288 32 292 36
rect 298 32 302 36
rect 308 32 312 36
rect 318 32 322 36
rect 328 32 332 36
rect 338 32 342 36
rect 566 33 570 37
<< labels >>
rlabel metal2 s 4 882 4 882 2 vdd
rlabel metal2 s 4 690 4 690 2 vss
rlabel metal2 s 2 494 2 494 2 vdd
rlabel metal2 s 2 2 2 2 2 vss
rlabel metal2 s 288 18 288 18 2 PAD
rlabel metal1 278 1352 278 1352 2 PAD
rlabel nwell s -4 -4 -4 -4 2 vdd
<< end >>
