module fill1 ();
endmodule
