magic
tech amic5n
timestamp 1623372921
<< nwell >>
rect -130 550 880 1495
<< ntransistor >>
rect 225 95 285 400
rect 465 95 525 400
<< ptransistor >>
rect 225 700 285 1345
rect 465 700 525 1345
<< nselect >>
rect -10 0 760 430
<< pselect >>
rect -10 670 760 1440
<< ndiffusion >>
rect 105 370 225 400
rect 105 320 135 370
rect 185 320 225 370
rect 105 175 225 320
rect 105 125 135 175
rect 185 125 225 175
rect 105 95 225 125
rect 285 95 465 400
rect 525 345 645 400
rect 525 295 565 345
rect 615 295 645 345
rect 525 175 645 295
rect 525 125 565 175
rect 615 125 645 175
rect 525 95 645 125
<< pdiffusion >>
rect 105 1315 225 1345
rect 105 1265 135 1315
rect 185 1265 225 1315
rect 105 1215 225 1265
rect 105 1165 135 1215
rect 185 1165 225 1215
rect 105 1115 225 1165
rect 105 1065 135 1115
rect 185 1065 225 1115
rect 105 1015 225 1065
rect 105 965 135 1015
rect 185 965 225 1015
rect 105 915 225 965
rect 105 865 135 915
rect 185 865 225 915
rect 105 700 225 865
rect 285 1315 465 1345
rect 285 1265 350 1315
rect 400 1265 465 1315
rect 285 1180 465 1265
rect 285 1130 350 1180
rect 400 1130 465 1180
rect 285 1080 465 1130
rect 285 1030 350 1080
rect 400 1030 465 1080
rect 285 980 465 1030
rect 285 930 350 980
rect 400 930 465 980
rect 285 880 465 930
rect 285 830 350 880
rect 400 830 465 880
rect 285 780 465 830
rect 285 730 350 780
rect 400 730 465 780
rect 285 700 465 730
rect 525 1315 645 1345
rect 525 1265 565 1315
rect 615 1265 645 1315
rect 525 1215 645 1265
rect 525 1165 565 1215
rect 615 1165 645 1215
rect 525 1115 645 1165
rect 525 1065 565 1115
rect 615 1065 645 1115
rect 525 1015 645 1065
rect 525 965 565 1015
rect 615 965 645 1015
rect 525 915 645 965
rect 525 865 565 915
rect 615 865 645 915
rect 525 815 645 865
rect 525 765 565 815
rect 615 765 645 815
rect 525 700 645 765
<< ndcontact >>
rect 135 320 185 370
rect 135 125 185 175
rect 565 295 615 345
rect 565 125 615 175
<< pdcontact >>
rect 135 1265 185 1315
rect 135 1165 185 1215
rect 135 1065 185 1115
rect 135 965 185 1015
rect 135 865 185 915
rect 350 1265 400 1315
rect 350 1130 400 1180
rect 350 1030 400 1080
rect 350 930 400 980
rect 350 830 400 880
rect 350 730 400 780
rect 565 1265 615 1315
rect 565 1165 615 1215
rect 565 1065 615 1115
rect 565 965 615 1015
rect 565 865 615 915
rect 565 765 615 815
<< polysilicon >>
rect 225 1345 285 1410
rect 465 1345 525 1410
rect 225 630 285 700
rect 115 610 285 630
rect 115 560 135 610
rect 185 560 285 610
rect 115 540 285 560
rect 225 400 285 540
rect 465 525 525 700
rect 465 505 635 525
rect 465 455 565 505
rect 615 455 635 505
rect 465 435 635 455
rect 465 400 525 435
rect 225 30 285 95
rect 465 30 525 95
<< polycontact >>
rect 135 560 185 610
rect 565 455 615 505
<< metal1 >>
rect 0 1395 750 1485
rect 115 1315 205 1395
rect 115 1265 135 1315
rect 185 1265 205 1315
rect 115 1215 205 1265
rect 115 1165 135 1215
rect 185 1165 205 1215
rect 115 1115 205 1165
rect 115 1065 135 1115
rect 185 1065 205 1115
rect 115 1015 205 1065
rect 115 965 135 1015
rect 185 965 205 1015
rect 115 915 205 965
rect 115 865 135 915
rect 185 865 205 915
rect 115 760 205 865
rect 330 1315 420 1335
rect 330 1265 350 1315
rect 400 1265 420 1315
rect 330 1180 420 1265
rect 330 1130 350 1180
rect 400 1130 420 1180
rect 330 1080 420 1130
rect 330 1030 350 1080
rect 400 1030 420 1080
rect 330 980 420 1030
rect 330 930 350 980
rect 400 930 420 980
rect 330 880 420 930
rect 330 830 350 880
rect 400 830 420 880
rect 330 780 420 830
rect 330 730 350 780
rect 400 730 420 780
rect 545 1315 635 1395
rect 545 1265 565 1315
rect 615 1265 635 1315
rect 545 1215 635 1265
rect 545 1165 565 1215
rect 615 1165 635 1215
rect 545 1115 635 1165
rect 545 1065 565 1115
rect 615 1065 635 1115
rect 545 1015 635 1065
rect 545 965 565 1015
rect 615 965 635 1015
rect 545 915 635 965
rect 545 865 565 915
rect 615 865 635 915
rect 545 815 635 865
rect 545 765 565 815
rect 615 765 635 815
rect 545 745 635 765
rect 115 610 205 685
rect 115 560 135 610
rect 185 560 205 610
rect 115 540 205 560
rect 115 370 205 390
rect 115 320 135 370
rect 185 320 205 370
rect 115 175 205 320
rect 330 365 420 730
rect 545 505 720 525
rect 545 455 565 505
rect 615 455 720 505
rect 545 435 720 455
rect 330 345 635 365
rect 330 295 565 345
rect 615 295 635 345
rect 330 275 635 295
rect 115 125 135 175
rect 185 125 205 175
rect 115 45 205 125
rect 545 175 635 275
rect 545 125 565 175
rect 615 125 635 175
rect 545 45 635 125
rect 0 -45 750 45
<< labels >>
flabel metal1 s 105 -25 105 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel metal1 s 135 550 135 550 2 FreeSans 400 0 0 0 a
port 7 ne
flabel nwell 0 585 0 585 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 360 470 360 470 2 FreeSans 400 0 0 0 z
port 20 ne
flabel metal1 s 616 445 616 445 2 FreeSans 400 0 0 0 b
port 7 ne
<< end >>
