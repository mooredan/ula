magic
tech scmos
timestamp 1591469683
<< metal1 >>
rect -10 -10 260 260
<< metal2 >>
rect -8 -8 258 258
<< gv1 >>
rect 4 244 6 246
rect 14 244 16 246
rect 24 244 26 246
rect 34 244 36 246
rect 44 244 46 246
rect 54 244 56 246
rect 64 244 66 246
rect 74 244 76 246
rect 84 244 86 246
rect 94 244 96 246
rect 104 244 106 246
rect 114 244 116 246
rect 124 244 126 246
rect 134 244 136 246
rect 144 244 146 246
rect 154 244 156 246
rect 164 244 166 246
rect 174 244 176 246
rect 184 244 186 246
rect 194 244 196 246
rect 204 244 206 246
rect 214 244 216 246
rect 224 244 226 246
rect 234 244 236 246
rect 244 244 246 246
rect 4 234 6 236
rect 14 234 16 236
rect 24 234 26 236
rect 34 234 36 236
rect 44 234 46 236
rect 54 234 56 236
rect 64 234 66 236
rect 74 234 76 236
rect 84 234 86 236
rect 94 234 96 236
rect 104 234 106 236
rect 114 234 116 236
rect 124 234 126 236
rect 134 234 136 236
rect 144 234 146 236
rect 154 234 156 236
rect 164 234 166 236
rect 174 234 176 236
rect 184 234 186 236
rect 194 234 196 236
rect 204 234 206 236
rect 214 234 216 236
rect 224 234 226 236
rect 234 234 236 236
rect 244 234 246 236
rect 4 224 6 226
rect 14 224 16 226
rect 24 224 26 226
rect 34 224 36 226
rect 44 224 46 226
rect 54 224 56 226
rect 64 224 66 226
rect 74 224 76 226
rect 84 224 86 226
rect 94 224 96 226
rect 104 224 106 226
rect 114 224 116 226
rect 124 224 126 226
rect 134 224 136 226
rect 144 224 146 226
rect 154 224 156 226
rect 164 224 166 226
rect 174 224 176 226
rect 184 224 186 226
rect 194 224 196 226
rect 204 224 206 226
rect 214 224 216 226
rect 224 224 226 226
rect 234 224 236 226
rect 244 224 246 226
rect 4 214 6 216
rect 14 214 16 216
rect 24 214 26 216
rect 34 214 36 216
rect 44 214 46 216
rect 54 214 56 216
rect 64 214 66 216
rect 74 214 76 216
rect 84 214 86 216
rect 94 214 96 216
rect 104 214 106 216
rect 114 214 116 216
rect 124 214 126 216
rect 134 214 136 216
rect 144 214 146 216
rect 154 214 156 216
rect 164 214 166 216
rect 174 214 176 216
rect 184 214 186 216
rect 194 214 196 216
rect 204 214 206 216
rect 214 214 216 216
rect 224 214 226 216
rect 234 214 236 216
rect 244 214 246 216
rect 4 204 6 206
rect 14 204 16 206
rect 24 204 26 206
rect 34 204 36 206
rect 44 204 46 206
rect 54 204 56 206
rect 64 204 66 206
rect 74 204 76 206
rect 84 204 86 206
rect 94 204 96 206
rect 104 204 106 206
rect 114 204 116 206
rect 124 204 126 206
rect 134 204 136 206
rect 144 204 146 206
rect 154 204 156 206
rect 164 204 166 206
rect 174 204 176 206
rect 184 204 186 206
rect 194 204 196 206
rect 204 204 206 206
rect 214 204 216 206
rect 224 204 226 206
rect 234 204 236 206
rect 244 204 246 206
rect 4 194 6 196
rect 14 194 16 196
rect 24 194 26 196
rect 34 194 36 196
rect 44 194 46 196
rect 54 194 56 196
rect 64 194 66 196
rect 74 194 76 196
rect 84 194 86 196
rect 94 194 96 196
rect 104 194 106 196
rect 114 194 116 196
rect 124 194 126 196
rect 134 194 136 196
rect 144 194 146 196
rect 154 194 156 196
rect 164 194 166 196
rect 174 194 176 196
rect 184 194 186 196
rect 194 194 196 196
rect 204 194 206 196
rect 214 194 216 196
rect 224 194 226 196
rect 234 194 236 196
rect 244 194 246 196
rect 4 184 6 186
rect 14 184 16 186
rect 24 184 26 186
rect 34 184 36 186
rect 44 184 46 186
rect 54 184 56 186
rect 64 184 66 186
rect 74 184 76 186
rect 84 184 86 186
rect 94 184 96 186
rect 104 184 106 186
rect 114 184 116 186
rect 124 184 126 186
rect 134 184 136 186
rect 144 184 146 186
rect 154 184 156 186
rect 164 184 166 186
rect 174 184 176 186
rect 184 184 186 186
rect 194 184 196 186
rect 204 184 206 186
rect 214 184 216 186
rect 224 184 226 186
rect 234 184 236 186
rect 244 184 246 186
rect 4 174 6 176
rect 14 174 16 176
rect 24 174 26 176
rect 34 174 36 176
rect 44 174 46 176
rect 54 174 56 176
rect 64 174 66 176
rect 74 174 76 176
rect 84 174 86 176
rect 94 174 96 176
rect 104 174 106 176
rect 114 174 116 176
rect 124 174 126 176
rect 134 174 136 176
rect 144 174 146 176
rect 154 174 156 176
rect 164 174 166 176
rect 174 174 176 176
rect 184 174 186 176
rect 194 174 196 176
rect 204 174 206 176
rect 214 174 216 176
rect 224 174 226 176
rect 234 174 236 176
rect 244 174 246 176
rect 4 164 6 166
rect 14 164 16 166
rect 24 164 26 166
rect 34 164 36 166
rect 44 164 46 166
rect 54 164 56 166
rect 64 164 66 166
rect 74 164 76 166
rect 84 164 86 166
rect 94 164 96 166
rect 104 164 106 166
rect 114 164 116 166
rect 124 164 126 166
rect 134 164 136 166
rect 144 164 146 166
rect 154 164 156 166
rect 164 164 166 166
rect 174 164 176 166
rect 184 164 186 166
rect 194 164 196 166
rect 204 164 206 166
rect 214 164 216 166
rect 224 164 226 166
rect 234 164 236 166
rect 244 164 246 166
rect 4 154 6 156
rect 14 154 16 156
rect 24 154 26 156
rect 34 154 36 156
rect 44 154 46 156
rect 54 154 56 156
rect 64 154 66 156
rect 74 154 76 156
rect 84 154 86 156
rect 94 154 96 156
rect 104 154 106 156
rect 114 154 116 156
rect 124 154 126 156
rect 134 154 136 156
rect 144 154 146 156
rect 154 154 156 156
rect 164 154 166 156
rect 174 154 176 156
rect 184 154 186 156
rect 194 154 196 156
rect 204 154 206 156
rect 214 154 216 156
rect 224 154 226 156
rect 234 154 236 156
rect 244 154 246 156
rect 4 144 6 146
rect 14 144 16 146
rect 24 144 26 146
rect 34 144 36 146
rect 44 144 46 146
rect 54 144 56 146
rect 64 144 66 146
rect 74 144 76 146
rect 84 144 86 146
rect 94 144 96 146
rect 104 144 106 146
rect 114 144 116 146
rect 124 144 126 146
rect 134 144 136 146
rect 144 144 146 146
rect 154 144 156 146
rect 164 144 166 146
rect 174 144 176 146
rect 184 144 186 146
rect 194 144 196 146
rect 204 144 206 146
rect 214 144 216 146
rect 224 144 226 146
rect 234 144 236 146
rect 244 144 246 146
rect 4 134 6 136
rect 14 134 16 136
rect 24 134 26 136
rect 34 134 36 136
rect 44 134 46 136
rect 54 134 56 136
rect 64 134 66 136
rect 74 134 76 136
rect 84 134 86 136
rect 94 134 96 136
rect 104 134 106 136
rect 114 134 116 136
rect 124 134 126 136
rect 134 134 136 136
rect 144 134 146 136
rect 154 134 156 136
rect 164 134 166 136
rect 174 134 176 136
rect 184 134 186 136
rect 194 134 196 136
rect 204 134 206 136
rect 214 134 216 136
rect 224 134 226 136
rect 234 134 236 136
rect 244 134 246 136
rect 4 124 6 126
rect 14 124 16 126
rect 24 124 26 126
rect 34 124 36 126
rect 44 124 46 126
rect 54 124 56 126
rect 64 124 66 126
rect 74 124 76 126
rect 84 124 86 126
rect 94 124 96 126
rect 104 124 106 126
rect 114 124 116 126
rect 124 124 126 126
rect 134 124 136 126
rect 144 124 146 126
rect 154 124 156 126
rect 164 124 166 126
rect 174 124 176 126
rect 184 124 186 126
rect 194 124 196 126
rect 204 124 206 126
rect 214 124 216 126
rect 224 124 226 126
rect 234 124 236 126
rect 244 124 246 126
rect 4 114 6 116
rect 14 114 16 116
rect 24 114 26 116
rect 34 114 36 116
rect 44 114 46 116
rect 54 114 56 116
rect 64 114 66 116
rect 74 114 76 116
rect 84 114 86 116
rect 94 114 96 116
rect 104 114 106 116
rect 114 114 116 116
rect 124 114 126 116
rect 134 114 136 116
rect 144 114 146 116
rect 154 114 156 116
rect 164 114 166 116
rect 174 114 176 116
rect 184 114 186 116
rect 194 114 196 116
rect 204 114 206 116
rect 214 114 216 116
rect 224 114 226 116
rect 234 114 236 116
rect 244 114 246 116
rect 4 104 6 106
rect 14 104 16 106
rect 24 104 26 106
rect 34 104 36 106
rect 44 104 46 106
rect 54 104 56 106
rect 64 104 66 106
rect 74 104 76 106
rect 84 104 86 106
rect 94 104 96 106
rect 104 104 106 106
rect 114 104 116 106
rect 124 104 126 106
rect 134 104 136 106
rect 144 104 146 106
rect 154 104 156 106
rect 164 104 166 106
rect 174 104 176 106
rect 184 104 186 106
rect 194 104 196 106
rect 204 104 206 106
rect 214 104 216 106
rect 224 104 226 106
rect 234 104 236 106
rect 244 104 246 106
rect 4 94 6 96
rect 14 94 16 96
rect 24 94 26 96
rect 34 94 36 96
rect 44 94 46 96
rect 54 94 56 96
rect 64 94 66 96
rect 74 94 76 96
rect 84 94 86 96
rect 94 94 96 96
rect 104 94 106 96
rect 114 94 116 96
rect 124 94 126 96
rect 134 94 136 96
rect 144 94 146 96
rect 154 94 156 96
rect 164 94 166 96
rect 174 94 176 96
rect 184 94 186 96
rect 194 94 196 96
rect 204 94 206 96
rect 214 94 216 96
rect 224 94 226 96
rect 234 94 236 96
rect 244 94 246 96
rect 4 84 6 86
rect 14 84 16 86
rect 24 84 26 86
rect 34 84 36 86
rect 44 84 46 86
rect 54 84 56 86
rect 64 84 66 86
rect 74 84 76 86
rect 84 84 86 86
rect 94 84 96 86
rect 104 84 106 86
rect 114 84 116 86
rect 124 84 126 86
rect 134 84 136 86
rect 144 84 146 86
rect 154 84 156 86
rect 164 84 166 86
rect 174 84 176 86
rect 184 84 186 86
rect 194 84 196 86
rect 204 84 206 86
rect 214 84 216 86
rect 224 84 226 86
rect 234 84 236 86
rect 244 84 246 86
rect 4 74 6 76
rect 14 74 16 76
rect 24 74 26 76
rect 34 74 36 76
rect 44 74 46 76
rect 54 74 56 76
rect 64 74 66 76
rect 74 74 76 76
rect 84 74 86 76
rect 94 74 96 76
rect 104 74 106 76
rect 114 74 116 76
rect 124 74 126 76
rect 134 74 136 76
rect 144 74 146 76
rect 154 74 156 76
rect 164 74 166 76
rect 174 74 176 76
rect 184 74 186 76
rect 194 74 196 76
rect 204 74 206 76
rect 214 74 216 76
rect 224 74 226 76
rect 234 74 236 76
rect 244 74 246 76
rect 4 64 6 66
rect 14 64 16 66
rect 24 64 26 66
rect 34 64 36 66
rect 44 64 46 66
rect 54 64 56 66
rect 64 64 66 66
rect 74 64 76 66
rect 84 64 86 66
rect 94 64 96 66
rect 104 64 106 66
rect 114 64 116 66
rect 124 64 126 66
rect 134 64 136 66
rect 144 64 146 66
rect 154 64 156 66
rect 164 64 166 66
rect 174 64 176 66
rect 184 64 186 66
rect 194 64 196 66
rect 204 64 206 66
rect 214 64 216 66
rect 224 64 226 66
rect 234 64 236 66
rect 244 64 246 66
rect 4 54 6 56
rect 14 54 16 56
rect 24 54 26 56
rect 34 54 36 56
rect 44 54 46 56
rect 54 54 56 56
rect 64 54 66 56
rect 74 54 76 56
rect 84 54 86 56
rect 94 54 96 56
rect 104 54 106 56
rect 114 54 116 56
rect 124 54 126 56
rect 134 54 136 56
rect 144 54 146 56
rect 154 54 156 56
rect 164 54 166 56
rect 174 54 176 56
rect 184 54 186 56
rect 194 54 196 56
rect 204 54 206 56
rect 214 54 216 56
rect 224 54 226 56
rect 234 54 236 56
rect 244 54 246 56
rect 4 44 6 46
rect 14 44 16 46
rect 24 44 26 46
rect 34 44 36 46
rect 44 44 46 46
rect 54 44 56 46
rect 64 44 66 46
rect 74 44 76 46
rect 84 44 86 46
rect 94 44 96 46
rect 104 44 106 46
rect 114 44 116 46
rect 124 44 126 46
rect 134 44 136 46
rect 144 44 146 46
rect 154 44 156 46
rect 164 44 166 46
rect 174 44 176 46
rect 184 44 186 46
rect 194 44 196 46
rect 204 44 206 46
rect 214 44 216 46
rect 224 44 226 46
rect 234 44 236 46
rect 244 44 246 46
rect 4 34 6 36
rect 14 34 16 36
rect 24 34 26 36
rect 34 34 36 36
rect 44 34 46 36
rect 54 34 56 36
rect 64 34 66 36
rect 74 34 76 36
rect 84 34 86 36
rect 94 34 96 36
rect 104 34 106 36
rect 114 34 116 36
rect 124 34 126 36
rect 134 34 136 36
rect 144 34 146 36
rect 154 34 156 36
rect 164 34 166 36
rect 174 34 176 36
rect 184 34 186 36
rect 194 34 196 36
rect 204 34 206 36
rect 214 34 216 36
rect 224 34 226 36
rect 234 34 236 36
rect 244 34 246 36
rect 4 24 6 26
rect 14 24 16 26
rect 24 24 26 26
rect 34 24 36 26
rect 44 24 46 26
rect 54 24 56 26
rect 64 24 66 26
rect 74 24 76 26
rect 84 24 86 26
rect 94 24 96 26
rect 104 24 106 26
rect 114 24 116 26
rect 124 24 126 26
rect 134 24 136 26
rect 144 24 146 26
rect 154 24 156 26
rect 164 24 166 26
rect 174 24 176 26
rect 184 24 186 26
rect 194 24 196 26
rect 204 24 206 26
rect 214 24 216 26
rect 224 24 226 26
rect 234 24 236 26
rect 244 24 246 26
rect 4 14 6 16
rect 14 14 16 16
rect 24 14 26 16
rect 34 14 36 16
rect 44 14 46 16
rect 54 14 56 16
rect 64 14 66 16
rect 74 14 76 16
rect 84 14 86 16
rect 94 14 96 16
rect 104 14 106 16
rect 114 14 116 16
rect 124 14 126 16
rect 134 14 136 16
rect 144 14 146 16
rect 154 14 156 16
rect 164 14 166 16
rect 174 14 176 16
rect 184 14 186 16
rect 194 14 196 16
rect 204 14 206 16
rect 214 14 216 16
rect 224 14 226 16
rect 234 14 236 16
rect 244 14 246 16
rect 4 4 6 6
rect 14 4 16 6
rect 24 4 26 6
rect 34 4 36 6
rect 44 4 46 6
rect 54 4 56 6
rect 64 4 66 6
rect 74 4 76 6
rect 84 4 86 6
rect 94 4 96 6
rect 104 4 106 6
rect 114 4 116 6
rect 124 4 126 6
rect 134 4 136 6
rect 144 4 146 6
rect 154 4 156 6
rect 164 4 166 6
rect 174 4 176 6
rect 184 4 186 6
rect 194 4 196 6
rect 204 4 206 6
rect 214 4 216 6
rect 224 4 226 6
rect 234 4 236 6
rect 244 4 246 6
<< metal3 >>
rect -4 250 254 254
rect -4 0 0 250
rect 250 0 254 250
rect -4 -4 254 0
<< gv2 >>
rect 9 239 11 241
rect 19 239 21 241
rect 29 239 31 241
rect 39 239 41 241
rect 49 239 51 241
rect 59 239 61 241
rect 69 239 71 241
rect 79 239 81 241
rect 89 239 91 241
rect 99 239 101 241
rect 109 239 111 241
rect 119 239 121 241
rect 129 239 131 241
rect 139 239 141 241
rect 149 239 151 241
rect 159 239 161 241
rect 169 239 171 241
rect 179 239 181 241
rect 189 239 191 241
rect 199 239 201 241
rect 209 239 211 241
rect 219 239 221 241
rect 229 239 231 241
rect 239 239 241 241
rect 9 229 11 231
rect 19 229 21 231
rect 29 229 31 231
rect 39 229 41 231
rect 49 229 51 231
rect 59 229 61 231
rect 69 229 71 231
rect 79 229 81 231
rect 89 229 91 231
rect 99 229 101 231
rect 109 229 111 231
rect 119 229 121 231
rect 129 229 131 231
rect 139 229 141 231
rect 149 229 151 231
rect 159 229 161 231
rect 169 229 171 231
rect 179 229 181 231
rect 189 229 191 231
rect 199 229 201 231
rect 209 229 211 231
rect 219 229 221 231
rect 229 229 231 231
rect 239 229 241 231
rect 9 219 11 221
rect 19 219 21 221
rect 29 219 31 221
rect 39 219 41 221
rect 49 219 51 221
rect 59 219 61 221
rect 69 219 71 221
rect 79 219 81 221
rect 89 219 91 221
rect 99 219 101 221
rect 109 219 111 221
rect 119 219 121 221
rect 129 219 131 221
rect 139 219 141 221
rect 149 219 151 221
rect 159 219 161 221
rect 169 219 171 221
rect 179 219 181 221
rect 189 219 191 221
rect 199 219 201 221
rect 209 219 211 221
rect 219 219 221 221
rect 229 219 231 221
rect 239 219 241 221
rect 9 209 11 211
rect 19 209 21 211
rect 29 209 31 211
rect 39 209 41 211
rect 49 209 51 211
rect 59 209 61 211
rect 69 209 71 211
rect 79 209 81 211
rect 89 209 91 211
rect 99 209 101 211
rect 109 209 111 211
rect 119 209 121 211
rect 129 209 131 211
rect 139 209 141 211
rect 149 209 151 211
rect 159 209 161 211
rect 169 209 171 211
rect 179 209 181 211
rect 189 209 191 211
rect 199 209 201 211
rect 209 209 211 211
rect 219 209 221 211
rect 229 209 231 211
rect 239 209 241 211
rect 9 199 11 201
rect 19 199 21 201
rect 29 199 31 201
rect 39 199 41 201
rect 49 199 51 201
rect 59 199 61 201
rect 69 199 71 201
rect 79 199 81 201
rect 89 199 91 201
rect 99 199 101 201
rect 109 199 111 201
rect 119 199 121 201
rect 129 199 131 201
rect 139 199 141 201
rect 149 199 151 201
rect 159 199 161 201
rect 169 199 171 201
rect 179 199 181 201
rect 189 199 191 201
rect 199 199 201 201
rect 209 199 211 201
rect 219 199 221 201
rect 229 199 231 201
rect 239 199 241 201
rect 9 189 11 191
rect 19 189 21 191
rect 29 189 31 191
rect 39 189 41 191
rect 49 189 51 191
rect 59 189 61 191
rect 69 189 71 191
rect 79 189 81 191
rect 89 189 91 191
rect 99 189 101 191
rect 109 189 111 191
rect 119 189 121 191
rect 129 189 131 191
rect 139 189 141 191
rect 149 189 151 191
rect 159 189 161 191
rect 169 189 171 191
rect 179 189 181 191
rect 189 189 191 191
rect 199 189 201 191
rect 209 189 211 191
rect 219 189 221 191
rect 229 189 231 191
rect 239 189 241 191
rect 9 179 11 181
rect 19 179 21 181
rect 29 179 31 181
rect 39 179 41 181
rect 49 179 51 181
rect 59 179 61 181
rect 69 179 71 181
rect 79 179 81 181
rect 89 179 91 181
rect 99 179 101 181
rect 109 179 111 181
rect 119 179 121 181
rect 129 179 131 181
rect 139 179 141 181
rect 149 179 151 181
rect 159 179 161 181
rect 169 179 171 181
rect 179 179 181 181
rect 189 179 191 181
rect 199 179 201 181
rect 209 179 211 181
rect 219 179 221 181
rect 229 179 231 181
rect 239 179 241 181
rect 9 169 11 171
rect 19 169 21 171
rect 29 169 31 171
rect 39 169 41 171
rect 49 169 51 171
rect 59 169 61 171
rect 69 169 71 171
rect 79 169 81 171
rect 89 169 91 171
rect 99 169 101 171
rect 109 169 111 171
rect 119 169 121 171
rect 129 169 131 171
rect 139 169 141 171
rect 149 169 151 171
rect 159 169 161 171
rect 169 169 171 171
rect 179 169 181 171
rect 189 169 191 171
rect 199 169 201 171
rect 209 169 211 171
rect 219 169 221 171
rect 229 169 231 171
rect 239 169 241 171
rect 9 159 11 161
rect 19 159 21 161
rect 29 159 31 161
rect 39 159 41 161
rect 49 159 51 161
rect 59 159 61 161
rect 69 159 71 161
rect 79 159 81 161
rect 89 159 91 161
rect 99 159 101 161
rect 109 159 111 161
rect 119 159 121 161
rect 129 159 131 161
rect 139 159 141 161
rect 149 159 151 161
rect 159 159 161 161
rect 169 159 171 161
rect 179 159 181 161
rect 189 159 191 161
rect 199 159 201 161
rect 209 159 211 161
rect 219 159 221 161
rect 229 159 231 161
rect 239 159 241 161
rect 9 149 11 151
rect 19 149 21 151
rect 29 149 31 151
rect 39 149 41 151
rect 49 149 51 151
rect 59 149 61 151
rect 69 149 71 151
rect 79 149 81 151
rect 89 149 91 151
rect 99 149 101 151
rect 109 149 111 151
rect 119 149 121 151
rect 129 149 131 151
rect 139 149 141 151
rect 149 149 151 151
rect 159 149 161 151
rect 169 149 171 151
rect 179 149 181 151
rect 189 149 191 151
rect 199 149 201 151
rect 209 149 211 151
rect 219 149 221 151
rect 229 149 231 151
rect 239 149 241 151
rect 9 139 11 141
rect 19 139 21 141
rect 29 139 31 141
rect 39 139 41 141
rect 49 139 51 141
rect 59 139 61 141
rect 69 139 71 141
rect 79 139 81 141
rect 89 139 91 141
rect 99 139 101 141
rect 109 139 111 141
rect 119 139 121 141
rect 129 139 131 141
rect 139 139 141 141
rect 149 139 151 141
rect 159 139 161 141
rect 169 139 171 141
rect 179 139 181 141
rect 189 139 191 141
rect 199 139 201 141
rect 209 139 211 141
rect 219 139 221 141
rect 229 139 231 141
rect 239 139 241 141
rect 9 129 11 131
rect 19 129 21 131
rect 29 129 31 131
rect 39 129 41 131
rect 49 129 51 131
rect 59 129 61 131
rect 69 129 71 131
rect 79 129 81 131
rect 89 129 91 131
rect 99 129 101 131
rect 109 129 111 131
rect 119 129 121 131
rect 129 129 131 131
rect 139 129 141 131
rect 149 129 151 131
rect 159 129 161 131
rect 169 129 171 131
rect 179 129 181 131
rect 189 129 191 131
rect 199 129 201 131
rect 209 129 211 131
rect 219 129 221 131
rect 229 129 231 131
rect 239 129 241 131
rect 9 119 11 121
rect 19 119 21 121
rect 29 119 31 121
rect 39 119 41 121
rect 49 119 51 121
rect 59 119 61 121
rect 69 119 71 121
rect 79 119 81 121
rect 89 119 91 121
rect 99 119 101 121
rect 109 119 111 121
rect 119 119 121 121
rect 129 119 131 121
rect 139 119 141 121
rect 149 119 151 121
rect 159 119 161 121
rect 169 119 171 121
rect 179 119 181 121
rect 189 119 191 121
rect 199 119 201 121
rect 209 119 211 121
rect 219 119 221 121
rect 229 119 231 121
rect 239 119 241 121
rect 9 109 11 111
rect 19 109 21 111
rect 29 109 31 111
rect 39 109 41 111
rect 49 109 51 111
rect 59 109 61 111
rect 69 109 71 111
rect 79 109 81 111
rect 89 109 91 111
rect 99 109 101 111
rect 109 109 111 111
rect 119 109 121 111
rect 129 109 131 111
rect 139 109 141 111
rect 149 109 151 111
rect 159 109 161 111
rect 169 109 171 111
rect 179 109 181 111
rect 189 109 191 111
rect 199 109 201 111
rect 209 109 211 111
rect 219 109 221 111
rect 229 109 231 111
rect 239 109 241 111
rect 9 99 11 101
rect 19 99 21 101
rect 29 99 31 101
rect 39 99 41 101
rect 49 99 51 101
rect 59 99 61 101
rect 69 99 71 101
rect 79 99 81 101
rect 89 99 91 101
rect 99 99 101 101
rect 109 99 111 101
rect 119 99 121 101
rect 129 99 131 101
rect 139 99 141 101
rect 149 99 151 101
rect 159 99 161 101
rect 169 99 171 101
rect 179 99 181 101
rect 189 99 191 101
rect 199 99 201 101
rect 209 99 211 101
rect 219 99 221 101
rect 229 99 231 101
rect 239 99 241 101
rect 9 89 11 91
rect 19 89 21 91
rect 29 89 31 91
rect 39 89 41 91
rect 49 89 51 91
rect 59 89 61 91
rect 69 89 71 91
rect 79 89 81 91
rect 89 89 91 91
rect 99 89 101 91
rect 109 89 111 91
rect 119 89 121 91
rect 129 89 131 91
rect 139 89 141 91
rect 149 89 151 91
rect 159 89 161 91
rect 169 89 171 91
rect 179 89 181 91
rect 189 89 191 91
rect 199 89 201 91
rect 209 89 211 91
rect 219 89 221 91
rect 229 89 231 91
rect 239 89 241 91
rect 9 79 11 81
rect 19 79 21 81
rect 29 79 31 81
rect 39 79 41 81
rect 49 79 51 81
rect 59 79 61 81
rect 69 79 71 81
rect 79 79 81 81
rect 89 79 91 81
rect 99 79 101 81
rect 109 79 111 81
rect 119 79 121 81
rect 129 79 131 81
rect 139 79 141 81
rect 149 79 151 81
rect 159 79 161 81
rect 169 79 171 81
rect 179 79 181 81
rect 189 79 191 81
rect 199 79 201 81
rect 209 79 211 81
rect 219 79 221 81
rect 229 79 231 81
rect 239 79 241 81
rect 9 69 11 71
rect 19 69 21 71
rect 29 69 31 71
rect 39 69 41 71
rect 49 69 51 71
rect 59 69 61 71
rect 69 69 71 71
rect 79 69 81 71
rect 89 69 91 71
rect 99 69 101 71
rect 109 69 111 71
rect 119 69 121 71
rect 129 69 131 71
rect 139 69 141 71
rect 149 69 151 71
rect 159 69 161 71
rect 169 69 171 71
rect 179 69 181 71
rect 189 69 191 71
rect 199 69 201 71
rect 209 69 211 71
rect 219 69 221 71
rect 229 69 231 71
rect 239 69 241 71
rect 9 59 11 61
rect 19 59 21 61
rect 29 59 31 61
rect 39 59 41 61
rect 49 59 51 61
rect 59 59 61 61
rect 69 59 71 61
rect 79 59 81 61
rect 89 59 91 61
rect 99 59 101 61
rect 109 59 111 61
rect 119 59 121 61
rect 129 59 131 61
rect 139 59 141 61
rect 149 59 151 61
rect 159 59 161 61
rect 169 59 171 61
rect 179 59 181 61
rect 189 59 191 61
rect 199 59 201 61
rect 209 59 211 61
rect 219 59 221 61
rect 229 59 231 61
rect 239 59 241 61
rect 9 49 11 51
rect 19 49 21 51
rect 29 49 31 51
rect 39 49 41 51
rect 49 49 51 51
rect 59 49 61 51
rect 69 49 71 51
rect 79 49 81 51
rect 89 49 91 51
rect 99 49 101 51
rect 109 49 111 51
rect 119 49 121 51
rect 129 49 131 51
rect 139 49 141 51
rect 149 49 151 51
rect 159 49 161 51
rect 169 49 171 51
rect 179 49 181 51
rect 189 49 191 51
rect 199 49 201 51
rect 209 49 211 51
rect 219 49 221 51
rect 229 49 231 51
rect 239 49 241 51
rect 9 39 11 41
rect 19 39 21 41
rect 29 39 31 41
rect 39 39 41 41
rect 49 39 51 41
rect 59 39 61 41
rect 69 39 71 41
rect 79 39 81 41
rect 89 39 91 41
rect 99 39 101 41
rect 109 39 111 41
rect 119 39 121 41
rect 129 39 131 41
rect 139 39 141 41
rect 149 39 151 41
rect 159 39 161 41
rect 169 39 171 41
rect 179 39 181 41
rect 189 39 191 41
rect 199 39 201 41
rect 209 39 211 41
rect 219 39 221 41
rect 229 39 231 41
rect 239 39 241 41
rect 9 29 11 31
rect 19 29 21 31
rect 29 29 31 31
rect 39 29 41 31
rect 49 29 51 31
rect 59 29 61 31
rect 69 29 71 31
rect 79 29 81 31
rect 89 29 91 31
rect 99 29 101 31
rect 109 29 111 31
rect 119 29 121 31
rect 129 29 131 31
rect 139 29 141 31
rect 149 29 151 31
rect 159 29 161 31
rect 169 29 171 31
rect 179 29 181 31
rect 189 29 191 31
rect 199 29 201 31
rect 209 29 211 31
rect 219 29 221 31
rect 229 29 231 31
rect 239 29 241 31
rect 9 19 11 21
rect 19 19 21 21
rect 29 19 31 21
rect 39 19 41 21
rect 49 19 51 21
rect 59 19 61 21
rect 69 19 71 21
rect 79 19 81 21
rect 89 19 91 21
rect 99 19 101 21
rect 109 19 111 21
rect 119 19 121 21
rect 129 19 131 21
rect 139 19 141 21
rect 149 19 151 21
rect 159 19 161 21
rect 169 19 171 21
rect 179 19 181 21
rect 189 19 191 21
rect 199 19 201 21
rect 209 19 211 21
rect 219 19 221 21
rect 229 19 231 21
rect 239 19 241 21
rect 9 9 11 11
rect 19 9 21 11
rect 29 9 31 11
rect 39 9 41 11
rect 49 9 51 11
rect 59 9 61 11
rect 69 9 71 11
rect 79 9 81 11
rect 89 9 91 11
rect 99 9 101 11
rect 109 9 111 11
rect 119 9 121 11
rect 129 9 131 11
rect 139 9 141 11
rect 149 9 151 11
rect 159 9 161 11
rect 169 9 171 11
rect 179 9 181 11
rect 189 9 191 11
rect 199 9 201 11
rect 209 9 211 11
rect 219 9 221 11
rect 229 9 231 11
rect 239 9 241 11
<< pad >>
rect 0 0 250 250
<< end >>
