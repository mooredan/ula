magic
tech amic5n
timestamp 1608937081
<< nwell >>
rect -160 850 830 2500
<< ntransistor >>
rect 110 450 170 700
rect 500 140 560 700
<< ptransistor >>
rect 110 1000 170 1510
rect 500 1000 560 2350
<< nselect >>
rect 70 1670 240 1900
rect -55 360 725 730
rect -55 190 70 360
rect 240 190 725 360
rect -55 45 725 190
<< pselect >>
rect -55 1900 725 2445
rect -55 1670 70 1900
rect 240 1670 725 1900
rect -55 970 725 1670
rect 70 190 240 360
<< ndiffusion >>
rect -10 670 110 700
rect -10 620 20 670
rect 70 620 110 670
rect -10 530 110 620
rect -10 480 20 530
rect 70 480 110 530
rect -10 450 110 480
rect 170 670 290 700
rect 170 620 210 670
rect 260 620 290 670
rect 170 530 290 620
rect 170 480 210 530
rect 260 480 290 530
rect 170 450 290 480
rect 380 670 500 700
rect 380 620 410 670
rect 460 620 500 670
rect 380 520 500 620
rect 380 470 410 520
rect 460 470 500 520
rect 380 420 500 470
rect 380 370 410 420
rect 460 370 500 420
rect 380 320 500 370
rect 380 270 410 320
rect 460 270 500 320
rect 380 220 500 270
rect 380 170 410 220
rect 460 170 500 220
rect 380 140 500 170
rect 560 670 680 700
rect 560 620 600 670
rect 650 620 680 670
rect 560 520 680 620
rect 560 470 600 520
rect 650 470 680 520
rect 560 420 680 470
rect 560 370 600 420
rect 650 370 680 420
rect 560 320 680 370
rect 560 270 600 320
rect 650 270 680 320
rect 560 220 680 270
rect 560 170 600 220
rect 650 170 680 220
rect 560 140 680 170
<< pdiffusion >>
rect 380 2320 500 2350
rect 380 2270 410 2320
rect 460 2270 500 2320
rect 380 2180 500 2270
rect 380 2130 410 2180
rect 460 2130 500 2180
rect 380 2080 500 2130
rect 380 2030 410 2080
rect 460 2030 500 2080
rect 380 1980 500 2030
rect 380 1930 410 1980
rect 460 1930 500 1980
rect 380 1880 500 1930
rect 380 1830 410 1880
rect 460 1830 500 1880
rect 380 1780 500 1830
rect 380 1730 410 1780
rect 460 1730 500 1780
rect 380 1680 500 1730
rect 380 1630 410 1680
rect 460 1630 500 1680
rect 380 1580 500 1630
rect 380 1530 410 1580
rect 460 1530 500 1580
rect -10 1480 110 1510
rect -10 1430 20 1480
rect 70 1430 110 1480
rect -10 1380 110 1430
rect -10 1330 20 1380
rect 70 1330 110 1380
rect -10 1280 110 1330
rect -10 1230 20 1280
rect 70 1230 110 1280
rect -10 1180 110 1230
rect -10 1130 20 1180
rect 70 1130 110 1180
rect -10 1080 110 1130
rect -10 1030 20 1080
rect 70 1030 110 1080
rect -10 1000 110 1030
rect 170 1480 290 1510
rect 170 1430 210 1480
rect 260 1430 290 1480
rect 170 1380 290 1430
rect 170 1330 210 1380
rect 260 1330 290 1380
rect 170 1280 290 1330
rect 170 1230 210 1280
rect 260 1230 290 1280
rect 170 1180 290 1230
rect 170 1130 210 1180
rect 260 1130 290 1180
rect 170 1080 290 1130
rect 170 1030 210 1080
rect 260 1030 290 1080
rect 170 1000 290 1030
rect 380 1480 500 1530
rect 380 1430 410 1480
rect 460 1430 500 1480
rect 380 1380 500 1430
rect 380 1330 410 1380
rect 460 1330 500 1380
rect 380 1280 500 1330
rect 380 1230 410 1280
rect 460 1230 500 1280
rect 380 1180 500 1230
rect 380 1130 410 1180
rect 460 1130 500 1180
rect 380 1080 500 1130
rect 380 1030 410 1080
rect 460 1030 500 1080
rect 380 1000 500 1030
rect 560 2320 680 2350
rect 560 2270 600 2320
rect 650 2270 680 2320
rect 560 2180 680 2270
rect 560 2130 600 2180
rect 650 2130 680 2180
rect 560 2080 680 2130
rect 560 2030 600 2080
rect 650 2030 680 2080
rect 560 1980 680 2030
rect 560 1930 600 1980
rect 650 1930 680 1980
rect 560 1880 680 1930
rect 560 1830 600 1880
rect 650 1830 680 1880
rect 560 1780 680 1830
rect 560 1730 600 1780
rect 650 1730 680 1780
rect 560 1680 680 1730
rect 560 1630 600 1680
rect 650 1630 680 1680
rect 560 1580 680 1630
rect 560 1530 600 1580
rect 650 1530 680 1580
rect 560 1480 680 1530
rect 560 1430 600 1480
rect 650 1430 680 1480
rect 560 1380 680 1430
rect 560 1330 600 1380
rect 650 1330 680 1380
rect 560 1280 680 1330
rect 560 1230 600 1280
rect 650 1230 680 1280
rect 560 1180 680 1230
rect 560 1130 600 1180
rect 650 1130 680 1180
rect 560 1080 680 1130
rect 560 1030 600 1080
rect 650 1030 680 1080
rect 560 1000 680 1030
<< psubstratepdiff >>
rect 100 300 210 330
rect 100 250 130 300
rect 180 250 210 300
rect 100 220 210 250
<< nsubstratendiff >>
rect 100 1780 210 1870
rect 100 1730 130 1780
rect 180 1730 210 1780
rect 100 1700 210 1730
<< nsubstratencontact >>
rect 130 1730 180 1780
<< psubstratepcontact >>
rect 130 250 180 300
<< ndcontact >>
rect 20 620 70 670
rect 20 480 70 530
rect 210 620 260 670
rect 210 480 260 530
rect 410 620 460 670
rect 410 470 460 520
rect 410 370 460 420
rect 410 270 460 320
rect 410 170 460 220
rect 600 620 650 670
rect 600 470 650 520
rect 600 370 650 420
rect 600 270 650 320
rect 600 170 650 220
<< pdcontact >>
rect 410 2270 460 2320
rect 410 2130 460 2180
rect 410 2030 460 2080
rect 410 1930 460 1980
rect 410 1830 460 1880
rect 410 1730 460 1780
rect 410 1630 460 1680
rect 410 1530 460 1580
rect 20 1430 70 1480
rect 20 1330 70 1380
rect 20 1230 70 1280
rect 20 1130 70 1180
rect 20 1030 70 1080
rect 210 1430 260 1480
rect 210 1330 260 1380
rect 210 1230 260 1280
rect 210 1130 260 1180
rect 210 1030 260 1080
rect 410 1430 460 1480
rect 410 1330 460 1380
rect 410 1230 460 1280
rect 410 1130 460 1180
rect 410 1030 460 1080
rect 600 2270 650 2320
rect 600 2130 650 2180
rect 600 2030 650 2080
rect 600 1930 650 1980
rect 600 1830 650 1880
rect 600 1730 650 1780
rect 600 1630 650 1680
rect 600 1530 650 1580
rect 600 1430 650 1480
rect 600 1330 650 1380
rect 600 1230 650 1280
rect 600 1130 650 1180
rect 600 1030 650 1080
<< polysilicon >>
rect 500 2350 560 2415
rect 110 1510 170 1575
rect 110 890 170 1000
rect 500 890 560 1000
rect 0 870 170 890
rect 0 820 20 870
rect 70 820 170 870
rect 0 800 170 820
rect 390 870 560 890
rect 390 820 410 870
rect 460 820 560 870
rect 390 800 560 820
rect 110 700 170 800
rect 500 700 560 800
rect 110 385 170 450
rect 500 75 560 140
<< polycontact >>
rect 20 820 70 870
rect 410 820 460 870
<< metal1 >>
rect 0 2400 670 2490
rect 0 1800 90 2400
rect 390 2320 480 2400
rect 390 2270 410 2320
rect 460 2270 480 2320
rect 390 2180 480 2270
rect 390 2130 410 2180
rect 460 2130 480 2180
rect 390 2080 480 2130
rect 390 2030 410 2080
rect 460 2030 480 2080
rect 390 1980 480 2030
rect 390 1930 410 1980
rect 460 1930 480 1980
rect 390 1880 480 1930
rect 390 1830 410 1880
rect 460 1830 480 1880
rect 0 1780 200 1800
rect 0 1730 130 1780
rect 180 1730 200 1780
rect 0 1710 200 1730
rect 390 1780 480 1830
rect 390 1730 410 1780
rect 460 1730 480 1780
rect 0 1480 90 1710
rect 390 1680 480 1730
rect 390 1630 410 1680
rect 460 1630 480 1680
rect 390 1580 480 1630
rect 390 1530 410 1580
rect 460 1530 480 1580
rect 0 1430 20 1480
rect 70 1430 90 1480
rect 0 1380 90 1430
rect 0 1330 20 1380
rect 70 1330 90 1380
rect 0 1280 90 1330
rect 0 1230 20 1280
rect 70 1230 90 1280
rect 0 1180 90 1230
rect 0 1130 20 1180
rect 70 1130 90 1180
rect 0 1080 90 1130
rect 0 1030 20 1080
rect 70 1030 90 1080
rect 0 1010 90 1030
rect 190 1480 280 1500
rect 190 1430 210 1480
rect 260 1430 280 1480
rect 190 1380 280 1430
rect 190 1330 210 1380
rect 260 1330 280 1380
rect 190 1280 280 1330
rect 190 1230 210 1280
rect 260 1230 280 1280
rect 190 1180 280 1230
rect 190 1130 210 1180
rect 260 1130 280 1180
rect 190 1080 280 1130
rect 190 1030 210 1080
rect 260 1030 280 1080
rect 190 890 280 1030
rect 390 1480 480 1530
rect 390 1430 410 1480
rect 460 1430 480 1480
rect 390 1380 480 1430
rect 390 1330 410 1380
rect 460 1330 480 1380
rect 390 1280 480 1330
rect 390 1230 410 1280
rect 460 1230 480 1280
rect 390 1180 480 1230
rect 390 1130 410 1180
rect 460 1130 480 1180
rect 390 1080 480 1130
rect 390 1030 410 1080
rect 460 1030 480 1080
rect 390 1010 480 1030
rect 580 2320 670 2340
rect 580 2270 600 2320
rect 650 2270 670 2320
rect 580 2180 670 2270
rect 580 2130 600 2180
rect 650 2130 670 2180
rect 580 2080 670 2130
rect 580 2030 600 2080
rect 650 2030 670 2080
rect 580 1980 670 2030
rect 580 1930 600 1980
rect 650 1930 670 1980
rect 580 1880 670 1930
rect 580 1830 600 1880
rect 650 1830 670 1880
rect 580 1780 670 1830
rect 580 1730 600 1780
rect 650 1730 670 1780
rect 580 1680 670 1730
rect 580 1630 600 1680
rect 650 1630 670 1680
rect 580 1580 670 1630
rect 580 1530 600 1580
rect 650 1530 670 1580
rect 580 1480 670 1530
rect 580 1430 600 1480
rect 650 1430 670 1480
rect 580 1380 670 1430
rect 580 1330 600 1380
rect 650 1330 670 1380
rect 580 1280 670 1330
rect 580 1230 600 1280
rect 650 1230 670 1280
rect 580 1180 670 1230
rect 580 1130 600 1180
rect 650 1130 670 1180
rect 580 1080 670 1130
rect 580 1030 600 1080
rect 650 1030 670 1080
rect 0 870 90 890
rect 0 820 20 870
rect 70 820 90 870
rect 0 800 90 820
rect 190 870 480 890
rect 190 820 410 870
rect 460 820 480 870
rect 190 800 480 820
rect 0 670 90 690
rect 0 620 20 670
rect 70 620 90 670
rect 0 530 90 620
rect 0 480 20 530
rect 70 480 90 530
rect 0 320 90 480
rect 190 670 280 800
rect 190 620 210 670
rect 260 620 280 670
rect 190 530 280 620
rect 190 480 210 530
rect 260 480 280 530
rect 190 460 280 480
rect 390 670 480 690
rect 390 620 410 670
rect 460 620 480 670
rect 390 520 480 620
rect 390 470 410 520
rect 460 470 480 520
rect 390 420 480 470
rect 390 370 410 420
rect 460 370 480 420
rect 390 320 480 370
rect 0 300 200 320
rect 0 250 130 300
rect 180 250 200 300
rect 0 230 200 250
rect 390 270 410 320
rect 460 270 480 320
rect 0 90 90 230
rect 390 220 480 270
rect 390 170 410 220
rect 460 170 480 220
rect 390 90 480 170
rect 580 670 670 1030
rect 580 620 600 670
rect 650 620 670 670
rect 580 520 670 620
rect 580 470 600 520
rect 650 470 670 520
rect 580 420 670 470
rect 580 370 600 420
rect 650 370 670 420
rect 580 320 670 370
rect 580 270 600 320
rect 650 270 670 320
rect 580 220 670 270
rect 580 170 600 220
rect 650 170 670 220
rect 580 150 670 170
rect 0 0 670 90
<< labels >>
flabel metal1 s 20 20 20 20 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 20 810 20 810 2 FreeSans 400 0 0 0 a
port 2 ne
flabel metal1 s 10 2430 10 2430 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel nwell 700 900 700 900 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 610 770 610 770 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 290 820 290 820 2 FreeSans 400 0 0 0 n1
<< end >>
