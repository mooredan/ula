magic
tech amic5n
timestamp 1624420999
<< nwell >>
rect -130 550 2080 1495
<< ntransistor >>
rect 165 95 225 400
rect 800 95 860 400
rect 1345 125 1405 400
rect 1535 125 1595 400
rect 1725 125 1785 400
<< ptransistor >>
rect 165 700 225 1345
rect 355 700 415 1345
rect 610 700 670 1345
rect 800 700 860 1345
rect 1345 705 1405 1290
rect 1535 705 1595 1290
rect 1725 705 1785 1290
<< nselect >>
rect 1060 765 1225 1290
rect -10 350 1960 430
rect -10 295 1060 350
rect -10 100 400 295
rect 630 125 1060 295
rect 1225 125 1960 350
rect 630 100 1960 125
rect -10 0 1960 100
<< pselect >>
rect -10 1290 1960 1440
rect -10 765 1060 1290
rect 1225 765 1960 1290
rect -10 670 1960 765
rect 400 100 630 295
rect 1060 125 1225 350
<< ndiffusion >>
rect 45 370 165 400
rect 45 320 75 370
rect 125 320 165 370
rect 45 175 165 320
rect 45 125 75 175
rect 125 125 165 175
rect 45 95 165 125
rect 225 370 345 400
rect 225 320 265 370
rect 315 320 345 370
rect 225 175 345 320
rect 680 370 800 400
rect 680 320 710 370
rect 760 320 800 370
rect 225 125 265 175
rect 315 125 345 175
rect 680 175 800 320
rect 225 95 345 125
rect 680 125 710 175
rect 760 125 800 175
rect 680 95 800 125
rect 860 355 980 400
rect 860 305 900 355
rect 950 305 980 355
rect 1225 370 1345 400
rect 860 175 980 305
rect 860 125 900 175
rect 950 125 980 175
rect 1225 320 1255 370
rect 1305 320 1345 370
rect 1225 205 1345 320
rect 1225 155 1255 205
rect 1305 155 1345 205
rect 1225 125 1345 155
rect 1405 370 1535 400
rect 1405 320 1445 370
rect 1495 320 1535 370
rect 1405 205 1535 320
rect 1405 155 1445 205
rect 1495 155 1535 205
rect 1405 125 1535 155
rect 1595 345 1725 400
rect 1595 295 1635 345
rect 1685 295 1725 345
rect 1595 205 1725 295
rect 1595 155 1635 205
rect 1685 155 1725 205
rect 1595 125 1725 155
rect 1785 370 1905 400
rect 1785 320 1825 370
rect 1875 320 1905 370
rect 1785 205 1905 320
rect 1785 155 1825 205
rect 1875 155 1905 205
rect 1785 125 1905 155
rect 860 95 980 125
<< pdiffusion >>
rect 45 1315 165 1345
rect 45 1265 75 1315
rect 125 1265 165 1315
rect 45 1200 165 1265
rect 45 1150 75 1200
rect 125 1150 165 1200
rect 45 1065 165 1150
rect 45 1015 75 1065
rect 125 1015 165 1065
rect 45 945 165 1015
rect 45 895 75 945
rect 125 895 165 945
rect 45 825 165 895
rect 45 775 75 825
rect 125 775 165 825
rect 45 700 165 775
rect 225 1315 355 1345
rect 225 1265 265 1315
rect 315 1265 355 1315
rect 225 1215 355 1265
rect 225 1165 265 1215
rect 315 1165 355 1215
rect 225 1115 355 1165
rect 225 1065 265 1115
rect 315 1065 355 1115
rect 225 985 355 1065
rect 225 935 265 985
rect 315 935 355 985
rect 225 700 355 935
rect 415 1315 610 1345
rect 415 1265 475 1315
rect 525 1265 610 1315
rect 415 1200 610 1265
rect 415 1150 475 1200
rect 525 1150 610 1200
rect 415 1065 610 1150
rect 415 1015 475 1065
rect 525 1015 610 1065
rect 415 945 610 1015
rect 415 895 475 945
rect 525 895 610 945
rect 415 825 610 895
rect 415 775 475 825
rect 525 775 610 825
rect 415 700 610 775
rect 670 1155 800 1345
rect 670 1105 710 1155
rect 760 1105 800 1155
rect 670 1015 800 1105
rect 670 965 710 1015
rect 760 965 800 1015
rect 670 915 800 965
rect 670 865 710 915
rect 760 865 800 915
rect 670 815 800 865
rect 670 765 710 815
rect 760 765 800 815
rect 670 700 800 765
rect 860 1315 980 1345
rect 860 1265 900 1315
rect 950 1265 980 1315
rect 860 1215 980 1265
rect 860 1165 900 1215
rect 950 1165 980 1215
rect 860 1115 980 1165
rect 860 1065 900 1115
rect 950 1065 980 1115
rect 860 1015 980 1065
rect 860 965 900 1015
rect 950 965 980 1015
rect 860 915 980 965
rect 860 865 900 915
rect 950 865 980 915
rect 860 815 980 865
rect 860 765 900 815
rect 950 765 980 815
rect 1225 1260 1345 1290
rect 1225 1210 1255 1260
rect 1305 1210 1345 1260
rect 1225 1115 1345 1210
rect 1225 1065 1255 1115
rect 1305 1065 1345 1115
rect 1225 1015 1345 1065
rect 1225 965 1255 1015
rect 1305 965 1345 1015
rect 1225 915 1345 965
rect 1225 865 1255 915
rect 1305 865 1345 915
rect 1225 815 1345 865
rect 1225 765 1255 815
rect 1305 765 1345 815
rect 860 700 980 765
rect 1225 705 1345 765
rect 1405 1260 1535 1290
rect 1405 1210 1445 1260
rect 1495 1210 1535 1260
rect 1405 1080 1535 1210
rect 1405 1030 1445 1080
rect 1495 1030 1535 1080
rect 1405 980 1535 1030
rect 1405 930 1445 980
rect 1495 930 1535 980
rect 1405 825 1535 930
rect 1405 775 1445 825
rect 1495 775 1535 825
rect 1405 705 1535 775
rect 1595 1260 1725 1290
rect 1595 1210 1635 1260
rect 1685 1210 1725 1260
rect 1595 1115 1725 1210
rect 1595 1065 1635 1115
rect 1685 1065 1725 1115
rect 1595 975 1725 1065
rect 1595 925 1635 975
rect 1685 925 1725 975
rect 1595 705 1725 925
rect 1785 1260 1905 1290
rect 1785 1210 1825 1260
rect 1875 1210 1905 1260
rect 1785 1085 1905 1210
rect 1785 1035 1825 1085
rect 1875 1035 1905 1085
rect 1785 985 1905 1035
rect 1785 935 1825 985
rect 1875 935 1905 985
rect 1785 885 1905 935
rect 1785 835 1825 885
rect 1875 835 1905 885
rect 1785 785 1905 835
rect 1785 735 1825 785
rect 1875 735 1905 785
rect 1785 705 1905 735
<< psubstratepdiff >>
rect 455 220 565 250
rect 455 170 485 220
rect 535 170 565 220
rect 455 140 565 170
rect 1110 320 1225 350
rect 1110 270 1140 320
rect 1190 270 1225 320
rect 1110 205 1225 270
rect 1110 155 1140 205
rect 1190 155 1225 205
rect 1110 125 1225 155
<< nsubstratendiff >>
rect 1110 1260 1225 1290
rect 1110 1210 1145 1260
rect 1195 1210 1225 1260
rect 1110 1160 1225 1210
rect 1110 1110 1140 1160
rect 1190 1110 1225 1160
rect 1110 1060 1225 1110
rect 1110 1010 1140 1060
rect 1190 1010 1225 1060
rect 1110 960 1225 1010
rect 1110 910 1140 960
rect 1190 910 1225 960
rect 1110 855 1225 910
rect 1110 805 1140 855
rect 1190 805 1225 855
rect 1110 765 1225 805
<< nsubstratencontact >>
rect 1145 1210 1195 1260
rect 1140 1110 1190 1160
rect 1140 1010 1190 1060
rect 1140 910 1190 960
rect 1140 805 1190 855
<< psubstratepcontact >>
rect 485 170 535 220
rect 1140 270 1190 320
rect 1140 155 1190 205
<< ndcontact >>
rect 75 320 125 370
rect 75 125 125 175
rect 265 320 315 370
rect 710 320 760 370
rect 265 125 315 175
rect 710 125 760 175
rect 900 305 950 355
rect 900 125 950 175
rect 1255 320 1305 370
rect 1255 155 1305 205
rect 1445 320 1495 370
rect 1445 155 1495 205
rect 1635 295 1685 345
rect 1635 155 1685 205
rect 1825 320 1875 370
rect 1825 155 1875 205
<< pdcontact >>
rect 75 1265 125 1315
rect 75 1150 125 1200
rect 75 1015 125 1065
rect 75 895 125 945
rect 75 775 125 825
rect 265 1265 315 1315
rect 265 1165 315 1215
rect 265 1065 315 1115
rect 265 935 315 985
rect 475 1265 525 1315
rect 475 1150 525 1200
rect 475 1015 525 1065
rect 475 895 525 945
rect 475 775 525 825
rect 710 1105 760 1155
rect 710 965 760 1015
rect 710 865 760 915
rect 710 765 760 815
rect 900 1265 950 1315
rect 900 1165 950 1215
rect 900 1065 950 1115
rect 900 965 950 1015
rect 900 865 950 915
rect 900 765 950 815
rect 1255 1210 1305 1260
rect 1255 1065 1305 1115
rect 1255 965 1305 1015
rect 1255 865 1305 915
rect 1255 765 1305 815
rect 1445 1210 1495 1260
rect 1445 1030 1495 1080
rect 1445 930 1495 980
rect 1445 775 1495 825
rect 1635 1210 1685 1260
rect 1635 1065 1685 1115
rect 1635 925 1685 975
rect 1825 1210 1875 1260
rect 1825 1035 1875 1085
rect 1825 935 1875 985
rect 1825 835 1875 885
rect 1825 735 1875 785
<< polysilicon >>
rect 165 1345 225 1410
rect 355 1345 415 1410
rect 610 1345 670 1410
rect 800 1345 860 1410
rect 1345 1290 1405 1355
rect 1535 1290 1595 1355
rect 1725 1290 1785 1355
rect 165 630 225 700
rect 355 630 415 700
rect 165 610 415 630
rect 165 560 225 610
rect 275 560 415 610
rect 165 540 415 560
rect 165 400 225 540
rect 610 525 670 700
rect 800 525 860 700
rect 1345 685 1405 705
rect 1535 685 1595 705
rect 1725 685 1785 705
rect 1235 665 1785 685
rect 1235 615 1255 665
rect 1305 615 1355 665
rect 1405 615 1455 665
rect 1505 615 1555 665
rect 1605 615 1655 665
rect 1705 615 1785 665
rect 1235 595 1785 615
rect 610 505 1020 525
rect 610 455 950 505
rect 1000 455 1020 505
rect 610 435 1020 455
rect 800 400 860 435
rect 1345 400 1405 595
rect 1535 400 1595 595
rect 1725 400 1785 595
rect 165 30 225 95
rect 800 30 860 95
rect 1345 60 1405 125
rect 1535 60 1595 125
rect 1725 60 1785 125
<< polycontact >>
rect 225 560 275 610
rect 1255 615 1305 665
rect 1355 615 1405 665
rect 1455 615 1505 665
rect 1555 615 1605 665
rect 1655 615 1705 665
rect 950 455 1000 505
<< metal1 >>
rect 0 1395 1950 1485
rect 55 1315 145 1335
rect 55 1265 75 1315
rect 125 1265 145 1315
rect 55 1200 145 1265
rect 55 1150 75 1200
rect 125 1150 145 1200
rect 55 1065 145 1150
rect 55 1015 75 1065
rect 125 1015 145 1065
rect 55 945 145 1015
rect 55 895 75 945
rect 125 895 145 945
rect 245 1315 335 1395
rect 245 1265 265 1315
rect 315 1265 335 1315
rect 245 1215 335 1265
rect 245 1165 265 1215
rect 315 1165 335 1215
rect 245 1115 335 1165
rect 245 1065 265 1115
rect 315 1065 335 1115
rect 245 985 335 1065
rect 245 935 265 985
rect 315 935 335 985
rect 245 915 335 935
rect 455 1325 545 1335
rect 880 1325 970 1335
rect 455 1315 970 1325
rect 455 1265 475 1315
rect 525 1265 900 1315
rect 950 1265 970 1315
rect 455 1235 970 1265
rect 455 1200 545 1235
rect 455 1150 475 1200
rect 525 1150 545 1200
rect 880 1215 970 1235
rect 455 1065 545 1150
rect 455 1015 475 1065
rect 525 1015 545 1065
rect 455 945 545 1015
rect 55 845 145 895
rect 455 895 475 945
rect 525 895 545 945
rect 455 845 545 895
rect 55 825 545 845
rect 55 775 75 825
rect 125 775 475 825
rect 525 775 545 825
rect 55 755 545 775
rect 690 1155 780 1175
rect 690 1105 710 1155
rect 760 1105 780 1155
rect 690 1015 780 1105
rect 690 965 710 1015
rect 760 965 780 1015
rect 690 915 780 965
rect 690 865 710 915
rect 760 865 780 915
rect 690 815 780 865
rect 690 765 710 815
rect 760 765 780 815
rect 690 685 780 765
rect 880 1165 900 1215
rect 950 1165 970 1215
rect 880 1115 970 1165
rect 880 1065 900 1115
rect 950 1065 970 1115
rect 880 1015 970 1065
rect 880 965 900 1015
rect 950 965 970 1015
rect 880 915 970 965
rect 880 865 900 915
rect 950 865 970 915
rect 880 815 970 865
rect 880 765 900 815
rect 950 765 970 815
rect 880 745 970 765
rect 1120 1260 1325 1395
rect 1120 1210 1145 1260
rect 1195 1210 1255 1260
rect 1305 1210 1325 1260
rect 1120 1160 1325 1210
rect 1120 1110 1140 1160
rect 1190 1115 1325 1160
rect 1190 1110 1255 1115
rect 1120 1065 1255 1110
rect 1305 1065 1325 1115
rect 1120 1060 1325 1065
rect 1120 1010 1140 1060
rect 1190 1015 1325 1060
rect 1190 1010 1255 1015
rect 1120 965 1255 1010
rect 1305 965 1325 1015
rect 1120 960 1325 965
rect 1120 910 1140 960
rect 1190 915 1325 960
rect 1190 910 1255 915
rect 1120 865 1255 910
rect 1305 865 1325 915
rect 1120 855 1325 865
rect 1120 805 1140 855
rect 1190 815 1325 855
rect 1190 805 1255 815
rect 1120 765 1255 805
rect 1305 765 1325 815
rect 1120 760 1325 765
rect 1230 745 1325 760
rect 1425 1260 1515 1280
rect 1425 1210 1445 1260
rect 1495 1210 1515 1260
rect 1425 1080 1515 1210
rect 1425 1030 1445 1080
rect 1495 1030 1515 1080
rect 1425 980 1515 1030
rect 1425 930 1445 980
rect 1495 930 1515 980
rect 1425 845 1515 930
rect 1615 1260 1705 1395
rect 1615 1210 1635 1260
rect 1685 1210 1705 1260
rect 1615 1115 1705 1210
rect 1615 1065 1635 1115
rect 1685 1065 1705 1115
rect 1615 975 1705 1065
rect 1615 925 1635 975
rect 1685 925 1705 975
rect 1615 905 1705 925
rect 1805 1260 1895 1280
rect 1805 1210 1825 1260
rect 1875 1210 1895 1260
rect 1805 1085 1895 1210
rect 1805 1035 1825 1085
rect 1875 1035 1895 1085
rect 1805 985 1895 1035
rect 1805 935 1825 985
rect 1875 935 1895 985
rect 1805 885 1895 935
rect 1805 845 1825 885
rect 1425 835 1825 845
rect 1875 835 1895 885
rect 1425 825 1895 835
rect 1425 775 1445 825
rect 1495 785 1895 825
rect 1495 775 1825 785
rect 1425 755 1825 775
rect 1805 735 1825 755
rect 1875 735 1895 785
rect 205 610 295 685
rect 205 560 225 610
rect 275 560 295 610
rect 205 540 295 560
rect 690 665 1725 685
rect 690 615 1255 665
rect 1305 615 1355 665
rect 1405 615 1455 665
rect 1505 615 1555 665
rect 1605 615 1655 665
rect 1705 615 1725 665
rect 690 595 1725 615
rect 690 390 780 595
rect 1805 525 1895 735
rect 930 505 1020 525
rect 930 455 950 505
rect 1000 455 1020 505
rect 930 435 1020 455
rect 1425 435 1895 525
rect 55 370 145 390
rect 55 320 75 370
rect 125 320 145 370
rect 55 175 145 320
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 245 370 780 390
rect 245 320 265 370
rect 315 320 710 370
rect 760 320 780 370
rect 245 300 780 320
rect 245 175 335 300
rect 245 125 265 175
rect 315 125 335 175
rect 245 105 335 125
rect 465 220 555 240
rect 465 170 485 220
rect 535 170 555 220
rect 465 45 555 170
rect 690 175 780 300
rect 690 125 710 175
rect 760 125 780 175
rect 690 105 780 125
rect 880 355 970 375
rect 880 305 900 355
rect 950 305 970 355
rect 1235 370 1325 390
rect 1235 340 1255 370
rect 880 175 970 305
rect 880 125 900 175
rect 950 125 970 175
rect 880 45 970 125
rect 1120 320 1255 340
rect 1305 320 1325 370
rect 1120 270 1140 320
rect 1190 270 1325 320
rect 1120 205 1325 270
rect 1120 155 1140 205
rect 1190 155 1255 205
rect 1305 155 1325 205
rect 1120 45 1325 155
rect 1425 370 1515 435
rect 1425 320 1445 370
rect 1495 320 1515 370
rect 1805 370 1895 435
rect 1425 205 1515 320
rect 1425 155 1445 205
rect 1495 155 1515 205
rect 1425 135 1515 155
rect 1615 345 1705 365
rect 1615 295 1635 345
rect 1685 295 1705 345
rect 1615 205 1705 295
rect 1615 155 1635 205
rect 1685 155 1705 205
rect 1615 45 1705 155
rect 1805 320 1825 370
rect 1875 320 1895 370
rect 1805 205 1895 320
rect 1805 155 1825 205
rect 1875 155 1895 205
rect 1805 135 1895 155
rect 0 -45 1950 45
<< labels >>
flabel metal1 s 120 1415 120 1415 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel nwell 55 600 55 600 8 FreeSans 400 180 0 0 vdd
flabel metal1 s 225 550 225 550 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 1455 470 1455 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 950 445 950 445 2 FreeSans 400 0 0 0 b
port 2 ne
<< properties >>
string FIXED_BBOX 0 0 1950 1440
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
<< end >>
