magic
tech scmos
timestamp 1591563829
<< metal1 >>
rect -23 -10 -19 -3
rect -16 -10 -12 -3
rect -9 -10 -5 -3
rect -2 -10 2 -3
rect 5 -10 9 -3
rect 12 -10 16 -3
rect 19 -10 23 -3
rect 26 -10 30 -3
rect 33 -10 37 -3
rect 40 -10 44 -3
rect 47 -10 51 -3
rect 54 -10 58 -3
rect 61 -10 65 -3
rect 68 -10 72 -3
rect 75 -10 79 -3
rect 82 -10 86 -3
rect 89 -10 93 -3
rect 96 -10 100 -3
rect 103 -10 107 -3
rect 110 -10 114 -3
rect 117 -6 121 166
rect 124 -10 128 -3
rect 131 -10 135 -3
rect 138 -10 142 -3
rect 145 -10 149 -3
rect 152 -10 156 -3
rect 159 -10 163 -3
rect 166 -10 170 -3
rect 173 -10 177 -3
rect 180 -10 184 -3
rect 187 -10 191 -3
rect 194 -10 198 -3
rect 201 -10 205 -3
<< metal2 >>
rect -24 155 -4 161
rect -22 148 -8 152
rect -22 141 -8 145
rect -22 134 -8 138
rect -22 127 -8 131
rect -22 120 -8 124
rect -22 113 -8 117
rect -22 106 -8 110
rect -22 99 -8 103
rect -22 92 -8 96
rect -22 85 -8 89
rect -25 76 -5 82
rect -22 69 -8 73
rect -22 62 -8 66
rect -22 55 -8 59
rect -22 48 -8 52
rect -22 41 -8 45
rect -22 34 -8 38
rect -22 27 -8 31
rect -22 20 -8 24
rect -22 13 -8 17
rect -22 6 -8 10
rect -23 -3 -3 3
use inv_c  inv_c_0 ~/projects/ula/mag
timestamp 1591543887
transform 1 0 119 0 1 0
box -1 0 29 81
use dff_d_v2  dff_d_v2_1
timestamp 1542931922
transform 1 0 0 0 -1 158
box -1 0 120 81
use nor2_c  nor2_c_0
timestamp 1543318314
transform 1 0 119 0 -1 158
box -1 0 50 81
use dff_d_v2  dff_d_v2_0
timestamp 1542931922
transform 1 0 0 0 1 0
box -1 0 120 81
use inv_b  inv_b_0 ~/projects/ula/mag
timestamp 1591543887
transform 1 0 217 0 -1 158
box -1 0 29 81
use inv_c  inv_c_1
timestamp 1591543887
transform 1 0 147 0 1 0
box -1 0 29 81
use inv_c  inv_c_2
timestamp 1591543887
transform -1 0 203 0 1 0
box -1 0 29 81
use inv_c  inv_c_3
timestamp 1591543887
transform 1 0 203 0 1 0
box -1 0 29 81
use nor2_c  nor2_c_1
timestamp 1543318314
transform 1 0 168 0 -1 158
box -1 0 50 81
use buf_c  buf_c_0
timestamp 1543573773
transform 1 0 230 0 1 0
box 0 0 51 81
use nand2_b  nand2_b_0 ~/projects/ula/mag
timestamp 1591563829
transform 1 0 245 0 -1 158
box -1 0 36 81
<< end >>
