magic
tech amic5n
timestamp 1608317706
<< poly2capcontact >>
rect 875 515 1405 625
<< poly2cap >>
rect 810 240 1470 900
<< polysilicon >>
rect 660 60 1620 1050
<< polycontact >>
rect 695 95 745 145
<< polycontact >>
rect 845 95 895 145
<< polycontact >>
rect 995 95 1045 145
<< polycontact >>
rect 1145 95 1195 145
<< polycontact >>
rect 1295 95 1345 145
<< polycontact >>
rect 1445 95 1495 145
<< metal1 >>
rect 720 2190 2850 2370
rect 1260 630 1410 810
rect 3480 180 3630 1500
rect 660 0 3630 180
<< labels >>
flabel metal1  2550 60 2550 60 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 1350 720 1350 720 2 FreeSans 400 0 0 0 n2x
port 2 ne
flabel metal1  750 2340 750 2340 2 FreeSans 400 0 0 0 vdd
port 3 ne
<< checkpaint >>
rect -10 -10 3640 2380
<< end >>
