`celldefine
module nwsx ();
  // empty
endmodule
`endcelldefine
