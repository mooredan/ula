* input impedance  
*
* this can be used to determine the input capacitance

.include cell.cir
.lib ../../device_models/AMI_C5N.lib TT

.param VDD_VAL=5.0
.csparam v_vdd = {VDD_VAL}
.param FREQ=10.0Meg
.param PER={1 / FREQ}

.param TT=50p
.param CA=1f
.param CB=1f
.param CZ=1f

* power supply
Vvdd vdd 0 DC VDD_VAL PWL( 0 0  1u 0  2u {VDD_VAL})
Vvss vss 0 DC 0

* input a
Va   a_s 0 DC 0 PWL (                  0      0 
+                    {3u + PER *  2}          0
+                    {3u + PER *  2 + TT}  {VDD_VAL}
+                    {3u + PER *  3}       {VDD_VAL} 
+                    {3u + PER *  3 + TT}     0
+                    {3u + PER *  5}          0
+                    {3u + PER *  5 + TT}  {VDD_VAL}
+                    {3u + PER *  6}       {VDD_VAL} 
+                    {3u + PER *  6 + TT}     0
+                    {3u + PER * 10}          0 
+                    {3u + PER * 10 + TT}  {VDD_VAL})
Ra_s a_s a 100
Ca   a   0 {CA} 


* input b
Vb   b_s 0 DC 0 PWL (                  0      0 
+                    {3u + PER *  4}          0
+                    {3u + PER *  4 + TT}  {VDD_VAL}
+                    {3u + PER *  8}       {VDD_VAL} 
+                    {3u + PER *  8 + TT}     0
+                    {3u + PER *  9}          0
+                    {3u + PER *  9 + TT}  {VDD_VAL}
+                    {3u + PER * 11}       {VDD_VAL} 
+                    {3u + PER * 11 + TT}     0
+                    {3u + PER * 12}          0
+                    {3u + PER * 12 + TT}  {VDD_VAL})

Rb_s b_s b 100
Cb   b   0 {CA} 

* DUT
Xdut z a b vdd vss xor2_a

* output load
Cz z 0 {CZ} 

.control

***********************************
* Do input capacitance measurement
***********************************
* let vol  = $&v_vdd * 0.20
* set vol  = "$&vol"

let vmid = $&v_vdd * 0.5
set vmid = "$&vmid"

alter ca 0
alter cb 0
alter cz 0

* alter vvdd  dc 5.0
alter vvdd  dc $&v_vdd
alter va    dc $vmid
alter vb    dc $vmid

let idx = 70
set idx = "$&idx"

***********************************
* set up and measure input pin a
***********************************
alter va ac 1.0

ac dec 10 1 100e6

let freq = real(frequency[$idx])
set freq = "$&freq"

let a_cap = '1.0 / (imag(v(a)[$idx] / i(va)[$idx]) * 2 * pi * real(frequency[$idx]))'
set a_cap = "$&a_cap"
echo incap: pin: a cap: $a_cap  freq: $freq

***********************************
* set up and measure input pin b
***********************************
alter va ac 0.0
alter vb ac 1.0

ac dec 10 1 100e6

let freq = real(frequency[$idx])
set freq = "$&freq"

let b_cap = '1.0 / (imag(v(b)[$idx] / i(vb)[$idx]) * 2 * pi * real(frequency[$idx]))'
set b_cap = "$&b_cap"
echo incap: pin: b cap: $b_cap  freq: $freq

quit 0

.endc

.end
