magic
tech amic5n
magscale 1 2
timestamp 1624239416
<< nwell >>
rect 1115 1100 2535 2990
<< ntransistor >>
rect 1825 190 1945 800
<< ptransistor >>
rect 1825 1400 1945 2690
<< nselect >>
rect 1355 0 2295 860
<< pselect >>
rect 1355 1340 2295 2880
<< ndiffusion >>
rect 1585 740 1825 800
rect 1585 640 1645 740
rect 1745 640 1825 740
rect 1585 350 1825 640
rect 1585 250 1645 350
rect 1745 250 1825 350
rect 1585 190 1825 250
rect 1945 740 2185 800
rect 1945 640 2025 740
rect 2125 640 2185 740
rect 1945 350 2185 640
rect 1945 250 2025 350
rect 2125 250 2185 350
rect 1945 190 2185 250
<< pdiffusion >>
rect 1585 2630 1825 2690
rect 1585 2530 1645 2630
rect 1745 2530 1825 2630
rect 1585 2430 1825 2530
rect 1585 2330 1645 2430
rect 1745 2330 1825 2430
rect 1585 2230 1825 2330
rect 1585 2130 1645 2230
rect 1745 2130 1825 2230
rect 1585 2030 1825 2130
rect 1585 1930 1645 2030
rect 1745 1930 1825 2030
rect 1585 1830 1825 1930
rect 1585 1730 1645 1830
rect 1745 1730 1825 1830
rect 1585 1630 1825 1730
rect 1585 1530 1645 1630
rect 1745 1530 1825 1630
rect 1585 1400 1825 1530
rect 1945 2630 2185 2690
rect 1945 2530 2025 2630
rect 2125 2530 2185 2630
rect 1945 2360 2185 2530
rect 1945 2260 2025 2360
rect 2125 2260 2185 2360
rect 1945 2160 2185 2260
rect 1945 2060 2025 2160
rect 2125 2060 2185 2160
rect 1945 1960 2185 2060
rect 1945 1860 2025 1960
rect 2125 1860 2185 1960
rect 1945 1760 2185 1860
rect 1945 1660 2025 1760
rect 2125 1660 2185 1760
rect 1945 1560 2185 1660
rect 1945 1460 2025 1560
rect 2125 1460 2185 1560
rect 1945 1400 2185 1460
<< ndcontact >>
rect 1645 640 1745 740
rect 1645 250 1745 350
rect 2025 640 2125 740
rect 2025 250 2125 350
<< pdcontact >>
rect 1645 2530 1745 2630
rect 1645 2330 1745 2430
rect 1645 2130 1745 2230
rect 1645 1930 1745 2030
rect 1645 1730 1745 1830
rect 1645 1530 1745 1630
rect 2025 2530 2125 2630
rect 2025 2260 2125 2360
rect 2025 2060 2125 2160
rect 2025 1860 2125 1960
rect 2025 1660 2125 1760
rect 2025 1460 2125 1560
<< polysilicon >>
rect 1825 2690 1945 2820
rect 1825 1260 1945 1400
rect 1605 1220 1945 1260
rect 1605 1120 1645 1220
rect 1745 1120 1945 1220
rect 1605 1080 1945 1120
rect 1825 800 1945 1080
rect 1825 60 1945 190
<< polycontact >>
rect 1645 1120 1745 1220
<< metal1 >>
rect 1375 2790 2275 2970
rect 1605 2630 1785 2790
rect 1605 2530 1645 2630
rect 1745 2530 1785 2630
rect 1605 2430 1785 2530
rect 1605 2330 1645 2430
rect 1745 2330 1785 2430
rect 1605 2230 1785 2330
rect 1605 2130 1645 2230
rect 1745 2130 1785 2230
rect 1605 2030 1785 2130
rect 1605 1930 1645 2030
rect 1745 1930 1785 2030
rect 1605 1830 1785 1930
rect 1605 1730 1645 1830
rect 1745 1730 1785 1830
rect 1605 1630 1785 1730
rect 1605 1530 1645 1630
rect 1745 1530 1785 1630
rect 1605 1490 1785 1530
rect 1985 2630 2165 2670
rect 1985 2530 2025 2630
rect 2125 2530 2165 2630
rect 1985 2360 2165 2530
rect 1985 2260 2025 2360
rect 2125 2260 2165 2360
rect 1985 2160 2165 2260
rect 1985 2060 2025 2160
rect 2125 2060 2165 2160
rect 1985 1960 2165 2060
rect 1985 1860 2025 1960
rect 2125 1860 2165 1960
rect 1985 1760 2165 1860
rect 1985 1660 2025 1760
rect 2125 1660 2165 1760
rect 1985 1560 2165 1660
rect 1985 1460 2025 1560
rect 2125 1460 2165 1560
rect 1605 1220 1785 1370
rect 1605 1120 1645 1220
rect 1745 1120 1785 1220
rect 1605 1080 1785 1120
rect 1605 740 1785 780
rect 1605 640 1645 740
rect 1745 640 1785 740
rect 1605 350 1785 640
rect 1605 250 1645 350
rect 1745 250 1785 350
rect 1605 90 1785 250
rect 1985 740 2165 1460
rect 1985 640 2025 740
rect 2125 640 2165 740
rect 1985 350 2165 640
rect 1985 250 2025 350
rect 2125 250 2165 350
rect 1985 210 2165 250
rect 1375 -90 2275 90
rect -90 -1230 90 -950
rect -90 -1330 -50 -1230
rect 50 -1330 90 -1230
rect -90 -1550 90 -1330
rect -90 -1650 -50 -1550
rect 50 -1650 90 -1550
rect -90 -1810 90 -1650
rect 210 -1230 390 -970
rect 210 -1330 250 -1230
rect 350 -1330 390 -1230
rect 210 -1550 390 -1330
rect 210 -1650 250 -1550
rect 350 -1650 390 -1550
rect 210 -1770 390 -1650
rect 1695 -1140 2560 -865
rect 1695 -1240 1845 -1140
rect 1945 -1240 2065 -1140
rect 2165 -1240 2560 -1140
rect 1695 -1360 2560 -1240
rect 1695 -1460 1845 -1360
rect 1945 -1460 2065 -1360
rect 2165 -1460 2560 -1360
rect 1695 -1775 2560 -1460
<< via1 >>
rect -50 -1330 50 -1230
rect -50 -1650 50 -1550
rect 250 -1330 350 -1230
rect 250 -1650 350 -1550
rect 1845 -1240 1945 -1140
rect 2065 -1240 2165 -1140
rect 1845 -1460 1945 -1360
rect 2065 -1460 2165 -1360
<< metal2 >>
rect -5570 5350 1010 5530
rect -5570 5030 1010 5210
rect -5530 4710 1010 4890
rect -5530 4390 1010 4570
rect -5530 4070 1010 4250
rect -5530 3750 1010 3930
rect -5530 3430 1010 3610
rect -5530 3110 1010 3290
rect -5530 2790 1010 2970
rect -5530 2470 1010 2650
rect -5530 2150 1010 2330
rect -5530 1830 1010 2010
rect -5530 1510 1010 1690
rect -5530 1190 1010 1370
rect -5530 870 1010 1050
rect -5530 550 1010 730
rect -5530 230 1010 410
rect -5530 -90 1010 90
rect -5530 -410 1010 -230
rect -5530 -730 1010 -550
rect -5530 -1050 1010 -870
rect 1415 -1140 4660 -965
rect -1270 -1230 890 -1190
rect -1270 -1330 -1080 -1230
rect -980 -1330 -760 -1230
rect -660 -1330 -50 -1230
rect 50 -1330 250 -1230
rect 350 -1330 890 -1230
rect -1270 -1370 890 -1330
rect 1415 -1240 1845 -1140
rect 1945 -1240 2065 -1140
rect 2165 -1240 3340 -1140
rect 3440 -1145 4660 -1140
rect 3440 -1240 3600 -1145
rect 1415 -1245 3600 -1240
rect 3700 -1245 4660 -1145
rect 1415 -1360 4660 -1245
rect 1415 -1460 1845 -1360
rect 1945 -1460 2065 -1360
rect 2165 -1400 4660 -1360
rect 2165 -1460 3340 -1400
rect 1415 -1500 3340 -1460
rect 3440 -1405 4660 -1400
rect 3440 -1500 3600 -1405
rect 1415 -1505 3600 -1500
rect 3700 -1505 4660 -1405
rect -1270 -1550 890 -1510
rect -1270 -1650 -1080 -1550
rect -980 -1650 -760 -1550
rect -660 -1650 -50 -1550
rect 50 -1650 250 -1550
rect 350 -1650 890 -1550
rect 1415 -1645 4660 -1505
rect -1270 -1690 890 -1650
<< via2 >>
rect -1080 -1330 -980 -1230
rect -760 -1330 -660 -1230
rect 3340 -1240 3440 -1140
rect 3600 -1245 3700 -1145
rect 3340 -1500 3440 -1400
rect 3600 -1505 3700 -1405
rect -1080 -1650 -980 -1550
rect -760 -1650 -660 -1550
<< metal3 >>
rect -1110 -1190 -950 -1050
rect -790 -1190 -630 -1050
rect 3115 -1140 4065 -675
rect -1120 -1230 -940 -1190
rect -1120 -1330 -1080 -1230
rect -980 -1330 -940 -1230
rect -1120 -1370 -940 -1330
rect -800 -1230 -620 -1190
rect -800 -1330 -760 -1230
rect -660 -1330 -620 -1230
rect -800 -1370 -620 -1330
rect 3115 -1240 3340 -1140
rect 3440 -1145 4065 -1140
rect 3440 -1240 3600 -1145
rect 3115 -1245 3600 -1240
rect 3700 -1245 4065 -1145
rect -1110 -1510 -950 -1370
rect -790 -1510 -630 -1370
rect 3115 -1400 4065 -1245
rect 3115 -1500 3340 -1400
rect 3440 -1405 4065 -1400
rect 3440 -1500 3600 -1405
rect 3115 -1505 3600 -1500
rect 3700 -1505 4065 -1405
rect -1120 -1550 -940 -1510
rect -1120 -1650 -1080 -1550
rect -980 -1650 -940 -1550
rect -1120 -1690 -940 -1650
rect -800 -1550 -620 -1510
rect -800 -1650 -760 -1550
rect -660 -1650 -620 -1550
rect -800 -1690 -620 -1650
rect -1110 -1810 -950 -1690
rect -790 -1810 -630 -1690
rect 3115 -1810 4065 -1505
<< labels >>
flabel metal1 s 1565 2830 1565 2830 2 FreeSans 800 0 0 0 vdd
port 2 ne
flabel nwell 2165 1200 2165 1200 2 FreeSans 800 0 0 0 vdd
flabel metal1 s 2045 940 2045 940 2 FreeSans 800 0 0 0 z
port 0 ne
flabel metal1 s 1645 1100 1645 1100 2 FreeSans 800 0 0 0 a
port 1 ne
flabel metal1 s 1385 10 1385 10 2 FreeSans 800 0 0 0 vss
port 3 ne
<< end >>
