magic
tech amic5n
timestamp 1608317707
<< nwell >>
rect -120 870 1320 2430
<< nselect >>
rect 0 60 1200 750
<< pselect >>
rect 0 990 1200 2310
rect 210 960 270 990
rect 930 960 990 990
<< ntransistor >>
rect 210 120 270 690
rect 450 120 510 690
rect 690 120 750 690
rect 930 120 990 690
<< ptransistor >>
rect 210 1050 270 2250
rect 450 1050 510 2250
rect 690 1050 750 2250
rect 930 1050 990 2250
<< ndiffusion >>
rect 60 120 210 690
rect 270 120 450 690
rect 510 120 690 690
rect 750 120 930 690
rect 990 120 1140 690
<< pdiffusion >>
rect 60 1050 210 2250
rect 270 1050 450 2250
rect 510 1050 690 2250
rect 750 1050 930 2250
rect 990 1050 1140 2250
<< polysilicon >>
rect 210 2250 270 2310
rect 450 2250 510 2310
rect 690 2250 750 2310
rect 930 2250 990 2310
rect 210 960 270 1050
rect 60 780 270 960
rect 210 690 270 780
rect 450 960 510 1050
rect 690 960 750 1050
rect 450 780 750 960
rect 450 690 510 780
rect 690 690 750 780
rect 930 960 990 1050
rect 930 780 1140 960
rect 930 690 990 780
rect 210 60 270 120
rect 450 60 510 120
rect 690 60 750 120
rect 930 60 990 120
<< pdcontact >>
rect 95 2165 145 2215
<< pdcontact >>
rect 1055 2165 1105 2215
<< pdcontact >>
rect 335 2105 385 2155
<< pdcontact >>
rect 575 2105 625 2155
<< pdcontact >>
rect 815 2105 865 2155
<< pdcontact >>
rect 95 1985 145 2035
<< pdcontact >>
rect 335 1955 385 2005
<< pdcontact >>
rect 575 1955 625 2005
<< pdcontact >>
rect 815 1955 865 2005
<< pdcontact >>
rect 1055 1985 1105 2035
<< pdcontact >>
rect 95 1835 145 1885
<< pdcontact >>
rect 1055 1835 1105 1885
<< pdcontact >>
rect 335 1775 385 1825
<< pdcontact >>
rect 575 1775 625 1825
<< pdcontact >>
rect 815 1775 865 1825
<< pdcontact >>
rect 95 1685 145 1735
<< pdcontact >>
rect 1055 1685 1105 1735
<< pdcontact >>
rect 95 1535 145 1585
<< pdcontact >>
rect 335 1565 385 1615
<< pdcontact >>
rect 575 1595 625 1645
<< pdcontact >>
rect 815 1565 865 1615
<< pdcontact >>
rect 1055 1535 1105 1585
<< pdcontact >>
rect 95 1385 145 1435
<< pdcontact >>
rect 335 1385 385 1435
<< pdcontact >>
rect 575 1415 625 1465
<< pdcontact >>
rect 815 1385 865 1435
<< pdcontact >>
rect 1055 1385 1105 1435
<< pdcontact >>
rect 95 1235 145 1285
<< pdcontact >>
rect 335 1235 385 1285
<< pdcontact >>
rect 575 1235 625 1285
<< pdcontact >>
rect 815 1235 865 1285
<< pdcontact >>
rect 1055 1235 1105 1285
<< pdcontact >>
rect 95 1085 145 1135
<< pdcontact >>
rect 335 1085 385 1135
<< pdcontact >>
rect 575 1085 625 1135
<< pdcontact >>
rect 815 1085 865 1135
<< pdcontact >>
rect 1055 1085 1105 1135
<< polycontact >>
rect 125 845 175 895
<< polycontact >>
rect 575 845 625 895
<< polycontact >>
rect 1025 845 1075 895
<< ndcontact >>
rect 95 605 145 655
<< ndcontact >>
rect 575 605 625 655
<< ndcontact >>
rect 1055 605 1105 655
<< ndcontact >>
rect 95 455 145 505
<< ndcontact >>
rect 575 425 625 475
<< ndcontact >>
rect 1055 455 1105 505
<< ndcontact >>
rect 95 305 145 355
<< ndcontact >>
rect 1055 305 1105 355
<< ndcontact >>
rect 575 215 625 265
<< ndcontact >>
rect 95 155 145 205
<< ndcontact >>
rect 1055 155 1105 205
<< metal1 >>
rect 0 2280 1200 2370
rect 60 1050 180 2280
rect 90 810 210 930
rect 300 690 420 2190
rect 540 1050 660 2280
rect 510 810 690 930
rect 780 690 900 2190
rect 1020 1050 1140 2280
rect 990 810 1110 930
rect 60 90 180 690
rect 300 570 900 690
rect 540 180 660 570
rect 1020 90 1140 690
rect 0 0 1200 90
<< metal2 >>
rect 90 690 210 930
rect 540 810 660 1170
rect 990 690 1110 930
rect 90 570 1110 690
<< via1 >>
rect 125 845 175 895
rect 575 845 625 895
rect 1025 845 1075 895
<< labels >>
flabel nwell  0 930 0 930 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 30 30 30 30 2 FreeSans 400 0 0 0 vss
port 5 ne
flabel metal1 s 30 2310 30 2310 2 FreeSans 400 0 0 0 vdd
port 4 ne
flabel metal1 s 630 870 630 870 8 FreeSans 400 0 0 0 b
port 3 ne
flabel metal1 s 150 870 150 870 2 FreeSans 400 0 0 0 a
port 2 ne
flabel metal1 s 360 780 360 780 2 FreeSans 400 0 0 0 z
port 1 ne
flabel ndiffusion s 360 330 360 330 2 FreeSans 400 0 0 0 x1
flabel ndiffusion s 810 330 810 330 2 FreeSans 400 0 0 0 x2
<< checkpaint >>
rect -130 -10 1330 2440
<< end >>
