magic
tech amic5n
timestamp 1624419743
<< nwell >>
rect -130 550 1630 1495
<< ntransistor >>
rect 225 275 285 400
rect 615 95 675 400
rect 825 95 885 400
rect 1215 275 1275 400
<< ptransistor >>
rect 225 745 285 930
rect 615 700 675 1345
rect 825 700 885 1345
rect 1215 745 1275 930
<< nselect >>
rect 110 1090 320 1300
rect 1130 1040 1390 1300
rect -10 0 1510 430
<< pselect >>
rect -10 1300 1510 1440
rect -10 1090 110 1300
rect 320 1090 1130 1300
rect -10 1040 1130 1090
rect 1390 1040 1510 1300
rect -10 670 1510 1040
<< ndiffusion >>
rect 75 370 225 400
rect 75 320 115 370
rect 165 320 225 370
rect 75 275 225 320
rect 285 370 405 400
rect 285 320 325 370
rect 375 320 405 370
rect 285 275 405 320
rect 495 370 615 400
rect 495 320 525 370
rect 575 320 615 370
rect 75 270 195 275
rect 75 220 115 270
rect 165 220 195 270
rect 75 190 195 220
rect 495 175 615 320
rect 495 125 525 175
rect 575 125 615 175
rect 495 95 615 125
rect 675 95 825 400
rect 885 345 1005 400
rect 885 295 925 345
rect 975 295 1005 345
rect 885 185 1005 295
rect 1095 370 1215 400
rect 1095 320 1125 370
rect 1175 320 1215 370
rect 1095 275 1215 320
rect 1275 370 1425 400
rect 1275 320 1335 370
rect 1385 320 1425 370
rect 1275 275 1425 320
rect 1305 270 1425 275
rect 1305 220 1335 270
rect 1385 220 1425 270
rect 1305 190 1425 220
rect 885 135 925 185
rect 975 135 1005 185
rect 885 95 1005 135
<< pdiffusion >>
rect 495 1315 615 1345
rect 495 1265 525 1315
rect 575 1265 615 1315
rect 495 1215 615 1265
rect 495 1165 525 1215
rect 575 1165 615 1215
rect 495 1115 615 1165
rect 495 1065 525 1115
rect 575 1065 615 1115
rect 495 1015 615 1065
rect 75 930 195 955
rect 495 965 525 1015
rect 575 965 615 1015
rect 75 925 225 930
rect 75 875 115 925
rect 165 875 225 925
rect 75 825 225 875
rect 75 775 115 825
rect 165 775 225 825
rect 75 745 225 775
rect 285 860 405 930
rect 285 810 325 860
rect 375 810 405 860
rect 285 745 405 810
rect 495 900 615 965
rect 495 850 525 900
rect 575 850 615 900
rect 495 780 615 850
rect 495 730 525 780
rect 575 730 615 780
rect 495 700 615 730
rect 675 1315 825 1345
rect 675 1265 725 1315
rect 775 1265 825 1315
rect 675 1180 825 1265
rect 675 1130 725 1180
rect 775 1130 825 1180
rect 675 1080 825 1130
rect 675 1030 725 1080
rect 775 1030 825 1080
rect 675 980 825 1030
rect 675 930 725 980
rect 775 930 825 980
rect 675 880 825 930
rect 675 830 725 880
rect 775 830 825 880
rect 675 780 825 830
rect 675 730 725 780
rect 775 730 825 780
rect 675 700 825 730
rect 885 1315 1005 1345
rect 885 1265 925 1315
rect 975 1265 1005 1315
rect 885 1215 1005 1265
rect 885 1165 925 1215
rect 975 1165 1005 1215
rect 885 1115 1005 1165
rect 885 1065 925 1115
rect 975 1065 1005 1115
rect 885 1015 1005 1065
rect 885 965 925 1015
rect 975 965 1005 1015
rect 885 915 1005 965
rect 1305 930 1425 955
rect 885 865 925 915
rect 975 865 1005 915
rect 885 780 1005 865
rect 885 730 925 780
rect 975 730 1005 780
rect 1095 860 1215 930
rect 1095 810 1125 860
rect 1175 810 1215 860
rect 1095 745 1215 810
rect 1275 925 1425 930
rect 1275 875 1335 925
rect 1385 875 1425 925
rect 1275 825 1425 875
rect 1275 775 1335 825
rect 1385 775 1425 825
rect 1275 745 1425 775
rect 885 700 1005 730
<< nsubstratendiff >>
rect 140 1225 280 1255
rect 140 1175 185 1225
rect 235 1175 280 1225
rect 140 1145 280 1175
rect 1170 1225 1360 1255
rect 1170 1175 1265 1225
rect 1315 1175 1360 1225
rect 1170 1095 1360 1175
<< nsubstratencontact >>
rect 185 1175 235 1225
rect 1265 1175 1315 1225
<< ndcontact >>
rect 115 320 165 370
rect 325 320 375 370
rect 525 320 575 370
rect 115 220 165 270
rect 525 125 575 175
rect 925 295 975 345
rect 1125 320 1175 370
rect 1335 320 1385 370
rect 1335 220 1385 270
rect 925 135 975 185
<< pdcontact >>
rect 525 1265 575 1315
rect 525 1165 575 1215
rect 525 1065 575 1115
rect 525 965 575 1015
rect 115 875 165 925
rect 115 775 165 825
rect 325 810 375 860
rect 525 850 575 900
rect 525 730 575 780
rect 725 1265 775 1315
rect 725 1130 775 1180
rect 725 1030 775 1080
rect 725 930 775 980
rect 725 830 775 880
rect 725 730 775 780
rect 925 1265 975 1315
rect 925 1165 975 1215
rect 925 1065 975 1115
rect 925 965 975 1015
rect 925 865 975 915
rect 925 730 975 780
rect 1125 810 1175 860
rect 1335 875 1385 925
rect 1335 775 1385 825
<< polysilicon >>
rect 615 1345 675 1410
rect 825 1345 885 1410
rect 225 930 285 995
rect 225 685 285 745
rect 1215 930 1275 995
rect 115 665 285 685
rect 115 615 135 665
rect 185 615 285 665
rect 615 630 675 700
rect 115 595 285 615
rect 225 400 285 595
rect 490 610 675 630
rect 490 560 510 610
rect 560 560 675 610
rect 490 540 675 560
rect 615 400 675 540
rect 825 525 885 700
rect 1215 685 1275 745
rect 1215 665 1385 685
rect 1215 615 1315 665
rect 1365 615 1385 665
rect 1215 595 1385 615
rect 825 505 1010 525
rect 825 455 940 505
rect 990 455 1010 505
rect 825 435 1010 455
rect 825 400 885 435
rect 1215 400 1275 595
rect 225 210 285 275
rect 1215 210 1275 275
rect 615 30 675 95
rect 825 30 885 95
<< polycontact >>
rect 135 615 185 665
rect 510 560 560 610
rect 1315 615 1365 665
rect 940 455 990 505
<< metal1 >>
rect 0 1395 1500 1485
rect 95 1245 185 1395
rect 505 1315 595 1395
rect 505 1265 525 1315
rect 575 1265 595 1315
rect 95 1225 255 1245
rect 95 1175 185 1225
rect 235 1175 255 1225
rect 95 1155 255 1175
rect 505 1215 595 1265
rect 505 1165 525 1215
rect 575 1165 595 1215
rect 95 925 185 1155
rect 95 875 115 925
rect 165 875 185 925
rect 505 1115 595 1165
rect 505 1065 525 1115
rect 575 1065 595 1115
rect 505 1015 595 1065
rect 505 965 525 1015
rect 575 965 595 1015
rect 505 900 595 965
rect 95 825 185 875
rect 95 775 115 825
rect 165 775 185 825
rect 95 745 185 775
rect 305 860 395 890
rect 305 810 325 860
rect 375 810 395 860
rect 30 665 205 685
rect 30 615 135 665
rect 185 615 205 665
rect 30 595 205 615
rect 305 630 395 810
rect 505 850 525 900
rect 575 850 595 900
rect 505 780 595 850
rect 505 730 525 780
rect 575 730 595 780
rect 505 710 595 730
rect 705 1315 795 1335
rect 705 1265 725 1315
rect 775 1265 795 1315
rect 705 1180 795 1265
rect 705 1130 725 1180
rect 775 1130 795 1180
rect 705 1080 795 1130
rect 705 1030 725 1080
rect 775 1030 795 1080
rect 705 980 795 1030
rect 705 930 725 980
rect 775 930 795 980
rect 705 880 795 930
rect 705 830 725 880
rect 775 830 795 880
rect 705 780 795 830
rect 705 730 725 780
rect 775 730 795 780
rect 305 610 580 630
rect 305 560 510 610
rect 560 560 580 610
rect 305 540 580 560
rect 95 370 185 390
rect 95 320 115 370
rect 165 320 185 370
rect 95 270 185 320
rect 305 370 395 540
rect 305 320 325 370
rect 375 320 395 370
rect 305 285 395 320
rect 505 370 595 390
rect 505 320 525 370
rect 575 320 595 370
rect 95 220 115 270
rect 165 220 185 270
rect 95 45 185 220
rect 505 175 595 320
rect 705 365 795 730
rect 905 1315 995 1395
rect 905 1265 925 1315
rect 975 1265 995 1315
rect 905 1215 995 1265
rect 1315 1245 1405 1395
rect 905 1165 925 1215
rect 975 1165 995 1215
rect 905 1115 995 1165
rect 1245 1225 1405 1245
rect 1245 1175 1265 1225
rect 1315 1175 1405 1225
rect 1245 1155 1405 1175
rect 905 1065 925 1115
rect 975 1065 995 1115
rect 905 1015 995 1065
rect 905 965 925 1015
rect 975 965 995 1015
rect 905 915 995 965
rect 905 865 925 915
rect 975 865 995 915
rect 1315 925 1405 1155
rect 905 780 995 865
rect 905 730 925 780
rect 975 730 995 780
rect 905 710 995 730
rect 1105 860 1195 890
rect 1105 810 1125 860
rect 1175 810 1195 860
rect 1105 525 1195 810
rect 1315 875 1335 925
rect 1385 875 1405 925
rect 1315 825 1405 875
rect 1315 775 1335 825
rect 1385 775 1405 825
rect 1315 745 1405 775
rect 1295 665 1470 685
rect 1295 615 1315 665
rect 1365 615 1470 665
rect 1295 595 1470 615
rect 920 505 1195 525
rect 920 455 940 505
rect 990 455 1195 505
rect 920 435 1195 455
rect 1105 370 1195 435
rect 705 345 995 365
rect 705 295 925 345
rect 975 295 995 345
rect 705 275 995 295
rect 1105 320 1125 370
rect 1175 320 1195 370
rect 1105 285 1195 320
rect 1315 370 1405 390
rect 1315 320 1335 370
rect 1385 320 1405 370
rect 505 125 525 175
rect 575 125 595 175
rect 505 45 595 125
rect 905 185 995 275
rect 905 135 925 185
rect 975 135 995 185
rect 905 105 995 135
rect 1315 270 1405 320
rect 1315 220 1335 270
rect 1385 220 1405 270
rect 1315 45 1405 220
rect 0 -45 1500 45
<< labels >>
flabel metal1 s 735 470 735 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 50 615 50 615 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 1426 620 1426 620 2 FreeSans 400 0 0 0 b
port 2 ne
flabel metal1 s 206 1415 206 1415 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 6 5 6 5 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel nwell 30 555 30 555 2 FreeSans 400 0 0 0 vdd
<< properties >>
string FIXED_BBOX 0 0 1500 1440
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
