magic
tech amic5n
timestamp 1625354305
<< nwell >>
rect -130 550 730 1495
<< ntransistor >>
rect 165 95 435 400
<< ptransistor >>
rect 165 710 435 1345
<< nselect >>
rect -10 0 610 430
<< pselect >>
rect -10 680 610 1440
rect -10 670 165 680
rect 435 670 610 680
<< ndiffusion >>
rect 45 370 165 400
rect 45 320 75 370
rect 125 320 165 370
rect 45 175 165 320
rect 45 125 75 175
rect 125 125 165 175
rect 45 95 165 125
rect 435 355 555 400
rect 435 305 475 355
rect 525 305 555 355
rect 435 175 555 305
rect 435 125 475 175
rect 525 125 555 175
rect 435 95 555 125
<< pdiffusion >>
rect 45 1315 165 1345
rect 45 1265 75 1315
rect 125 1265 165 1315
rect 45 1190 165 1265
rect 45 1140 75 1190
rect 125 1140 165 1190
rect 45 1090 165 1140
rect 45 1040 75 1090
rect 125 1040 165 1090
rect 45 990 165 1040
rect 45 940 75 990
rect 125 940 165 990
rect 45 890 165 940
rect 45 840 75 890
rect 125 840 165 890
rect 45 710 165 840
rect 435 1315 555 1345
rect 435 1265 475 1315
rect 525 1265 555 1315
rect 435 1190 555 1265
rect 435 1140 475 1190
rect 525 1140 555 1190
rect 435 1090 555 1140
rect 435 1040 475 1090
rect 525 1040 555 1090
rect 435 990 555 1040
rect 435 940 475 990
rect 525 940 555 990
rect 435 890 555 940
rect 435 840 475 890
rect 525 840 555 890
rect 435 790 555 840
rect 435 740 475 790
rect 525 740 555 790
rect 435 710 555 740
<< ndcontact >>
rect 75 320 125 370
rect 75 125 125 175
rect 475 305 525 355
rect 475 125 525 175
<< pdcontact >>
rect 75 1265 125 1315
rect 75 1140 125 1190
rect 75 1040 125 1090
rect 75 940 125 990
rect 75 840 125 890
rect 475 1265 525 1315
rect 475 1140 525 1190
rect 475 1040 525 1090
rect 475 940 525 990
rect 475 840 525 890
rect 475 740 525 790
<< polysilicon >>
rect 165 1345 435 1410
rect 165 675 435 710
rect 105 655 435 675
rect 105 605 125 655
rect 175 605 225 655
rect 275 605 325 655
rect 375 605 435 655
rect 105 585 435 605
rect 165 505 495 525
rect 165 455 225 505
rect 275 455 325 505
rect 375 455 425 505
rect 475 455 495 505
rect 165 435 495 455
rect 165 400 435 435
rect 165 30 435 95
<< polycontact >>
rect 125 605 175 655
rect 225 605 275 655
rect 325 605 375 655
rect 225 455 275 505
rect 325 455 375 505
rect 425 455 475 505
<< metal1 >>
rect 0 1395 600 1485
rect 55 1315 145 1395
rect 55 1265 75 1315
rect 125 1265 145 1315
rect 55 1190 145 1265
rect 55 1140 75 1190
rect 125 1140 145 1190
rect 55 1090 145 1140
rect 55 1040 75 1090
rect 125 1040 145 1090
rect 55 990 145 1040
rect 55 940 75 990
rect 125 940 145 990
rect 55 890 145 940
rect 55 840 75 890
rect 125 840 145 890
rect 55 735 145 840
rect 205 675 395 1335
rect 55 655 395 675
rect 55 605 125 655
rect 175 605 225 655
rect 275 605 325 655
rect 375 605 395 655
rect 55 585 395 605
rect 455 1315 545 1395
rect 455 1265 475 1315
rect 525 1265 545 1315
rect 455 1190 545 1265
rect 455 1140 475 1190
rect 525 1140 545 1190
rect 455 1090 545 1140
rect 455 1040 475 1090
rect 525 1040 545 1090
rect 455 990 545 1040
rect 455 940 475 990
rect 525 940 545 990
rect 455 890 545 940
rect 455 840 475 890
rect 525 840 545 890
rect 455 790 545 840
rect 455 740 475 790
rect 525 740 545 790
rect 55 370 145 585
rect 455 525 545 740
rect 55 320 75 370
rect 125 320 145 370
rect 55 175 145 320
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 205 505 545 525
rect 205 455 225 505
rect 275 455 325 505
rect 375 455 425 505
rect 475 455 545 505
rect 205 435 545 455
rect 205 105 395 435
rect 455 355 545 375
rect 455 305 475 355
rect 525 305 545 355
rect 455 175 545 305
rect 455 125 475 175
rect 525 125 545 175
rect 455 45 545 125
rect 0 -45 600 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 1 ne
flabel metal1 s 20 1415 20 1415 2 FreeSans 400 0 0 0 vdd
port 0 ne
flabel nwell 5 600 5 600 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFclass CORE
string LEFsite core
string FIXED_BBOX 0 0 600 1440
string LEFsymmetry X Y
<< end >>
