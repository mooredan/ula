module fill2 ();
endmodule
