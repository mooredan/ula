magic
tech scmos
timestamp 1607032420
<< poly2capcontact >>
rect 935 1835 2245 1945
<< poly2capcontact >>
rect 3095 1835 3985 1945
<< poly2capcontact >>
rect 875 515 1405 625
<< poly2cap >>
rect 870 1650 2310 2130
rect 3030 1650 4050 2130
rect 810 240 1470 900
<< psubstratepdiff >>
rect 2370 390 2730 690
<< polysilicon >>
rect 720 1500 2460 2310
rect 2850 1500 4200 2310
rect 660 60 1620 1050
<< polycontact >>
rect 755 2225 805 2275
<< polycontact >>
rect 905 2225 955 2275
<< polycontact >>
rect 1055 2225 1105 2275
<< polycontact >>
rect 1205 2225 1255 2275
<< polycontact >>
rect 1355 2225 1405 2275
<< polycontact >>
rect 1535 2225 1585 2275
<< polycontact >>
rect 1685 2225 1735 2275
<< polycontact >>
rect 1835 2225 1885 2275
<< polycontact >>
rect 1985 2225 2035 2275
<< polycontact >>
rect 2135 2225 2185 2275
<< polycontact >>
rect 2285 2225 2335 2275
<< polycontact >>
rect 3095 2225 3145 2275
<< polycontact >>
rect 3275 2225 3325 2275
<< polycontact >>
rect 3425 2225 3475 2275
<< polycontact >>
rect 3575 2225 3625 2275
<< polycontact >>
rect 3725 2225 3775 2275
<< polycontact >>
rect 3875 2225 3925 2275
<< polycontact >>
rect 4025 2225 4075 2275
<< psubstratepcontact >>
rect 2525 515 2575 565
<< polycontact >>
rect 695 95 745 145
<< polycontact >>
rect 845 95 895 145
<< polycontact >>
rect 995 95 1045 145
<< polycontact >>
rect 1145 95 1195 145
<< polycontact >>
rect 1295 95 1345 145
<< polycontact >>
rect 1445 95 1495 145
<< metal1 >>
rect 720 2190 4200 2370
rect 2100 1650 2250 1830
rect 1260 630 1410 810
rect 2490 180 2610 600
rect 3480 180 3630 1830
rect 660 0 3630 180
<< labels >>
flabel metal1 s 2160 1710 2160 1710 2 FreeSans 400 0 0 0 n2
port 1 ne
flabel metal1  750 2340 750 2340 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1  2550 60 2550 60 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 1350 720 1350 720 2 FreeSans 400 0 0 0 n2x
port 2 ne
<< checkpaint >>
rect -10 -10 4210 2380
<< end >>
