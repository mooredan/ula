magic
tech amic5n
timestamp 1608317706
<< nwell >>
rect 0 870 810 2370
<< poly2 >>
rect 780 1200 930 1350
rect 4020 1200 4200 1350
