magic
tech scmos
magscale 1 2
timestamp 1570494029
<< error_p >>
rect 20 1320 22 1322
rect 578 1320 580 1322
rect 18 1318 20 1320
rect 580 1318 582 1320
rect 80 1296 90 1298
rect 78 1294 90 1296
rect 510 1296 520 1298
rect 510 1294 522 1296
rect 80 1290 82 1294
rect 518 1290 520 1294
rect 80 1286 90 1290
rect 78 1284 90 1286
rect 510 1286 520 1290
rect 510 1284 522 1286
rect 80 1282 82 1284
rect 518 1282 520 1284
rect 82 1280 84 1282
rect 516 1280 518 1282
rect 50 1279 52 1280
rect 548 1279 550 1280
rect 48 1277 50 1278
rect 550 1277 552 1278
rect 50 1259 52 1260
rect 548 1259 550 1260
rect 48 1257 50 1258
rect 550 1257 552 1258
rect 96 1242 98 1244
rect 502 1242 504 1244
rect 94 1240 96 1242
rect 504 1240 506 1242
rect 50 1239 52 1240
rect 548 1239 550 1240
rect 48 1237 50 1238
rect 550 1237 552 1238
rect 50 1219 52 1220
rect 548 1219 550 1220
rect 48 1217 50 1218
rect 550 1217 552 1218
rect 50 1199 52 1200
rect 548 1199 550 1200
rect 48 1197 50 1198
rect 550 1197 552 1198
rect 94 1180 96 1182
rect 504 1180 506 1182
rect 50 1179 52 1180
rect 96 1178 98 1180
rect 502 1178 504 1180
rect 548 1179 550 1180
rect 48 1177 50 1178
rect 550 1177 552 1178
rect 50 1159 52 1160
rect 548 1159 550 1160
rect 48 1157 50 1158
rect 550 1157 552 1158
rect 50 1139 52 1140
rect 548 1139 550 1140
rect 48 1137 50 1138
rect 550 1137 552 1138
rect 50 1119 52 1120
rect 548 1119 550 1120
rect 48 1117 50 1118
rect 550 1117 552 1118
rect 96 1114 98 1116
rect 502 1114 504 1116
rect 94 1112 96 1114
rect 504 1112 506 1114
rect 50 1099 52 1100
rect 548 1099 550 1100
rect 48 1097 50 1098
rect 550 1097 552 1098
rect 50 1079 52 1080
rect 548 1079 550 1080
rect 48 1077 50 1078
rect 550 1077 552 1078
rect 50 1059 52 1060
rect 548 1059 550 1060
rect 48 1057 50 1058
rect 550 1057 552 1058
rect 94 1052 96 1054
rect 504 1052 506 1054
rect 96 1050 98 1052
rect 502 1050 504 1052
rect 50 1039 52 1040
rect 548 1039 550 1040
rect 48 1037 50 1038
rect 550 1037 552 1038
rect 50 1019 52 1020
rect 548 1019 550 1020
rect 48 1017 50 1018
rect 550 1017 552 1018
rect 50 999 52 1000
rect 548 999 550 1000
rect 48 997 50 998
rect 550 997 552 998
rect 96 984 98 986
rect 502 984 504 986
rect 94 982 96 984
rect 504 982 506 984
rect 50 979 52 980
rect 548 979 550 980
rect 48 977 50 978
rect 550 977 552 978
rect 50 959 52 960
rect 548 959 550 960
rect 48 957 50 958
rect 550 957 552 958
rect 50 939 52 940
rect 548 939 550 940
rect 48 937 50 938
rect 550 937 552 938
rect 94 922 96 924
rect 504 922 506 924
rect 96 920 98 922
rect 502 920 504 922
rect 50 919 52 920
rect 548 919 550 920
rect 48 917 50 918
rect 550 917 552 918
rect 50 899 52 900
rect 548 899 550 900
rect 48 897 50 898
rect 550 897 552 898
rect 294 895 296 897
rect 304 895 306 897
rect 292 893 294 895
rect 306 893 308 895
rect 62 873 64 875
rect 536 873 538 875
rect 60 871 62 873
rect 538 871 540 873
rect 32 828 34 830
rect 62 828 64 830
rect 92 828 94 830
rect 122 828 124 830
rect 152 828 154 830
rect 182 828 184 830
rect 416 828 418 830
rect 446 828 448 830
rect 476 828 478 830
rect 506 828 508 830
rect 536 828 538 830
rect 566 828 568 830
rect 34 826 36 828
rect 40 826 42 828
rect 64 826 66 828
rect 70 826 72 828
rect 94 826 96 828
rect 100 826 102 828
rect 124 826 126 828
rect 130 826 132 828
rect 154 826 156 828
rect 160 826 162 828
rect 184 826 186 828
rect 414 826 416 828
rect 438 826 440 828
rect 444 826 446 828
rect 468 826 470 828
rect 474 826 476 828
rect 498 826 500 828
rect 504 826 506 828
rect 528 826 530 828
rect 534 826 536 828
rect 558 826 560 828
rect 564 826 566 828
rect 42 824 44 826
rect 72 824 74 826
rect 102 824 104 826
rect 132 824 134 826
rect 162 824 164 826
rect 436 824 438 826
rect 466 824 468 826
rect 496 824 498 826
rect 526 824 528 826
rect 556 824 558 826
rect 42 818 44 820
rect 72 818 74 820
rect 102 818 104 820
rect 132 818 134 820
rect 162 818 164 820
rect 436 818 438 820
rect 466 818 468 820
rect 496 818 498 820
rect 526 818 528 820
rect 556 818 558 820
rect 34 816 36 818
rect 40 816 42 818
rect 64 816 66 818
rect 70 816 72 818
rect 94 816 96 818
rect 100 816 102 818
rect 124 816 126 818
rect 130 816 132 818
rect 154 816 156 818
rect 160 816 162 818
rect 184 816 186 818
rect 414 816 416 818
rect 438 816 440 818
rect 444 816 446 818
rect 468 816 470 818
rect 474 816 476 818
rect 498 816 500 818
rect 504 816 506 818
rect 528 816 530 818
rect 534 816 536 818
rect 558 816 560 818
rect 564 816 566 818
rect 32 814 34 816
rect 62 814 64 816
rect 92 814 94 816
rect 122 814 124 816
rect 152 814 154 816
rect 182 814 184 816
rect 416 814 418 816
rect 446 814 448 816
rect 476 814 478 816
rect 506 814 508 816
rect 536 814 538 816
rect 566 814 568 816
rect 32 808 34 810
rect 62 808 64 810
rect 92 808 94 810
rect 122 808 124 810
rect 152 808 154 810
rect 182 808 184 810
rect 416 808 418 810
rect 446 808 448 810
rect 476 808 478 810
rect 506 808 508 810
rect 536 808 538 810
rect 566 808 568 810
rect 34 806 36 808
rect 40 806 42 808
rect 64 806 66 808
rect 70 806 72 808
rect 94 806 96 808
rect 100 806 102 808
rect 124 806 126 808
rect 130 806 132 808
rect 154 806 156 808
rect 160 806 162 808
rect 184 806 186 808
rect 414 806 416 808
rect 438 806 440 808
rect 444 806 446 808
rect 468 806 470 808
rect 474 806 476 808
rect 498 806 500 808
rect 504 806 506 808
rect 528 806 530 808
rect 534 806 536 808
rect 558 806 560 808
rect 564 806 566 808
rect 42 804 44 806
rect 72 804 74 806
rect 102 804 104 806
rect 132 804 134 806
rect 162 804 164 806
rect 436 804 438 806
rect 466 804 468 806
rect 496 804 498 806
rect 526 804 528 806
rect 556 804 558 806
rect 42 798 44 800
rect 72 798 74 800
rect 102 798 104 800
rect 132 798 134 800
rect 162 798 164 800
rect 436 798 438 800
rect 466 798 468 800
rect 496 798 498 800
rect 526 798 528 800
rect 556 798 558 800
rect 34 796 36 798
rect 40 796 42 798
rect 64 796 66 798
rect 70 796 72 798
rect 94 796 96 798
rect 100 796 102 798
rect 124 796 126 798
rect 130 796 132 798
rect 154 796 156 798
rect 160 796 162 798
rect 184 796 186 798
rect 414 796 416 798
rect 438 796 440 798
rect 444 796 446 798
rect 468 796 470 798
rect 474 796 476 798
rect 498 796 500 798
rect 504 796 506 798
rect 528 796 530 798
rect 534 796 536 798
rect 558 796 560 798
rect 564 796 566 798
rect 32 794 34 796
rect 62 794 64 796
rect 92 794 94 796
rect 122 794 124 796
rect 152 794 154 796
rect 182 794 184 796
rect 416 794 418 796
rect 446 794 448 796
rect 476 794 478 796
rect 506 794 508 796
rect 536 794 538 796
rect 566 794 568 796
rect 32 788 34 790
rect 62 788 64 790
rect 92 788 94 790
rect 122 788 124 790
rect 152 788 154 790
rect 182 788 184 790
rect 416 788 418 790
rect 446 788 448 790
rect 476 788 478 790
rect 506 788 508 790
rect 536 788 538 790
rect 566 788 568 790
rect 34 786 36 788
rect 40 786 42 788
rect 64 786 66 788
rect 70 786 72 788
rect 94 786 96 788
rect 100 786 102 788
rect 124 786 126 788
rect 130 786 132 788
rect 154 786 156 788
rect 160 786 162 788
rect 184 786 186 788
rect 414 786 416 788
rect 438 786 440 788
rect 444 786 446 788
rect 468 786 470 788
rect 474 786 476 788
rect 498 786 500 788
rect 504 786 506 788
rect 528 786 530 788
rect 534 786 536 788
rect 558 786 560 788
rect 564 786 566 788
rect 42 784 44 786
rect 72 784 74 786
rect 102 784 104 786
rect 132 784 134 786
rect 162 784 164 786
rect 436 784 438 786
rect 466 784 468 786
rect 496 784 498 786
rect 526 784 528 786
rect 556 784 558 786
rect 42 778 44 780
rect 72 778 74 780
rect 526 778 528 780
rect 556 778 558 780
rect 34 776 36 778
rect 40 776 42 778
rect 64 776 66 778
rect 70 776 72 778
rect 94 776 96 778
rect 110 776 112 778
rect 124 776 126 778
rect 140 776 142 778
rect 154 776 156 778
rect 170 776 172 778
rect 184 776 186 778
rect 414 776 416 778
rect 428 776 430 778
rect 444 776 446 778
rect 458 776 460 778
rect 474 776 476 778
rect 488 776 490 778
rect 504 776 506 778
rect 528 776 530 778
rect 534 776 536 778
rect 558 776 560 778
rect 564 776 566 778
rect 32 774 34 776
rect 62 774 64 776
rect 92 774 94 776
rect 112 774 114 776
rect 122 774 124 776
rect 142 774 144 776
rect 152 774 154 776
rect 172 774 174 776
rect 182 774 184 776
rect 416 774 418 776
rect 426 774 428 776
rect 446 774 448 776
rect 456 774 458 776
rect 476 774 478 776
rect 486 774 488 776
rect 506 774 508 776
rect 536 774 538 776
rect 566 774 568 776
rect 32 768 34 770
rect 62 768 64 770
rect 92 768 94 770
rect 112 768 114 770
rect 122 768 124 770
rect 142 768 144 770
rect 152 768 154 770
rect 172 768 174 770
rect 182 768 184 770
rect 416 768 418 770
rect 426 768 428 770
rect 446 768 448 770
rect 456 768 458 770
rect 476 768 478 770
rect 486 768 488 770
rect 506 768 508 770
rect 536 768 538 770
rect 566 768 568 770
rect 34 766 36 768
rect 40 766 42 768
rect 64 766 66 768
rect 70 766 72 768
rect 94 766 96 768
rect 110 766 112 768
rect 124 766 126 768
rect 140 766 142 768
rect 154 766 156 768
rect 170 766 172 768
rect 184 766 186 768
rect 414 766 416 768
rect 428 766 430 768
rect 444 766 446 768
rect 458 766 460 768
rect 474 766 476 768
rect 488 766 490 768
rect 504 766 506 768
rect 528 766 530 768
rect 534 766 536 768
rect 558 766 560 768
rect 564 766 566 768
rect 42 764 44 766
rect 72 764 74 766
rect 526 764 528 766
rect 556 764 558 766
rect 42 758 44 760
rect 72 758 74 760
rect 102 758 104 760
rect 132 758 134 760
rect 162 758 164 760
rect 436 758 438 760
rect 466 758 468 760
rect 496 758 498 760
rect 526 758 528 760
rect 556 758 558 760
rect 34 756 36 758
rect 40 756 42 758
rect 64 756 66 758
rect 70 756 72 758
rect 94 756 96 758
rect 100 756 102 758
rect 124 756 126 758
rect 130 756 132 758
rect 154 756 156 758
rect 160 756 162 758
rect 184 756 186 758
rect 414 756 416 758
rect 438 756 440 758
rect 444 756 446 758
rect 468 756 470 758
rect 474 756 476 758
rect 498 756 500 758
rect 504 756 506 758
rect 528 756 530 758
rect 534 756 536 758
rect 558 756 560 758
rect 564 756 566 758
rect 32 754 34 756
rect 62 754 64 756
rect 92 754 94 756
rect 122 754 124 756
rect 152 754 154 756
rect 182 754 184 756
rect 416 754 418 756
rect 446 754 448 756
rect 476 754 478 756
rect 506 754 508 756
rect 536 754 538 756
rect 566 754 568 756
rect 32 748 34 750
rect 62 748 64 750
rect 92 748 94 750
rect 122 748 124 750
rect 152 748 154 750
rect 182 748 184 750
rect 416 748 418 750
rect 446 748 448 750
rect 476 748 478 750
rect 506 748 508 750
rect 536 748 538 750
rect 566 748 568 750
rect 34 746 36 748
rect 40 746 42 748
rect 64 746 66 748
rect 70 746 72 748
rect 94 746 96 748
rect 100 746 102 748
rect 124 746 126 748
rect 130 746 132 748
rect 154 746 156 748
rect 160 746 162 748
rect 184 746 186 748
rect 414 746 416 748
rect 438 746 440 748
rect 444 746 446 748
rect 468 746 470 748
rect 474 746 476 748
rect 498 746 500 748
rect 504 746 506 748
rect 528 746 530 748
rect 534 746 536 748
rect 558 746 560 748
rect 564 746 566 748
rect 42 744 44 746
rect 72 744 74 746
rect 102 744 104 746
rect 132 744 134 746
rect 162 744 164 746
rect 436 744 438 746
rect 466 744 468 746
rect 496 744 498 746
rect 526 744 528 746
rect 556 744 558 746
rect 42 718 44 720
rect 72 718 74 720
rect 102 718 104 720
rect 132 718 134 720
rect 162 718 164 720
rect 436 718 438 720
rect 466 718 468 720
rect 496 718 498 720
rect 526 718 528 720
rect 556 718 558 720
rect 34 716 36 718
rect 40 716 42 718
rect 64 716 66 718
rect 70 716 72 718
rect 94 716 96 718
rect 100 716 102 718
rect 124 716 126 718
rect 130 716 132 718
rect 154 716 156 718
rect 160 716 162 718
rect 184 716 186 718
rect 414 716 416 718
rect 438 716 440 718
rect 444 716 446 718
rect 468 716 470 718
rect 474 716 476 718
rect 498 716 500 718
rect 504 716 506 718
rect 528 716 530 718
rect 534 716 536 718
rect 558 716 560 718
rect 564 716 566 718
rect 32 714 34 716
rect 62 714 64 716
rect 92 714 94 716
rect 122 714 124 716
rect 152 714 154 716
rect 182 714 184 716
rect 416 714 418 716
rect 446 714 448 716
rect 476 714 478 716
rect 506 714 508 716
rect 536 714 538 716
rect 566 714 568 716
rect 32 708 34 710
rect 62 708 64 710
rect 92 708 94 710
rect 122 708 124 710
rect 152 708 154 710
rect 182 708 184 710
rect 416 708 418 710
rect 446 708 448 710
rect 476 708 478 710
rect 506 708 508 710
rect 536 708 538 710
rect 566 708 568 710
rect 34 706 36 708
rect 40 706 42 708
rect 64 706 66 708
rect 70 706 72 708
rect 94 706 96 708
rect 100 706 102 708
rect 124 706 126 708
rect 130 706 132 708
rect 154 706 156 708
rect 160 706 162 708
rect 184 706 186 708
rect 414 706 416 708
rect 438 706 440 708
rect 444 706 446 708
rect 468 706 470 708
rect 474 706 476 708
rect 498 706 500 708
rect 504 706 506 708
rect 528 706 530 708
rect 534 706 536 708
rect 558 706 560 708
rect 564 706 566 708
rect 42 704 44 706
rect 72 704 74 706
rect 102 704 104 706
rect 132 704 134 706
rect 162 704 164 706
rect 436 704 438 706
rect 466 704 468 706
rect 496 704 498 706
rect 526 704 528 706
rect 556 704 558 706
rect 42 698 44 700
rect 72 698 74 700
rect 102 698 104 700
rect 132 698 134 700
rect 162 698 164 700
rect 436 698 438 700
rect 466 698 468 700
rect 496 698 498 700
rect 526 698 528 700
rect 556 698 558 700
rect 34 696 36 698
rect 40 696 42 698
rect 64 696 66 698
rect 70 696 72 698
rect 94 696 96 698
rect 100 696 102 698
rect 124 696 126 698
rect 130 696 132 698
rect 154 696 156 698
rect 160 696 162 698
rect 184 696 186 698
rect 414 696 416 698
rect 438 696 440 698
rect 444 696 446 698
rect 468 696 470 698
rect 474 696 476 698
rect 498 696 500 698
rect 504 696 506 698
rect 528 696 530 698
rect 534 696 536 698
rect 558 696 560 698
rect 564 696 566 698
rect 32 694 34 696
rect 62 694 64 696
rect 92 694 94 696
rect 122 694 124 696
rect 152 694 154 696
rect 182 694 184 696
rect 416 694 418 696
rect 446 694 448 696
rect 476 694 478 696
rect 506 694 508 696
rect 536 694 538 696
rect 566 694 568 696
rect 32 644 34 646
rect 62 644 64 646
rect 92 644 94 646
rect 122 644 124 646
rect 152 644 154 646
rect 182 644 184 646
rect 416 644 418 646
rect 446 644 448 646
rect 476 644 478 646
rect 506 644 508 646
rect 536 644 538 646
rect 566 644 568 646
rect 34 642 36 644
rect 40 642 42 644
rect 64 642 66 644
rect 70 642 72 644
rect 94 642 96 644
rect 100 642 102 644
rect 124 642 126 644
rect 130 642 132 644
rect 154 642 156 644
rect 160 642 162 644
rect 184 642 186 644
rect 414 642 416 644
rect 438 642 440 644
rect 444 642 446 644
rect 468 642 470 644
rect 474 642 476 644
rect 498 642 500 644
rect 504 642 506 644
rect 528 642 530 644
rect 534 642 536 644
rect 558 642 560 644
rect 564 642 566 644
rect 42 640 44 642
rect 72 640 74 642
rect 102 640 104 642
rect 132 640 134 642
rect 162 640 164 642
rect 436 640 438 642
rect 466 640 468 642
rect 496 640 498 642
rect 526 640 528 642
rect 556 640 558 642
rect 42 634 44 636
rect 72 634 74 636
rect 102 634 104 636
rect 132 634 134 636
rect 162 634 164 636
rect 436 634 438 636
rect 466 634 468 636
rect 496 634 498 636
rect 526 634 528 636
rect 556 634 558 636
rect 34 632 36 634
rect 40 632 42 634
rect 64 632 66 634
rect 70 632 72 634
rect 94 632 96 634
rect 100 632 102 634
rect 124 632 126 634
rect 130 632 132 634
rect 154 632 156 634
rect 160 632 162 634
rect 184 632 186 634
rect 414 632 416 634
rect 438 632 440 634
rect 444 632 446 634
rect 468 632 470 634
rect 474 632 476 634
rect 498 632 500 634
rect 504 632 506 634
rect 528 632 530 634
rect 534 632 536 634
rect 558 632 560 634
rect 564 632 566 634
rect 32 630 34 632
rect 62 630 64 632
rect 92 630 94 632
rect 122 630 124 632
rect 152 630 154 632
rect 182 630 184 632
rect 416 630 418 632
rect 446 630 448 632
rect 476 630 478 632
rect 506 630 508 632
rect 536 630 538 632
rect 566 630 568 632
rect 32 624 34 626
rect 62 624 64 626
rect 92 624 94 626
rect 122 624 124 626
rect 152 624 154 626
rect 182 624 184 626
rect 416 624 418 626
rect 446 624 448 626
rect 476 624 478 626
rect 506 624 508 626
rect 536 624 538 626
rect 566 624 568 626
rect 34 622 36 624
rect 40 622 42 624
rect 64 622 66 624
rect 70 622 72 624
rect 94 622 96 624
rect 100 622 102 624
rect 124 622 126 624
rect 130 622 132 624
rect 154 622 156 624
rect 160 622 162 624
rect 184 622 186 624
rect 414 622 416 624
rect 438 622 440 624
rect 444 622 446 624
rect 468 622 470 624
rect 474 622 476 624
rect 498 622 500 624
rect 504 622 506 624
rect 528 622 530 624
rect 534 622 536 624
rect 558 622 560 624
rect 564 622 566 624
rect 42 620 44 622
rect 72 620 74 622
rect 102 620 104 622
rect 132 620 134 622
rect 162 620 164 622
rect 436 620 438 622
rect 466 620 468 622
rect 496 620 498 622
rect 526 620 528 622
rect 556 620 558 622
rect 42 594 44 596
rect 72 594 74 596
rect 102 594 104 596
rect 132 594 134 596
rect 162 594 164 596
rect 436 594 438 596
rect 466 594 468 596
rect 496 594 498 596
rect 526 594 528 596
rect 556 594 558 596
rect 34 592 36 594
rect 40 592 42 594
rect 64 592 66 594
rect 70 592 72 594
rect 94 592 96 594
rect 100 592 102 594
rect 124 592 126 594
rect 130 592 132 594
rect 154 592 156 594
rect 160 592 162 594
rect 184 592 186 594
rect 414 592 416 594
rect 438 592 440 594
rect 444 592 446 594
rect 468 592 470 594
rect 474 592 476 594
rect 498 592 500 594
rect 504 592 506 594
rect 528 592 530 594
rect 534 592 536 594
rect 558 592 560 594
rect 564 592 566 594
rect 32 590 34 592
rect 62 590 64 592
rect 92 590 94 592
rect 122 590 124 592
rect 152 590 154 592
rect 182 590 184 592
rect 416 590 418 592
rect 446 590 448 592
rect 476 590 478 592
rect 506 590 508 592
rect 536 590 538 592
rect 566 590 568 592
rect 32 584 34 586
rect 62 584 64 586
rect 92 584 94 586
rect 506 584 508 586
rect 536 584 538 586
rect 566 584 568 586
rect 34 582 36 584
rect 40 582 42 584
rect 64 582 66 584
rect 70 582 72 584
rect 94 582 96 584
rect 100 582 102 584
rect 114 582 116 584
rect 130 582 132 584
rect 144 582 146 584
rect 160 582 162 584
rect 174 582 176 584
rect 424 582 426 584
rect 438 582 440 584
rect 454 582 456 584
rect 468 582 470 584
rect 484 582 486 584
rect 498 582 500 584
rect 504 582 506 584
rect 528 582 530 584
rect 534 582 536 584
rect 558 582 560 584
rect 564 582 566 584
rect 42 580 44 582
rect 72 580 74 582
rect 102 580 104 582
rect 112 580 114 582
rect 132 580 134 582
rect 142 580 144 582
rect 162 580 164 582
rect 172 580 174 582
rect 426 580 428 582
rect 436 580 438 582
rect 456 580 458 582
rect 466 580 468 582
rect 486 580 488 582
rect 496 580 498 582
rect 526 580 528 582
rect 556 580 558 582
rect 42 574 44 576
rect 72 574 74 576
rect 102 574 104 576
rect 112 574 114 576
rect 132 574 134 576
rect 142 574 144 576
rect 162 574 164 576
rect 172 574 174 576
rect 426 574 428 576
rect 436 574 438 576
rect 456 574 458 576
rect 466 574 468 576
rect 486 574 488 576
rect 496 574 498 576
rect 526 574 528 576
rect 556 574 558 576
rect 34 572 36 574
rect 40 572 42 574
rect 64 572 66 574
rect 70 572 72 574
rect 94 572 96 574
rect 100 572 102 574
rect 114 572 116 574
rect 130 572 132 574
rect 144 572 146 574
rect 160 572 162 574
rect 174 572 176 574
rect 424 572 426 574
rect 438 572 440 574
rect 454 572 456 574
rect 468 572 470 574
rect 484 572 486 574
rect 498 572 500 574
rect 504 572 506 574
rect 528 572 530 574
rect 534 572 536 574
rect 558 572 560 574
rect 564 572 566 574
rect 32 570 34 572
rect 62 570 64 572
rect 92 570 94 572
rect 506 570 508 572
rect 536 570 538 572
rect 566 570 568 572
rect 32 564 34 566
rect 62 564 64 566
rect 92 564 94 566
rect 122 564 124 566
rect 152 564 154 566
rect 182 564 184 566
rect 416 564 418 566
rect 446 564 448 566
rect 476 564 478 566
rect 506 564 508 566
rect 536 564 538 566
rect 566 564 568 566
rect 34 562 36 564
rect 40 562 42 564
rect 64 562 66 564
rect 70 562 72 564
rect 94 562 96 564
rect 100 562 102 564
rect 124 562 126 564
rect 130 562 132 564
rect 154 562 156 564
rect 160 562 162 564
rect 184 562 186 564
rect 414 562 416 564
rect 438 562 440 564
rect 444 562 446 564
rect 468 562 470 564
rect 474 562 476 564
rect 498 562 500 564
rect 504 562 506 564
rect 528 562 530 564
rect 534 562 536 564
rect 558 562 560 564
rect 564 562 566 564
rect 42 560 44 562
rect 72 560 74 562
rect 102 560 104 562
rect 132 560 134 562
rect 162 560 164 562
rect 436 560 438 562
rect 466 560 468 562
rect 496 560 498 562
rect 526 560 528 562
rect 556 560 558 562
rect 42 554 44 556
rect 72 554 74 556
rect 102 554 104 556
rect 132 554 134 556
rect 162 554 164 556
rect 436 554 438 556
rect 466 554 468 556
rect 496 554 498 556
rect 526 554 528 556
rect 556 554 558 556
rect 34 552 36 554
rect 40 552 42 554
rect 64 552 66 554
rect 70 552 72 554
rect 94 552 96 554
rect 100 552 102 554
rect 124 552 126 554
rect 130 552 132 554
rect 154 552 156 554
rect 160 552 162 554
rect 184 552 186 554
rect 414 552 416 554
rect 438 552 440 554
rect 444 552 446 554
rect 468 552 470 554
rect 474 552 476 554
rect 498 552 500 554
rect 504 552 506 554
rect 528 552 530 554
rect 534 552 536 554
rect 558 552 560 554
rect 564 552 566 554
rect 32 550 34 552
rect 62 550 64 552
rect 92 550 94 552
rect 122 550 124 552
rect 152 550 154 552
rect 182 550 184 552
rect 416 550 418 552
rect 446 550 448 552
rect 476 550 478 552
rect 506 550 508 552
rect 536 550 538 552
rect 566 550 568 552
rect 32 544 34 546
rect 62 544 64 546
rect 92 544 94 546
rect 122 544 124 546
rect 152 544 154 546
rect 182 544 184 546
rect 416 544 418 546
rect 446 544 448 546
rect 476 544 478 546
rect 506 544 508 546
rect 536 544 538 546
rect 566 544 568 546
rect 34 542 36 544
rect 40 542 42 544
rect 64 542 66 544
rect 70 542 72 544
rect 94 542 96 544
rect 100 542 102 544
rect 124 542 126 544
rect 130 542 132 544
rect 154 542 156 544
rect 160 542 162 544
rect 184 542 186 544
rect 414 542 416 544
rect 438 542 440 544
rect 444 542 446 544
rect 468 542 470 544
rect 474 542 476 544
rect 498 542 500 544
rect 504 542 506 544
rect 528 542 530 544
rect 534 542 536 544
rect 558 542 560 544
rect 564 542 566 544
rect 42 540 44 542
rect 72 540 74 542
rect 102 540 104 542
rect 132 540 134 542
rect 162 540 164 542
rect 436 540 438 542
rect 466 540 468 542
rect 496 540 498 542
rect 526 540 528 542
rect 556 540 558 542
rect 42 534 44 536
rect 72 534 74 536
rect 102 534 104 536
rect 132 534 134 536
rect 162 534 164 536
rect 436 534 438 536
rect 466 534 468 536
rect 496 534 498 536
rect 526 534 528 536
rect 556 534 558 536
rect 34 532 36 534
rect 40 532 42 534
rect 64 532 66 534
rect 70 532 72 534
rect 94 532 96 534
rect 100 532 102 534
rect 124 532 126 534
rect 130 532 132 534
rect 154 532 156 534
rect 160 532 162 534
rect 184 532 186 534
rect 414 532 416 534
rect 438 532 440 534
rect 444 532 446 534
rect 468 532 470 534
rect 474 532 476 534
rect 498 532 500 534
rect 504 532 506 534
rect 528 532 530 534
rect 534 532 536 534
rect 558 532 560 534
rect 564 532 566 534
rect 32 530 34 532
rect 62 530 64 532
rect 92 530 94 532
rect 122 530 124 532
rect 152 530 154 532
rect 182 530 184 532
rect 416 530 418 532
rect 446 530 448 532
rect 476 530 478 532
rect 506 530 508 532
rect 536 530 538 532
rect 566 530 568 532
rect 504 466 506 468
rect 502 464 504 466
rect 106 422 108 424
rect 492 422 494 424
rect 104 420 106 422
rect 494 420 496 422
rect 104 358 106 360
rect 494 358 496 360
rect 106 356 108 358
rect 492 356 494 358
rect 106 290 108 292
rect 492 290 494 292
rect 104 288 106 290
rect 494 288 496 290
rect 104 228 106 230
rect 494 228 496 230
rect 106 226 108 228
rect 492 226 494 228
rect 106 160 108 162
rect 492 160 494 162
rect 104 158 106 160
rect 494 158 496 160
rect 104 98 106 100
rect 494 98 496 100
rect 106 96 108 98
rect 492 96 494 98
rect 10 12 12 14
rect 588 12 590 14
rect 12 10 14 12
rect 586 10 588 12
<< error_s >>
rect 110 1598 118 1600
rect 134 1598 142 1600
rect 158 1598 166 1600
rect 182 1598 190 1600
rect 206 1598 214 1600
rect 230 1598 238 1600
rect 254 1598 262 1600
rect 278 1598 286 1600
rect 302 1598 310 1600
rect 326 1598 334 1600
rect 350 1598 358 1600
rect 374 1598 382 1600
rect 398 1598 406 1600
rect 422 1598 430 1600
rect 446 1598 454 1600
rect 470 1598 478 1600
rect 494 1598 502 1600
rect 98 1592 106 1594
rect 98 1588 100 1592
rect 104 1588 106 1592
rect 98 1586 106 1588
rect 122 1592 130 1594
rect 122 1588 124 1592
rect 128 1588 130 1592
rect 122 1586 130 1588
rect 146 1592 154 1594
rect 146 1588 148 1592
rect 152 1588 154 1592
rect 146 1586 154 1588
rect 170 1592 178 1594
rect 170 1588 172 1592
rect 176 1588 178 1592
rect 170 1586 178 1588
rect 194 1592 202 1594
rect 194 1588 196 1592
rect 200 1588 202 1592
rect 194 1586 202 1588
rect 218 1592 226 1594
rect 218 1588 220 1592
rect 224 1588 226 1592
rect 218 1586 226 1588
rect 242 1592 250 1594
rect 242 1588 244 1592
rect 248 1588 250 1592
rect 242 1586 250 1588
rect 266 1592 274 1594
rect 266 1588 268 1592
rect 272 1588 274 1592
rect 266 1586 274 1588
rect 290 1592 298 1594
rect 290 1588 292 1592
rect 296 1588 298 1592
rect 290 1586 298 1588
rect 314 1592 322 1594
rect 314 1588 316 1592
rect 320 1588 322 1592
rect 314 1586 322 1588
rect 338 1592 346 1594
rect 338 1588 340 1592
rect 344 1588 346 1592
rect 338 1586 346 1588
rect 362 1592 370 1594
rect 362 1588 364 1592
rect 368 1588 370 1592
rect 362 1586 370 1588
rect 386 1592 394 1594
rect 386 1588 388 1592
rect 392 1588 394 1592
rect 386 1586 394 1588
rect 410 1592 418 1594
rect 410 1588 412 1592
rect 416 1588 418 1592
rect 410 1586 418 1588
rect 434 1592 442 1594
rect 434 1588 436 1592
rect 440 1588 442 1592
rect 434 1586 442 1588
rect 458 1592 466 1594
rect 458 1588 460 1592
rect 464 1588 466 1592
rect 458 1586 466 1588
rect 482 1592 490 1594
rect 482 1588 484 1592
rect 488 1588 490 1592
rect 482 1586 490 1588
rect 110 1580 118 1582
rect 110 1576 112 1580
rect 116 1576 118 1580
rect 110 1574 118 1576
rect 134 1580 142 1582
rect 134 1576 136 1580
rect 140 1576 142 1580
rect 134 1574 142 1576
rect 158 1580 166 1582
rect 158 1576 160 1580
rect 164 1576 166 1580
rect 158 1574 166 1576
rect 182 1580 190 1582
rect 182 1576 184 1580
rect 188 1576 190 1580
rect 182 1574 190 1576
rect 206 1580 214 1582
rect 206 1576 208 1580
rect 212 1576 214 1580
rect 206 1574 214 1576
rect 230 1580 238 1582
rect 230 1576 232 1580
rect 236 1576 238 1580
rect 230 1574 238 1576
rect 254 1580 262 1582
rect 254 1576 256 1580
rect 260 1576 262 1580
rect 254 1574 262 1576
rect 278 1580 286 1582
rect 278 1576 280 1580
rect 284 1576 286 1580
rect 278 1574 286 1576
rect 302 1580 310 1582
rect 302 1576 304 1580
rect 308 1576 310 1580
rect 302 1574 310 1576
rect 326 1580 334 1582
rect 326 1576 328 1580
rect 332 1576 334 1580
rect 326 1574 334 1576
rect 350 1580 358 1582
rect 350 1576 352 1580
rect 356 1576 358 1580
rect 350 1574 358 1576
rect 374 1580 382 1582
rect 374 1576 376 1580
rect 380 1576 382 1580
rect 374 1574 382 1576
rect 398 1580 406 1582
rect 398 1576 400 1580
rect 404 1576 406 1580
rect 398 1574 406 1576
rect 422 1580 430 1582
rect 422 1576 424 1580
rect 428 1576 430 1580
rect 422 1574 430 1576
rect 446 1580 454 1582
rect 446 1576 448 1580
rect 452 1576 454 1580
rect 446 1574 454 1576
rect 470 1580 478 1582
rect 470 1576 472 1580
rect 476 1576 478 1580
rect 470 1574 478 1576
rect 494 1580 502 1582
rect 494 1576 496 1580
rect 500 1576 502 1580
rect 494 1574 502 1576
rect 98 1568 106 1570
rect 98 1564 100 1568
rect 104 1564 106 1568
rect 98 1562 106 1564
rect 122 1568 130 1570
rect 122 1564 124 1568
rect 128 1564 130 1568
rect 122 1562 130 1564
rect 146 1568 154 1570
rect 146 1564 148 1568
rect 152 1564 154 1568
rect 146 1562 154 1564
rect 170 1568 178 1570
rect 170 1564 172 1568
rect 176 1564 178 1568
rect 170 1562 178 1564
rect 194 1568 202 1570
rect 194 1564 196 1568
rect 200 1564 202 1568
rect 194 1562 202 1564
rect 218 1568 226 1570
rect 218 1564 220 1568
rect 224 1564 226 1568
rect 218 1562 226 1564
rect 242 1568 250 1570
rect 242 1564 244 1568
rect 248 1564 250 1568
rect 242 1562 250 1564
rect 266 1568 274 1570
rect 266 1564 268 1568
rect 272 1564 274 1568
rect 266 1562 274 1564
rect 290 1568 298 1570
rect 290 1564 292 1568
rect 296 1564 298 1568
rect 290 1562 298 1564
rect 314 1568 322 1570
rect 314 1564 316 1568
rect 320 1564 322 1568
rect 314 1562 322 1564
rect 338 1568 346 1570
rect 338 1564 340 1568
rect 344 1564 346 1568
rect 338 1562 346 1564
rect 362 1568 370 1570
rect 362 1564 364 1568
rect 368 1564 370 1568
rect 362 1562 370 1564
rect 386 1568 394 1570
rect 386 1564 388 1568
rect 392 1564 394 1568
rect 386 1562 394 1564
rect 410 1568 418 1570
rect 410 1564 412 1568
rect 416 1564 418 1568
rect 410 1562 418 1564
rect 434 1568 442 1570
rect 434 1564 436 1568
rect 440 1564 442 1568
rect 434 1562 442 1564
rect 458 1568 466 1570
rect 458 1564 460 1568
rect 464 1564 466 1568
rect 458 1562 466 1564
rect 482 1568 490 1570
rect 482 1564 484 1568
rect 488 1564 490 1568
rect 482 1562 490 1564
rect 110 1556 118 1558
rect 110 1552 112 1556
rect 116 1552 118 1556
rect 110 1550 118 1552
rect 134 1556 142 1558
rect 134 1552 136 1556
rect 140 1552 142 1556
rect 134 1550 142 1552
rect 158 1556 166 1558
rect 158 1552 160 1556
rect 164 1552 166 1556
rect 158 1550 166 1552
rect 182 1556 190 1558
rect 182 1552 184 1556
rect 188 1552 190 1556
rect 182 1550 190 1552
rect 206 1556 214 1558
rect 206 1552 208 1556
rect 212 1552 214 1556
rect 206 1550 214 1552
rect 230 1556 238 1558
rect 230 1552 232 1556
rect 236 1552 238 1556
rect 230 1550 238 1552
rect 254 1556 262 1558
rect 254 1552 256 1556
rect 260 1552 262 1556
rect 254 1550 262 1552
rect 278 1556 286 1558
rect 278 1552 280 1556
rect 284 1552 286 1556
rect 278 1550 286 1552
rect 302 1556 310 1558
rect 302 1552 304 1556
rect 308 1552 310 1556
rect 302 1550 310 1552
rect 326 1556 334 1558
rect 326 1552 328 1556
rect 332 1552 334 1556
rect 326 1550 334 1552
rect 350 1556 358 1558
rect 350 1552 352 1556
rect 356 1552 358 1556
rect 350 1550 358 1552
rect 374 1556 382 1558
rect 374 1552 376 1556
rect 380 1552 382 1556
rect 374 1550 382 1552
rect 398 1556 406 1558
rect 398 1552 400 1556
rect 404 1552 406 1556
rect 398 1550 406 1552
rect 422 1556 430 1558
rect 422 1552 424 1556
rect 428 1552 430 1556
rect 422 1550 430 1552
rect 446 1556 454 1558
rect 446 1552 448 1556
rect 452 1552 454 1556
rect 446 1550 454 1552
rect 470 1556 478 1558
rect 470 1552 472 1556
rect 476 1552 478 1556
rect 470 1550 478 1552
rect 494 1556 502 1558
rect 494 1552 496 1556
rect 500 1552 502 1556
rect 494 1550 502 1552
rect 98 1544 106 1546
rect 98 1540 100 1544
rect 104 1540 106 1544
rect 98 1538 106 1540
rect 122 1544 130 1546
rect 122 1540 124 1544
rect 128 1540 130 1544
rect 122 1538 130 1540
rect 146 1544 154 1546
rect 146 1540 148 1544
rect 152 1540 154 1544
rect 146 1538 154 1540
rect 170 1544 178 1546
rect 170 1540 172 1544
rect 176 1540 178 1544
rect 170 1538 178 1540
rect 194 1544 202 1546
rect 194 1540 196 1544
rect 200 1540 202 1544
rect 194 1538 202 1540
rect 218 1544 226 1546
rect 218 1540 220 1544
rect 224 1540 226 1544
rect 218 1538 226 1540
rect 242 1544 250 1546
rect 242 1540 244 1544
rect 248 1540 250 1544
rect 242 1538 250 1540
rect 266 1544 274 1546
rect 266 1540 268 1544
rect 272 1540 274 1544
rect 266 1538 274 1540
rect 290 1544 298 1546
rect 290 1540 292 1544
rect 296 1540 298 1544
rect 290 1538 298 1540
rect 314 1544 322 1546
rect 314 1540 316 1544
rect 320 1540 322 1544
rect 314 1538 322 1540
rect 338 1544 346 1546
rect 338 1540 340 1544
rect 344 1540 346 1544
rect 338 1538 346 1540
rect 362 1544 370 1546
rect 362 1540 364 1544
rect 368 1540 370 1544
rect 362 1538 370 1540
rect 386 1544 394 1546
rect 386 1540 388 1544
rect 392 1540 394 1544
rect 386 1538 394 1540
rect 410 1544 418 1546
rect 410 1540 412 1544
rect 416 1540 418 1544
rect 410 1538 418 1540
rect 434 1544 442 1546
rect 434 1540 436 1544
rect 440 1540 442 1544
rect 434 1538 442 1540
rect 458 1544 466 1546
rect 458 1540 460 1544
rect 464 1540 466 1544
rect 458 1538 466 1540
rect 482 1544 490 1546
rect 482 1540 484 1544
rect 488 1540 490 1544
rect 482 1538 490 1540
<< nwell >>
rect 34 858 566 1306
rect -6 498 606 660
rect -6 22 22 498
rect 578 22 606 498
rect -6 -6 606 22
<< ntransistor >>
rect 76 432 276 438
rect 324 432 524 438
rect 76 342 276 348
rect 76 300 276 306
rect 324 342 524 348
rect 324 300 524 306
rect 76 212 276 218
rect 76 170 276 176
rect 324 212 524 218
rect 324 170 524 176
rect 76 82 276 88
rect 324 82 524 88
<< ptransistor >>
rect 76 1252 276 1258
rect 324 1252 524 1258
rect 76 1164 276 1170
rect 76 1124 276 1130
rect 324 1164 524 1170
rect 324 1124 524 1130
rect 76 1036 276 1042
rect 76 994 276 1000
rect 76 906 276 912
rect 324 1036 524 1042
rect 324 994 524 1000
rect 324 906 524 912
<< ndiffusion >>
rect 76 454 276 456
rect 76 446 82 454
rect 190 446 276 454
rect 76 438 276 446
rect 76 400 276 432
rect 76 392 112 400
rect 240 392 276 400
rect 76 388 276 392
rect 76 380 112 388
rect 240 380 276 388
rect 76 348 276 380
rect 324 454 524 456
rect 324 446 410 454
rect 518 446 524 454
rect 324 438 524 446
rect 76 334 276 342
rect 76 326 82 334
rect 240 326 276 334
rect 76 322 276 326
rect 76 314 82 322
rect 240 314 276 322
rect 76 306 276 314
rect 76 268 276 300
rect 76 250 112 268
rect 240 250 276 268
rect 76 218 276 250
rect 324 400 524 432
rect 324 392 360 400
rect 488 392 524 400
rect 324 388 524 392
rect 324 380 360 388
rect 488 380 524 388
rect 324 348 524 380
rect 324 334 524 342
rect 324 326 360 334
rect 518 326 524 334
rect 324 322 524 326
rect 324 314 360 322
rect 518 314 524 322
rect 324 306 524 314
rect 76 204 276 212
rect 76 196 82 204
rect 240 196 276 204
rect 76 192 276 196
rect 76 184 82 192
rect 240 184 276 192
rect 76 176 276 184
rect 76 138 276 170
rect 76 120 112 138
rect 240 120 276 138
rect 76 88 276 120
rect 324 268 524 300
rect 324 250 360 268
rect 488 250 524 268
rect 324 218 524 250
rect 324 204 524 212
rect 324 196 360 204
rect 518 196 524 204
rect 324 192 524 196
rect 324 184 360 192
rect 518 184 524 192
rect 324 176 524 184
rect 324 138 524 170
rect 324 120 360 138
rect 488 120 524 138
rect 324 88 524 120
rect 76 74 276 82
rect 76 66 82 74
rect 190 66 276 74
rect 76 64 276 66
rect 324 74 524 82
rect 324 66 410 74
rect 518 66 524 74
rect 324 64 524 66
<< pdiffusion >>
rect 76 1274 276 1276
rect 76 1266 82 1274
rect 240 1266 276 1274
rect 76 1258 276 1266
rect 76 1220 276 1252
rect 76 1202 112 1220
rect 240 1202 276 1220
rect 76 1170 276 1202
rect 324 1274 524 1276
rect 324 1266 360 1274
rect 518 1266 524 1274
rect 324 1258 524 1266
rect 76 1156 276 1164
rect 76 1138 82 1156
rect 240 1138 276 1156
rect 76 1130 276 1138
rect 76 1092 276 1124
rect 76 1074 112 1092
rect 240 1074 276 1092
rect 76 1042 276 1074
rect 324 1220 524 1252
rect 324 1202 360 1220
rect 488 1202 524 1220
rect 324 1170 524 1202
rect 324 1156 524 1164
rect 324 1138 360 1156
rect 518 1138 524 1156
rect 324 1130 524 1138
rect 76 1028 276 1036
rect 76 1020 82 1028
rect 240 1020 276 1028
rect 76 1016 276 1020
rect 76 1008 82 1016
rect 240 1008 276 1016
rect 76 1000 276 1008
rect 76 962 276 994
rect 76 944 112 962
rect 240 944 276 962
rect 76 912 276 944
rect 76 898 276 906
rect 76 890 82 898
rect 190 890 276 898
rect 76 888 276 890
rect 324 1092 524 1124
rect 324 1074 360 1092
rect 488 1074 524 1092
rect 324 1042 524 1074
rect 324 1028 524 1036
rect 324 1020 360 1028
rect 518 1020 524 1028
rect 324 1016 524 1020
rect 324 1008 360 1016
rect 518 1008 524 1016
rect 324 1000 524 1008
rect 324 962 524 994
rect 324 944 360 962
rect 488 944 524 962
rect 324 912 524 944
rect 324 898 524 906
rect 324 890 410 898
rect 518 890 524 898
rect 324 888 524 890
<< ndcontact >>
rect 82 446 190 454
rect 112 392 240 400
rect 112 380 240 388
rect 410 446 518 454
rect 82 326 240 334
rect 82 314 240 322
rect 112 250 240 268
rect 360 392 488 400
rect 360 380 488 388
rect 360 326 518 334
rect 360 314 518 322
rect 82 196 240 204
rect 82 184 240 192
rect 112 120 240 138
rect 360 250 488 268
rect 360 196 518 204
rect 360 184 518 192
rect 360 120 488 138
rect 82 66 190 74
rect 410 66 518 74
<< pdcontact >>
rect 82 1266 240 1274
rect 112 1202 240 1220
rect 360 1266 518 1274
rect 82 1138 240 1156
rect 112 1074 240 1092
rect 360 1202 488 1220
rect 360 1138 518 1156
rect 82 1020 240 1028
rect 82 1008 240 1016
rect 112 944 240 962
rect 82 890 190 898
rect 360 1074 488 1092
rect 360 1020 518 1028
rect 360 1008 518 1016
rect 360 944 488 962
rect 410 890 518 898
<< psubstratepdiff >>
rect 0 1338 600 1340
rect 0 840 2 1338
rect 190 1320 410 1338
rect 20 1318 580 1320
rect 20 846 22 1318
rect 578 846 580 1318
rect 20 844 580 846
rect 20 840 44 844
rect 0 836 44 840
rect 52 836 74 844
rect 82 836 104 844
rect 112 836 134 844
rect 142 836 164 844
rect 172 836 428 844
rect 436 836 458 844
rect 466 836 488 844
rect 496 836 518 844
rect 526 836 548 844
rect 556 840 580 844
rect 598 840 600 1338
rect 556 836 600 840
rect 0 828 4 836
rect 12 828 24 836
rect 42 828 54 836
rect 72 828 84 836
rect 102 828 114 836
rect 132 828 144 836
rect 162 828 174 836
rect 192 834 408 836
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 184 828
rect 0 818 14 826
rect 22 818 34 826
rect 52 818 64 826
rect 82 818 94 826
rect 112 818 124 826
rect 142 818 154 826
rect 172 818 184 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 184 818
rect 192 826 286 834
rect 314 826 408 834
rect 426 828 438 836
rect 456 828 468 836
rect 486 828 498 836
rect 516 828 528 836
rect 546 828 558 836
rect 576 828 588 836
rect 596 828 600 836
rect 0 808 4 816
rect 12 808 24 816
rect 42 808 54 816
rect 72 808 84 816
rect 102 808 114 816
rect 132 808 144 816
rect 162 808 174 816
rect 192 814 408 826
rect 416 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 416 818 428 826
rect 446 818 458 826
rect 476 818 488 826
rect 506 818 518 826
rect 536 818 548 826
rect 566 818 578 826
rect 586 818 600 826
rect 416 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 184 808
rect 0 798 14 806
rect 22 798 34 806
rect 52 798 64 806
rect 82 798 94 806
rect 112 798 124 806
rect 142 798 154 806
rect 172 798 184 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 184 798
rect 192 806 286 814
rect 314 806 408 814
rect 426 808 438 816
rect 456 808 468 816
rect 486 808 498 816
rect 516 808 528 816
rect 546 808 558 816
rect 576 808 588 816
rect 596 808 600 816
rect 0 788 4 796
rect 12 788 24 796
rect 42 788 54 796
rect 72 788 84 796
rect 102 788 114 796
rect 132 788 144 796
rect 162 788 174 796
rect 192 794 408 806
rect 416 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 416 798 428 806
rect 446 798 458 806
rect 476 798 488 806
rect 506 798 518 806
rect 536 798 548 806
rect 566 798 578 806
rect 586 798 600 806
rect 416 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 184 788
rect 0 778 14 786
rect 22 778 34 786
rect 52 778 64 786
rect 82 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 776 124 786
rect 142 776 154 786
rect 172 776 184 786
rect 192 786 286 794
rect 314 786 408 794
rect 426 788 438 796
rect 456 788 468 796
rect 486 788 498 796
rect 516 788 528 796
rect 546 788 558 796
rect 576 788 588 796
rect 596 788 600 796
rect 192 776 408 786
rect 416 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 416 776 428 786
rect 446 776 458 786
rect 476 776 488 786
rect 506 778 518 786
rect 536 778 548 786
rect 566 778 578 786
rect 586 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 0 768 4 776
rect 12 768 24 776
rect 42 768 54 776
rect 72 768 84 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 14 766
rect 22 758 34 766
rect 52 758 64 766
rect 82 758 94 766
rect 112 758 124 768
rect 142 758 154 768
rect 172 758 184 768
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 184 758
rect 192 758 286 776
rect 314 758 408 776
rect 516 768 528 776
rect 546 768 558 776
rect 576 768 588 776
rect 596 768 600 776
rect 0 748 4 756
rect 12 748 24 756
rect 42 748 54 756
rect 72 748 84 756
rect 102 748 114 756
rect 132 748 144 756
rect 162 748 174 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 184 748
rect 0 738 14 746
rect 22 738 34 746
rect 52 738 64 746
rect 82 738 94 746
rect 112 738 124 746
rect 142 738 154 746
rect 172 738 184 746
rect 192 746 408 758
rect 416 758 428 768
rect 446 758 458 768
rect 476 758 488 768
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 518 766
rect 536 758 548 766
rect 566 758 578 766
rect 586 758 600 766
rect 416 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 426 748 438 756
rect 456 748 468 756
rect 486 748 498 756
rect 516 748 528 756
rect 546 748 558 756
rect 576 748 588 756
rect 596 748 600 756
rect 192 738 286 746
rect 314 738 408 746
rect 416 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 416 738 428 746
rect 446 738 458 746
rect 476 738 488 746
rect 506 738 518 746
rect 536 738 548 746
rect 566 738 578 746
rect 586 738 600 746
rect 0 736 600 738
rect 0 728 4 736
rect 12 728 24 736
rect 32 728 568 736
rect 576 728 588 736
rect 596 728 600 736
rect 0 726 600 728
rect 0 718 14 726
rect 22 718 34 726
rect 52 718 64 726
rect 82 718 94 726
rect 112 718 124 726
rect 142 718 154 726
rect 172 718 184 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 184 718
rect 192 718 286 726
rect 314 718 408 726
rect 0 708 4 716
rect 12 708 24 716
rect 42 708 54 716
rect 72 708 84 716
rect 102 708 114 716
rect 132 708 144 716
rect 162 708 174 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 184 708
rect 0 698 14 706
rect 22 698 34 706
rect 52 698 64 706
rect 82 698 94 706
rect 112 698 124 706
rect 142 698 154 706
rect 172 698 184 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 184 698
rect 192 706 408 718
rect 416 718 428 726
rect 446 718 458 726
rect 476 718 488 726
rect 506 718 518 726
rect 536 718 548 726
rect 566 718 578 726
rect 586 718 600 726
rect 416 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 426 708 438 716
rect 456 708 468 716
rect 486 708 498 716
rect 516 708 528 716
rect 546 708 558 716
rect 576 708 588 716
rect 596 708 600 716
rect 192 698 286 706
rect 314 698 408 706
rect 0 688 4 696
rect 12 688 24 696
rect 42 688 54 696
rect 72 688 84 696
rect 102 688 114 696
rect 132 688 144 696
rect 162 688 174 696
rect 192 688 408 698
rect 416 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 416 698 428 706
rect 446 698 458 706
rect 476 698 488 706
rect 506 698 518 706
rect 536 698 548 706
rect 566 698 578 706
rect 586 698 600 706
rect 416 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 426 688 438 696
rect 456 688 468 696
rect 486 688 498 696
rect 516 688 528 696
rect 546 688 558 696
rect 576 688 588 696
rect 596 688 600 696
rect 0 686 600 688
rect 28 486 572 492
rect 28 484 286 486
rect 28 466 36 484
rect 74 466 82 484
rect 28 462 82 466
rect 28 454 36 462
rect 54 460 82 462
rect 54 454 60 460
rect 28 442 60 454
rect 28 434 36 442
rect 54 434 60 442
rect 76 456 82 460
rect 190 460 286 484
rect 190 456 276 460
rect 284 458 286 460
rect 314 474 572 486
rect 314 460 416 474
rect 564 466 572 474
rect 314 458 316 460
rect 28 422 60 434
rect 28 414 36 422
rect 54 414 60 422
rect 28 402 60 414
rect 28 394 36 402
rect 54 394 60 402
rect 28 382 60 394
rect 28 374 36 382
rect 54 374 60 382
rect 28 362 60 374
rect 28 354 36 362
rect 54 354 60 362
rect 28 342 60 354
rect 28 334 36 342
rect 54 334 60 342
rect 28 322 60 334
rect 28 314 36 322
rect 54 314 60 322
rect 28 302 60 314
rect 28 294 36 302
rect 54 294 60 302
rect 28 282 60 294
rect 28 274 36 282
rect 54 274 60 282
rect 28 262 60 274
rect 28 254 36 262
rect 54 254 60 262
rect 28 242 60 254
rect 28 234 36 242
rect 54 234 60 242
rect 28 222 60 234
rect 28 214 36 222
rect 54 214 60 222
rect 28 202 60 214
rect 28 194 36 202
rect 54 194 60 202
rect 28 182 60 194
rect 28 174 36 182
rect 54 174 60 182
rect 28 162 60 174
rect 28 154 36 162
rect 54 154 60 162
rect 28 142 60 154
rect 28 134 36 142
rect 54 134 60 142
rect 28 122 60 134
rect 28 114 36 122
rect 54 114 60 122
rect 28 102 60 114
rect 28 94 36 102
rect 54 94 60 102
rect 28 82 60 94
rect 284 400 316 458
rect 324 456 416 460
rect 504 462 572 466
rect 504 460 546 462
rect 504 456 524 460
rect 540 454 546 460
rect 564 454 572 462
rect 540 442 572 454
rect 284 392 291 400
rect 309 392 316 400
rect 284 384 316 392
rect 284 376 291 384
rect 309 376 316 384
rect 284 272 316 376
rect 284 264 291 272
rect 309 264 316 272
rect 284 256 316 264
rect 284 248 291 256
rect 309 248 316 256
rect 284 144 316 248
rect 284 136 291 144
rect 309 136 316 144
rect 284 128 316 136
rect 284 120 291 128
rect 309 120 316 128
rect 284 112 316 120
rect 284 104 291 112
rect 309 104 316 112
rect 284 96 316 104
rect 284 88 291 96
rect 309 88 316 96
rect 28 74 36 82
rect 54 74 60 82
rect 28 62 60 74
rect 28 54 36 62
rect 54 60 60 62
rect 76 62 276 64
rect 76 60 88 62
rect 54 54 88 60
rect 28 42 88 54
rect 28 34 36 42
rect 84 34 88 42
rect 96 34 108 62
rect 116 34 128 62
rect 136 34 148 62
rect 156 34 168 62
rect 176 34 188 62
rect 196 60 276 62
rect 284 60 316 88
rect 540 434 546 442
rect 564 434 572 442
rect 540 422 572 434
rect 540 414 546 422
rect 564 414 572 422
rect 540 402 572 414
rect 540 394 546 402
rect 564 394 572 402
rect 540 382 572 394
rect 540 374 546 382
rect 564 374 572 382
rect 540 362 572 374
rect 540 354 546 362
rect 564 354 572 362
rect 540 342 572 354
rect 540 334 546 342
rect 564 334 572 342
rect 540 322 572 334
rect 540 314 546 322
rect 564 314 572 322
rect 540 302 572 314
rect 540 294 546 302
rect 564 294 572 302
rect 540 282 572 294
rect 540 274 546 282
rect 564 274 572 282
rect 540 262 572 274
rect 540 254 546 262
rect 564 254 572 262
rect 540 242 572 254
rect 540 234 546 242
rect 564 234 572 242
rect 540 222 572 234
rect 540 214 546 222
rect 564 214 572 222
rect 540 202 572 214
rect 540 194 546 202
rect 564 194 572 202
rect 540 182 572 194
rect 540 174 546 182
rect 564 174 572 182
rect 540 162 572 174
rect 540 154 546 162
rect 564 154 572 162
rect 540 142 572 154
rect 540 134 546 142
rect 564 134 572 142
rect 540 122 572 134
rect 540 114 546 122
rect 564 114 572 122
rect 540 102 572 114
rect 540 94 546 102
rect 564 94 572 102
rect 540 82 572 94
rect 324 62 524 64
rect 324 60 404 62
rect 196 34 404 60
rect 412 34 424 62
rect 432 34 444 62
rect 452 34 464 62
rect 472 34 484 62
rect 492 34 504 62
rect 512 60 524 62
rect 540 74 546 82
rect 564 74 572 82
rect 540 62 572 74
rect 540 60 546 62
rect 512 54 546 60
rect 564 54 572 62
rect 512 42 572 54
rect 512 34 516 42
rect 564 34 572 42
rect 28 28 572 34
<< nsubstratendiff >>
rect 40 1298 560 1300
rect 40 1290 51 1298
rect 59 1290 72 1298
rect 80 1294 520 1298
rect 40 1289 82 1290
rect 40 1288 62 1289
rect 40 1280 41 1288
rect 49 1281 62 1288
rect 70 1286 82 1289
rect 90 1286 102 1294
rect 110 1286 122 1294
rect 130 1286 142 1294
rect 150 1286 162 1294
rect 170 1286 182 1294
rect 190 1286 202 1294
rect 210 1286 222 1294
rect 230 1286 370 1294
rect 378 1286 390 1294
rect 398 1286 410 1294
rect 418 1286 430 1294
rect 438 1286 450 1294
rect 458 1286 470 1294
rect 478 1286 490 1294
rect 498 1286 510 1294
rect 528 1290 541 1298
rect 549 1290 560 1298
rect 518 1289 560 1290
rect 518 1286 530 1289
rect 70 1284 530 1286
rect 70 1281 92 1284
rect 49 1280 92 1281
rect 40 1278 60 1280
rect 40 1270 51 1278
rect 59 1270 60 1278
rect 40 1268 60 1270
rect 40 1260 41 1268
rect 49 1260 60 1268
rect 40 1258 60 1260
rect 76 1276 92 1280
rect 100 1276 112 1284
rect 120 1276 132 1284
rect 140 1276 152 1284
rect 160 1276 172 1284
rect 180 1276 192 1284
rect 200 1276 212 1284
rect 220 1276 232 1284
rect 240 1280 360 1284
rect 240 1276 276 1280
rect 40 1250 51 1258
rect 59 1250 60 1258
rect 40 1248 60 1250
rect 40 1240 41 1248
rect 49 1240 60 1248
rect 40 1238 60 1240
rect 40 1230 51 1238
rect 59 1230 60 1238
rect 40 1228 60 1230
rect 40 1220 41 1228
rect 49 1220 60 1228
rect 40 1218 60 1220
rect 40 1210 51 1218
rect 59 1210 60 1218
rect 40 1208 60 1210
rect 40 1200 41 1208
rect 49 1200 60 1208
rect 40 1198 60 1200
rect 40 1190 51 1198
rect 59 1190 60 1198
rect 40 1188 60 1190
rect 40 1180 41 1188
rect 49 1180 60 1188
rect 40 1178 60 1180
rect 40 1170 51 1178
rect 59 1170 60 1178
rect 40 1168 60 1170
rect 40 1160 41 1168
rect 49 1160 60 1168
rect 40 1158 60 1160
rect 40 1150 51 1158
rect 59 1150 60 1158
rect 40 1148 60 1150
rect 40 1140 41 1148
rect 49 1140 60 1148
rect 40 1138 60 1140
rect 40 1130 51 1138
rect 59 1130 60 1138
rect 40 1128 60 1130
rect 40 1120 41 1128
rect 49 1120 60 1128
rect 40 1118 60 1120
rect 40 1110 51 1118
rect 59 1110 60 1118
rect 40 1108 60 1110
rect 40 1100 41 1108
rect 49 1100 60 1108
rect 40 1098 60 1100
rect 40 1090 51 1098
rect 59 1090 60 1098
rect 40 1088 60 1090
rect 40 1080 41 1088
rect 49 1080 60 1088
rect 40 1078 60 1080
rect 40 1070 51 1078
rect 59 1070 60 1078
rect 40 1068 60 1070
rect 40 1060 41 1068
rect 49 1060 60 1068
rect 40 1058 60 1060
rect 40 1050 51 1058
rect 59 1050 60 1058
rect 40 1048 60 1050
rect 40 1040 41 1048
rect 49 1040 60 1048
rect 40 1038 60 1040
rect 40 1030 51 1038
rect 59 1030 60 1038
rect 40 1028 60 1030
rect 40 1020 41 1028
rect 49 1020 60 1028
rect 40 1018 60 1020
rect 40 1010 51 1018
rect 59 1010 60 1018
rect 40 1008 60 1010
rect 40 1000 41 1008
rect 49 1000 60 1008
rect 40 998 60 1000
rect 40 990 51 998
rect 59 990 60 998
rect 40 988 60 990
rect 40 980 41 988
rect 49 980 60 988
rect 40 978 60 980
rect 40 970 51 978
rect 59 970 60 978
rect 40 968 60 970
rect 40 960 41 968
rect 49 960 60 968
rect 40 958 60 960
rect 40 950 51 958
rect 59 950 60 958
rect 40 948 60 950
rect 40 940 41 948
rect 49 940 60 948
rect 40 938 60 940
rect 40 930 51 938
rect 59 930 60 938
rect 40 928 60 930
rect 40 920 41 928
rect 49 920 60 928
rect 40 918 60 920
rect 40 910 51 918
rect 59 910 60 918
rect 40 908 60 910
rect 40 900 41 908
rect 49 900 60 908
rect 284 1226 316 1280
rect 324 1276 360 1280
rect 368 1276 380 1284
rect 388 1276 400 1284
rect 408 1276 420 1284
rect 428 1276 440 1284
rect 448 1276 460 1284
rect 468 1276 480 1284
rect 488 1276 500 1284
rect 508 1281 530 1284
rect 538 1288 560 1289
rect 538 1281 551 1288
rect 508 1280 551 1281
rect 559 1280 560 1288
rect 508 1276 524 1280
rect 540 1278 560 1280
rect 540 1270 541 1278
rect 549 1270 560 1278
rect 540 1268 560 1270
rect 540 1260 551 1268
rect 559 1260 560 1268
rect 540 1258 560 1260
rect 284 1218 291 1226
rect 309 1218 316 1226
rect 284 1210 316 1218
rect 284 1202 291 1210
rect 309 1202 316 1210
rect 284 1098 316 1202
rect 284 1090 291 1098
rect 309 1090 316 1098
rect 284 1082 316 1090
rect 284 1074 291 1082
rect 309 1074 316 1082
rect 40 898 60 900
rect 40 890 51 898
rect 59 890 60 898
rect 40 888 60 890
rect 40 880 41 888
rect 49 884 60 888
rect 76 884 276 888
rect 284 884 316 1074
rect 540 1250 541 1258
rect 549 1250 560 1258
rect 540 1248 560 1250
rect 540 1240 551 1248
rect 559 1240 560 1248
rect 540 1238 560 1240
rect 540 1230 541 1238
rect 549 1230 560 1238
rect 540 1228 560 1230
rect 540 1220 551 1228
rect 559 1220 560 1228
rect 540 1218 560 1220
rect 540 1210 541 1218
rect 549 1210 560 1218
rect 540 1208 560 1210
rect 540 1200 551 1208
rect 559 1200 560 1208
rect 540 1198 560 1200
rect 540 1190 541 1198
rect 549 1190 560 1198
rect 540 1188 560 1190
rect 540 1180 551 1188
rect 559 1180 560 1188
rect 540 1178 560 1180
rect 540 1170 541 1178
rect 549 1170 560 1178
rect 540 1168 560 1170
rect 540 1160 551 1168
rect 559 1160 560 1168
rect 540 1158 560 1160
rect 540 1150 541 1158
rect 549 1150 560 1158
rect 540 1148 560 1150
rect 540 1140 551 1148
rect 559 1140 560 1148
rect 540 1138 560 1140
rect 540 1130 541 1138
rect 549 1130 560 1138
rect 540 1128 560 1130
rect 540 1120 551 1128
rect 559 1120 560 1128
rect 540 1118 560 1120
rect 540 1110 541 1118
rect 549 1110 560 1118
rect 540 1108 560 1110
rect 540 1100 551 1108
rect 559 1100 560 1108
rect 540 1098 560 1100
rect 540 1090 541 1098
rect 549 1090 560 1098
rect 540 1088 560 1090
rect 540 1080 551 1088
rect 559 1080 560 1088
rect 540 1078 560 1080
rect 540 1070 541 1078
rect 549 1070 560 1078
rect 540 1068 560 1070
rect 540 1060 551 1068
rect 559 1060 560 1068
rect 540 1058 560 1060
rect 540 1050 541 1058
rect 549 1050 560 1058
rect 540 1048 560 1050
rect 540 1040 551 1048
rect 559 1040 560 1048
rect 540 1038 560 1040
rect 540 1030 541 1038
rect 549 1030 560 1038
rect 540 1028 560 1030
rect 540 1020 551 1028
rect 559 1020 560 1028
rect 540 1018 560 1020
rect 540 1010 541 1018
rect 549 1010 560 1018
rect 540 1008 560 1010
rect 540 1000 551 1008
rect 559 1000 560 1008
rect 540 998 560 1000
rect 540 990 541 998
rect 549 990 560 998
rect 540 988 560 990
rect 540 980 551 988
rect 559 980 560 988
rect 540 978 560 980
rect 540 970 541 978
rect 549 970 560 978
rect 540 968 560 970
rect 540 960 551 968
rect 559 960 560 968
rect 540 958 560 960
rect 540 950 541 958
rect 549 950 560 958
rect 540 948 560 950
rect 540 940 551 948
rect 559 940 560 948
rect 540 938 560 940
rect 540 930 541 938
rect 549 930 560 938
rect 540 928 560 930
rect 540 920 551 928
rect 559 920 560 928
rect 540 918 560 920
rect 540 910 541 918
rect 549 910 560 918
rect 540 908 560 910
rect 324 884 524 888
rect 540 900 551 908
rect 559 900 560 908
rect 540 898 560 900
rect 540 890 541 898
rect 549 890 560 898
rect 540 888 560 890
rect 540 884 551 888
rect 49 883 551 884
rect 49 880 62 883
rect 40 873 62 880
rect 40 865 42 873
rect 190 865 286 883
rect 314 865 410 883
rect 538 880 551 883
rect 559 880 560 888
rect 538 873 560 880
rect 558 865 560 873
rect 40 864 560 865
rect 0 652 600 654
rect 0 644 4 652
rect 12 644 24 652
rect 42 644 54 652
rect 72 644 84 652
rect 102 644 114 652
rect 132 644 144 652
rect 162 644 174 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 0 634 14 642
rect 22 634 34 642
rect 52 634 64 642
rect 82 634 94 642
rect 112 634 124 642
rect 142 634 154 642
rect 172 634 184 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 192 642 408 652
rect 426 644 438 652
rect 456 644 468 652
rect 486 644 498 652
rect 516 644 528 652
rect 546 644 558 652
rect 576 644 588 652
rect 596 644 600 652
rect 192 634 286 642
rect 314 634 408 642
rect 0 624 4 632
rect 12 624 24 632
rect 42 624 54 632
rect 72 624 84 632
rect 102 624 114 632
rect 132 624 144 632
rect 162 624 174 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 0 614 14 622
rect 22 614 34 622
rect 52 614 64 622
rect 82 614 94 622
rect 112 614 124 622
rect 142 614 154 622
rect 172 614 184 622
rect 192 622 408 634
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 416 634 428 642
rect 446 634 458 642
rect 476 634 488 642
rect 506 634 518 642
rect 536 634 548 642
rect 566 634 578 642
rect 586 634 600 642
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 426 624 438 632
rect 456 624 468 632
rect 486 624 498 632
rect 516 624 528 632
rect 546 624 558 632
rect 576 624 588 632
rect 596 624 600 632
rect 192 614 286 622
rect 314 614 408 622
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 416 614 428 622
rect 446 614 458 622
rect 476 614 488 622
rect 506 614 518 622
rect 536 614 548 622
rect 566 614 578 622
rect 586 614 600 622
rect 0 612 600 614
rect 0 604 4 612
rect 12 604 24 612
rect 32 604 568 612
rect 576 604 588 612
rect 596 604 600 612
rect 0 602 600 604
rect 0 594 14 602
rect 22 594 34 602
rect 52 594 64 602
rect 82 594 94 602
rect 112 594 124 602
rect 142 594 154 602
rect 172 594 184 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 192 594 286 602
rect 314 594 408 602
rect 0 584 4 592
rect 12 584 24 592
rect 42 584 54 592
rect 72 584 84 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 592
rect 132 582 144 592
rect 162 582 174 592
rect 0 574 14 582
rect 22 574 34 582
rect 52 574 64 582
rect 82 574 94 582
rect 192 574 408 594
rect 416 594 428 602
rect 446 594 458 602
rect 476 594 488 602
rect 506 594 518 602
rect 536 594 548 602
rect 566 594 578 602
rect 586 594 600 602
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 426 582 438 592
rect 456 582 468 592
rect 486 582 498 592
rect 516 584 528 592
rect 546 584 558 592
rect 576 584 588 592
rect 596 584 600 592
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 506 574 518 582
rect 536 574 548 582
rect 566 574 578 582
rect 586 574 600 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 0 564 4 572
rect 12 564 24 572
rect 42 564 54 572
rect 72 564 84 572
rect 102 564 114 574
rect 132 564 144 574
rect 162 564 174 574
rect 192 566 286 574
rect 314 566 408 574
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 0 554 14 562
rect 22 554 34 562
rect 52 554 64 562
rect 82 554 94 562
rect 112 554 124 562
rect 142 554 154 562
rect 172 554 184 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 192 554 408 566
rect 426 564 438 574
rect 456 564 468 574
rect 486 564 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 516 564 528 572
rect 546 564 558 572
rect 576 564 588 572
rect 596 564 600 572
rect 0 544 4 552
rect 12 544 24 552
rect 42 544 54 552
rect 72 544 84 552
rect 102 544 114 552
rect 132 544 144 552
rect 162 544 174 552
rect 192 546 286 554
rect 314 546 408 554
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 416 554 428 562
rect 446 554 458 562
rect 476 554 488 562
rect 506 554 518 562
rect 536 554 548 562
rect 566 554 578 562
rect 586 554 600 562
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 0 534 14 542
rect 22 534 34 542
rect 52 534 64 542
rect 82 534 94 542
rect 112 534 124 542
rect 142 534 154 542
rect 172 534 184 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 192 534 408 546
rect 426 544 438 552
rect 456 544 468 552
rect 486 544 498 552
rect 516 544 528 552
rect 546 544 558 552
rect 576 544 588 552
rect 596 544 600 552
rect 0 524 4 532
rect 12 524 24 532
rect 42 524 54 532
rect 72 524 84 532
rect 102 524 114 532
rect 132 524 144 532
rect 162 524 174 532
rect 192 526 286 534
rect 314 526 408 534
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 416 534 428 542
rect 446 534 458 542
rect 476 534 488 542
rect 506 534 518 542
rect 536 534 548 542
rect 566 534 578 542
rect 586 534 600 542
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 192 524 408 526
rect 426 524 438 532
rect 456 524 468 532
rect 486 524 498 532
rect 516 524 528 532
rect 546 524 558 532
rect 576 524 588 532
rect 596 524 600 532
rect 0 516 600 524
rect 0 512 24 516
rect 0 4 4 512
rect 12 508 24 512
rect 32 508 44 516
rect 52 508 64 516
rect 72 508 84 516
rect 92 508 104 516
rect 112 508 124 516
rect 132 508 144 516
rect 152 508 164 516
rect 172 508 184 516
rect 192 514 408 516
rect 192 508 286 514
rect 12 506 286 508
rect 314 508 408 514
rect 416 508 428 516
rect 436 508 448 516
rect 456 508 468 516
rect 476 508 488 516
rect 496 508 508 516
rect 516 508 528 516
rect 536 508 548 516
rect 556 508 568 516
rect 576 512 600 516
rect 576 508 588 512
rect 314 506 588 508
rect 12 504 588 506
rect 12 16 16 504
rect 584 16 588 504
rect 12 12 588 16
rect 192 4 196 12
rect 404 4 408 12
rect 596 4 600 512
rect 0 0 600 4
<< psubstratepcontact >>
rect 2 1320 190 1338
rect 410 1320 598 1338
rect 2 840 20 1320
rect 44 836 52 844
rect 74 836 82 844
rect 104 836 112 844
rect 134 836 142 844
rect 164 836 172 844
rect 428 836 436 844
rect 458 836 466 844
rect 488 836 496 844
rect 518 836 526 844
rect 548 836 556 844
rect 580 840 598 1320
rect 4 828 12 836
rect 24 828 42 836
rect 54 828 72 836
rect 84 828 102 836
rect 114 828 132 836
rect 144 828 162 836
rect 174 828 192 836
rect 34 826 42 828
rect 64 826 72 828
rect 94 826 102 828
rect 124 826 132 828
rect 154 826 162 828
rect 14 818 22 826
rect 34 818 52 826
rect 64 818 82 826
rect 94 818 112 826
rect 124 818 142 826
rect 154 818 172 826
rect 34 816 42 818
rect 64 816 72 818
rect 94 816 102 818
rect 124 816 132 818
rect 154 816 162 818
rect 184 816 192 828
rect 286 826 314 834
rect 408 828 426 836
rect 438 828 456 836
rect 468 828 486 836
rect 498 828 516 836
rect 528 828 546 836
rect 558 828 576 836
rect 588 828 596 836
rect 4 808 12 816
rect 24 808 42 816
rect 54 808 72 816
rect 84 808 102 816
rect 114 808 132 816
rect 144 808 162 816
rect 174 808 192 816
rect 408 816 416 828
rect 438 826 446 828
rect 468 826 476 828
rect 498 826 506 828
rect 528 826 536 828
rect 558 826 566 828
rect 428 818 446 826
rect 458 818 476 826
rect 488 818 506 826
rect 518 818 536 826
rect 548 818 566 826
rect 578 818 586 826
rect 438 816 446 818
rect 468 816 476 818
rect 498 816 506 818
rect 528 816 536 818
rect 558 816 566 818
rect 34 806 42 808
rect 64 806 72 808
rect 94 806 102 808
rect 124 806 132 808
rect 154 806 162 808
rect 14 798 22 806
rect 34 798 52 806
rect 64 798 82 806
rect 94 798 112 806
rect 124 798 142 806
rect 154 798 172 806
rect 34 796 42 798
rect 64 796 72 798
rect 94 796 102 798
rect 124 796 132 798
rect 154 796 162 798
rect 184 796 192 808
rect 286 806 314 814
rect 408 808 426 816
rect 438 808 456 816
rect 468 808 486 816
rect 498 808 516 816
rect 528 808 546 816
rect 558 808 576 816
rect 588 808 596 816
rect 4 788 12 796
rect 24 788 42 796
rect 54 788 72 796
rect 84 788 102 796
rect 114 788 132 796
rect 144 788 162 796
rect 174 788 192 796
rect 408 796 416 808
rect 438 806 446 808
rect 468 806 476 808
rect 498 806 506 808
rect 528 806 536 808
rect 558 806 566 808
rect 428 798 446 806
rect 458 798 476 806
rect 488 798 506 806
rect 518 798 536 806
rect 548 798 566 806
rect 578 798 586 806
rect 438 796 446 798
rect 468 796 476 798
rect 498 796 506 798
rect 528 796 536 798
rect 558 796 566 798
rect 34 786 42 788
rect 64 786 72 788
rect 94 786 102 788
rect 124 786 132 788
rect 154 786 162 788
rect 14 778 22 786
rect 34 778 52 786
rect 64 778 82 786
rect 34 776 42 778
rect 64 776 72 778
rect 94 776 112 786
rect 124 776 142 786
rect 154 776 172 786
rect 184 776 192 788
rect 286 786 314 794
rect 408 788 426 796
rect 438 788 456 796
rect 468 788 486 796
rect 498 788 516 796
rect 528 788 546 796
rect 558 788 576 796
rect 588 788 596 796
rect 408 776 416 788
rect 438 786 446 788
rect 468 786 476 788
rect 498 786 506 788
rect 528 786 536 788
rect 558 786 566 788
rect 428 776 446 786
rect 458 776 476 786
rect 488 776 506 786
rect 518 778 536 786
rect 548 778 566 786
rect 578 778 586 786
rect 528 776 536 778
rect 558 776 566 778
rect 4 768 12 776
rect 24 768 42 776
rect 54 768 72 776
rect 84 768 192 776
rect 34 766 42 768
rect 64 766 72 768
rect 14 758 22 766
rect 34 758 52 766
rect 64 758 82 766
rect 94 758 112 768
rect 124 758 142 768
rect 154 758 172 768
rect 34 756 42 758
rect 64 756 72 758
rect 94 756 102 758
rect 124 756 132 758
rect 154 756 162 758
rect 184 756 192 768
rect 286 758 314 776
rect 408 768 516 776
rect 528 768 546 776
rect 558 768 576 776
rect 588 768 596 776
rect 4 748 12 756
rect 24 748 42 756
rect 54 748 72 756
rect 84 748 102 756
rect 114 748 132 756
rect 144 748 162 756
rect 174 748 192 756
rect 34 746 42 748
rect 64 746 72 748
rect 94 746 102 748
rect 124 746 132 748
rect 154 746 162 748
rect 14 738 22 746
rect 34 738 52 746
rect 64 738 82 746
rect 94 738 112 746
rect 124 738 142 746
rect 154 738 172 746
rect 184 738 192 748
rect 408 756 416 768
rect 428 758 446 768
rect 458 758 476 768
rect 488 758 506 768
rect 528 766 536 768
rect 558 766 566 768
rect 518 758 536 766
rect 548 758 566 766
rect 578 758 586 766
rect 438 756 446 758
rect 468 756 476 758
rect 498 756 506 758
rect 528 756 536 758
rect 558 756 566 758
rect 408 748 426 756
rect 438 748 456 756
rect 468 748 486 756
rect 498 748 516 756
rect 528 748 546 756
rect 558 748 576 756
rect 588 748 596 756
rect 286 738 314 746
rect 408 738 416 748
rect 438 746 446 748
rect 468 746 476 748
rect 498 746 506 748
rect 528 746 536 748
rect 558 746 566 748
rect 428 738 446 746
rect 458 738 476 746
rect 488 738 506 746
rect 518 738 536 746
rect 548 738 566 746
rect 578 738 586 746
rect 4 728 12 736
rect 24 728 32 736
rect 568 728 576 736
rect 588 728 596 736
rect 14 718 22 726
rect 34 718 52 726
rect 64 718 82 726
rect 94 718 112 726
rect 124 718 142 726
rect 154 718 172 726
rect 34 716 42 718
rect 64 716 72 718
rect 94 716 102 718
rect 124 716 132 718
rect 154 716 162 718
rect 184 716 192 726
rect 286 718 314 726
rect 4 708 12 716
rect 24 708 42 716
rect 54 708 72 716
rect 84 708 102 716
rect 114 708 132 716
rect 144 708 162 716
rect 174 708 192 716
rect 34 706 42 708
rect 64 706 72 708
rect 94 706 102 708
rect 124 706 132 708
rect 154 706 162 708
rect 14 698 22 706
rect 34 698 52 706
rect 64 698 82 706
rect 94 698 112 706
rect 124 698 142 706
rect 154 698 172 706
rect 34 696 42 698
rect 64 696 72 698
rect 94 696 102 698
rect 124 696 132 698
rect 154 696 162 698
rect 184 696 192 708
rect 408 716 416 726
rect 428 718 446 726
rect 458 718 476 726
rect 488 718 506 726
rect 518 718 536 726
rect 548 718 566 726
rect 578 718 586 726
rect 438 716 446 718
rect 468 716 476 718
rect 498 716 506 718
rect 528 716 536 718
rect 558 716 566 718
rect 408 708 426 716
rect 438 708 456 716
rect 468 708 486 716
rect 498 708 516 716
rect 528 708 546 716
rect 558 708 576 716
rect 588 708 596 716
rect 286 698 314 706
rect 4 688 12 696
rect 24 688 42 696
rect 54 688 72 696
rect 84 688 102 696
rect 114 688 132 696
rect 144 688 162 696
rect 174 688 192 696
rect 408 696 416 708
rect 438 706 446 708
rect 468 706 476 708
rect 498 706 506 708
rect 528 706 536 708
rect 558 706 566 708
rect 428 698 446 706
rect 458 698 476 706
rect 488 698 506 706
rect 518 698 536 706
rect 548 698 566 706
rect 578 698 586 706
rect 438 696 446 698
rect 468 696 476 698
rect 498 696 506 698
rect 528 696 536 698
rect 558 696 566 698
rect 408 688 426 696
rect 438 688 456 696
rect 468 688 486 696
rect 498 688 516 696
rect 528 688 546 696
rect 558 688 576 696
rect 588 688 596 696
rect 36 466 74 484
rect 36 454 54 462
rect 36 434 54 442
rect 82 456 190 484
rect 286 458 314 486
rect 416 466 564 474
rect 36 414 54 422
rect 36 394 54 402
rect 36 374 54 382
rect 36 354 54 362
rect 36 334 54 342
rect 36 314 54 322
rect 36 294 54 302
rect 36 274 54 282
rect 36 254 54 262
rect 36 234 54 242
rect 36 214 54 222
rect 36 194 54 202
rect 36 174 54 182
rect 36 154 54 162
rect 36 134 54 142
rect 36 114 54 122
rect 36 94 54 102
rect 416 456 504 466
rect 546 454 564 462
rect 291 392 309 400
rect 291 376 309 384
rect 291 264 309 272
rect 291 248 309 256
rect 291 136 309 144
rect 291 120 309 128
rect 291 104 309 112
rect 291 88 309 96
rect 36 74 54 82
rect 36 54 54 62
rect 36 34 84 42
rect 88 34 96 62
rect 108 34 116 62
rect 128 34 136 62
rect 148 34 156 62
rect 168 34 176 62
rect 188 34 196 62
rect 546 434 564 442
rect 546 414 564 422
rect 546 394 564 402
rect 546 374 564 382
rect 546 354 564 362
rect 546 334 564 342
rect 546 314 564 322
rect 546 294 564 302
rect 546 274 564 282
rect 546 254 564 262
rect 546 234 564 242
rect 546 214 564 222
rect 546 194 564 202
rect 546 174 564 182
rect 546 154 564 162
rect 546 134 564 142
rect 546 114 564 122
rect 546 94 564 102
rect 404 34 412 62
rect 424 34 432 62
rect 444 34 452 62
rect 464 34 472 62
rect 484 34 492 62
rect 504 34 512 62
rect 546 74 564 82
rect 546 54 564 62
rect 516 34 564 42
<< nsubstratencontact >>
rect 51 1290 59 1298
rect 72 1294 80 1298
rect 520 1294 528 1298
rect 72 1290 90 1294
rect 41 1280 49 1288
rect 62 1281 70 1289
rect 82 1286 90 1290
rect 102 1286 110 1294
rect 122 1286 130 1294
rect 142 1286 150 1294
rect 162 1286 170 1294
rect 182 1286 190 1294
rect 202 1286 210 1294
rect 222 1286 230 1294
rect 370 1286 378 1294
rect 390 1286 398 1294
rect 410 1286 418 1294
rect 430 1286 438 1294
rect 450 1286 458 1294
rect 470 1286 478 1294
rect 490 1286 498 1294
rect 510 1290 528 1294
rect 541 1290 549 1298
rect 510 1286 518 1290
rect 51 1270 59 1278
rect 41 1260 49 1268
rect 92 1276 100 1284
rect 112 1276 120 1284
rect 132 1276 140 1284
rect 152 1276 160 1284
rect 172 1276 180 1284
rect 192 1276 200 1284
rect 212 1276 220 1284
rect 232 1276 240 1284
rect 51 1250 59 1258
rect 41 1240 49 1248
rect 51 1230 59 1238
rect 41 1220 49 1228
rect 51 1210 59 1218
rect 41 1200 49 1208
rect 51 1190 59 1198
rect 41 1180 49 1188
rect 51 1170 59 1178
rect 41 1160 49 1168
rect 51 1150 59 1158
rect 41 1140 49 1148
rect 51 1130 59 1138
rect 41 1120 49 1128
rect 51 1110 59 1118
rect 41 1100 49 1108
rect 51 1090 59 1098
rect 41 1080 49 1088
rect 51 1070 59 1078
rect 41 1060 49 1068
rect 51 1050 59 1058
rect 41 1040 49 1048
rect 51 1030 59 1038
rect 41 1020 49 1028
rect 51 1010 59 1018
rect 41 1000 49 1008
rect 51 990 59 998
rect 41 980 49 988
rect 51 970 59 978
rect 41 960 49 968
rect 51 950 59 958
rect 41 940 49 948
rect 51 930 59 938
rect 41 920 49 928
rect 51 910 59 918
rect 41 900 49 908
rect 360 1276 368 1284
rect 380 1276 388 1284
rect 400 1276 408 1284
rect 420 1276 428 1284
rect 440 1276 448 1284
rect 460 1276 468 1284
rect 480 1276 488 1284
rect 500 1276 508 1284
rect 530 1281 538 1289
rect 551 1280 559 1288
rect 541 1270 549 1278
rect 551 1260 559 1268
rect 291 1218 309 1226
rect 291 1202 309 1210
rect 291 1090 309 1098
rect 291 1074 309 1082
rect 51 890 59 898
rect 41 880 49 888
rect 541 1250 549 1258
rect 551 1240 559 1248
rect 541 1230 549 1238
rect 551 1220 559 1228
rect 541 1210 549 1218
rect 551 1200 559 1208
rect 541 1190 549 1198
rect 551 1180 559 1188
rect 541 1170 549 1178
rect 551 1160 559 1168
rect 541 1150 549 1158
rect 551 1140 559 1148
rect 541 1130 549 1138
rect 551 1120 559 1128
rect 541 1110 549 1118
rect 551 1100 559 1108
rect 541 1090 549 1098
rect 551 1080 559 1088
rect 541 1070 549 1078
rect 551 1060 559 1068
rect 541 1050 549 1058
rect 551 1040 559 1048
rect 541 1030 549 1038
rect 551 1020 559 1028
rect 541 1010 549 1018
rect 551 1000 559 1008
rect 541 990 549 998
rect 551 980 559 988
rect 541 970 549 978
rect 551 960 559 968
rect 541 950 549 958
rect 551 940 559 948
rect 541 930 549 938
rect 551 920 559 928
rect 541 910 549 918
rect 551 900 559 908
rect 541 890 549 898
rect 62 873 190 883
rect 42 865 190 873
rect 286 865 314 883
rect 410 873 538 883
rect 551 880 559 888
rect 410 865 558 873
rect 4 644 12 652
rect 24 644 42 652
rect 54 644 72 652
rect 84 644 102 652
rect 114 644 132 652
rect 144 644 162 652
rect 174 644 192 652
rect 34 642 42 644
rect 64 642 72 644
rect 94 642 102 644
rect 124 642 132 644
rect 154 642 162 644
rect 14 634 22 642
rect 34 634 52 642
rect 64 634 82 642
rect 94 634 112 642
rect 124 634 142 642
rect 154 634 172 642
rect 34 632 42 634
rect 64 632 72 634
rect 94 632 102 634
rect 124 632 132 634
rect 154 632 162 634
rect 184 632 192 644
rect 408 644 426 652
rect 438 644 456 652
rect 468 644 486 652
rect 498 644 516 652
rect 528 644 546 652
rect 558 644 576 652
rect 588 644 596 652
rect 286 634 314 642
rect 4 624 12 632
rect 24 624 42 632
rect 54 624 72 632
rect 84 624 102 632
rect 114 624 132 632
rect 144 624 162 632
rect 174 624 192 632
rect 34 622 42 624
rect 64 622 72 624
rect 94 622 102 624
rect 124 622 132 624
rect 154 622 162 624
rect 14 614 22 622
rect 34 614 52 622
rect 64 614 82 622
rect 94 614 112 622
rect 124 614 142 622
rect 154 614 172 622
rect 184 614 192 624
rect 408 632 416 644
rect 438 642 446 644
rect 468 642 476 644
rect 498 642 506 644
rect 528 642 536 644
rect 558 642 566 644
rect 428 634 446 642
rect 458 634 476 642
rect 488 634 506 642
rect 518 634 536 642
rect 548 634 566 642
rect 578 634 586 642
rect 438 632 446 634
rect 468 632 476 634
rect 498 632 506 634
rect 528 632 536 634
rect 558 632 566 634
rect 408 624 426 632
rect 438 624 456 632
rect 468 624 486 632
rect 498 624 516 632
rect 528 624 546 632
rect 558 624 576 632
rect 588 624 596 632
rect 286 614 314 622
rect 408 614 416 624
rect 438 622 446 624
rect 468 622 476 624
rect 498 622 506 624
rect 528 622 536 624
rect 558 622 566 624
rect 428 614 446 622
rect 458 614 476 622
rect 488 614 506 622
rect 518 614 536 622
rect 548 614 566 622
rect 578 614 586 622
rect 4 604 12 612
rect 24 604 32 612
rect 568 604 576 612
rect 588 604 596 612
rect 14 594 22 602
rect 34 594 52 602
rect 64 594 82 602
rect 94 594 112 602
rect 124 594 142 602
rect 154 594 172 602
rect 34 592 42 594
rect 64 592 72 594
rect 94 592 102 594
rect 124 592 132 594
rect 154 592 162 594
rect 184 592 192 602
rect 286 594 314 602
rect 4 584 12 592
rect 24 584 42 592
rect 54 584 72 592
rect 84 584 102 592
rect 34 582 42 584
rect 64 582 72 584
rect 94 582 102 584
rect 114 582 132 592
rect 144 582 162 592
rect 174 582 192 592
rect 14 574 22 582
rect 34 574 52 582
rect 64 574 82 582
rect 94 574 192 582
rect 408 592 416 602
rect 428 594 446 602
rect 458 594 476 602
rect 488 594 506 602
rect 518 594 536 602
rect 548 594 566 602
rect 578 594 586 602
rect 438 592 446 594
rect 468 592 476 594
rect 498 592 506 594
rect 528 592 536 594
rect 558 592 566 594
rect 408 582 426 592
rect 438 582 456 592
rect 468 582 486 592
rect 498 584 516 592
rect 528 584 546 592
rect 558 584 576 592
rect 588 584 596 592
rect 498 582 506 584
rect 528 582 536 584
rect 558 582 566 584
rect 408 574 506 582
rect 518 574 536 582
rect 548 574 566 582
rect 578 574 586 582
rect 34 572 42 574
rect 64 572 72 574
rect 94 572 102 574
rect 4 564 12 572
rect 24 564 42 572
rect 54 564 72 572
rect 84 564 102 572
rect 114 564 132 574
rect 144 564 162 574
rect 174 564 192 574
rect 286 566 314 574
rect 34 562 42 564
rect 64 562 72 564
rect 94 562 102 564
rect 124 562 132 564
rect 154 562 162 564
rect 14 554 22 562
rect 34 554 52 562
rect 64 554 82 562
rect 94 554 112 562
rect 124 554 142 562
rect 154 554 172 562
rect 34 552 42 554
rect 64 552 72 554
rect 94 552 102 554
rect 124 552 132 554
rect 154 552 162 554
rect 184 552 192 564
rect 408 564 426 574
rect 438 564 456 574
rect 468 564 486 574
rect 498 572 506 574
rect 528 572 536 574
rect 558 572 566 574
rect 498 564 516 572
rect 528 564 546 572
rect 558 564 576 572
rect 588 564 596 572
rect 4 544 12 552
rect 24 544 42 552
rect 54 544 72 552
rect 84 544 102 552
rect 114 544 132 552
rect 144 544 162 552
rect 174 544 192 552
rect 286 546 314 554
rect 408 552 416 564
rect 438 562 446 564
rect 468 562 476 564
rect 498 562 506 564
rect 528 562 536 564
rect 558 562 566 564
rect 428 554 446 562
rect 458 554 476 562
rect 488 554 506 562
rect 518 554 536 562
rect 548 554 566 562
rect 578 554 586 562
rect 438 552 446 554
rect 468 552 476 554
rect 498 552 506 554
rect 528 552 536 554
rect 558 552 566 554
rect 34 542 42 544
rect 64 542 72 544
rect 94 542 102 544
rect 124 542 132 544
rect 154 542 162 544
rect 14 534 22 542
rect 34 534 52 542
rect 64 534 82 542
rect 94 534 112 542
rect 124 534 142 542
rect 154 534 172 542
rect 34 532 42 534
rect 64 532 72 534
rect 94 532 102 534
rect 124 532 132 534
rect 154 532 162 534
rect 184 532 192 544
rect 408 544 426 552
rect 438 544 456 552
rect 468 544 486 552
rect 498 544 516 552
rect 528 544 546 552
rect 558 544 576 552
rect 588 544 596 552
rect 4 524 12 532
rect 24 524 42 532
rect 54 524 72 532
rect 84 524 102 532
rect 114 524 132 532
rect 144 524 162 532
rect 174 524 192 532
rect 286 526 314 534
rect 408 532 416 544
rect 438 542 446 544
rect 468 542 476 544
rect 498 542 506 544
rect 528 542 536 544
rect 558 542 566 544
rect 428 534 446 542
rect 458 534 476 542
rect 488 534 506 542
rect 518 534 536 542
rect 548 534 566 542
rect 578 534 586 542
rect 438 532 446 534
rect 468 532 476 534
rect 498 532 506 534
rect 528 532 536 534
rect 558 532 566 534
rect 408 524 426 532
rect 438 524 456 532
rect 468 524 486 532
rect 498 524 516 532
rect 528 524 546 532
rect 558 524 576 532
rect 588 524 596 532
rect 4 12 12 512
rect 24 508 32 516
rect 44 508 52 516
rect 64 508 72 516
rect 84 508 92 516
rect 104 508 112 516
rect 124 508 132 516
rect 144 508 152 516
rect 164 508 172 516
rect 184 508 192 516
rect 286 506 314 514
rect 408 508 416 516
rect 428 508 436 516
rect 448 508 456 516
rect 468 508 476 516
rect 488 508 496 516
rect 508 508 516 516
rect 528 508 536 516
rect 548 508 556 516
rect 568 508 576 516
rect 588 12 596 512
rect 4 4 192 12
rect 196 4 404 12
rect 408 4 596 12
<< polysilicon >>
rect 62 1252 76 1258
rect 276 1252 280 1258
rect 62 914 64 1252
rect 72 1170 74 1252
rect 320 1252 324 1258
rect 524 1252 538 1258
rect 72 1164 76 1170
rect 276 1164 280 1170
rect 72 1130 74 1164
rect 72 1124 76 1130
rect 276 1124 280 1130
rect 72 1042 74 1124
rect 526 1170 528 1252
rect 320 1164 324 1170
rect 524 1164 528 1170
rect 526 1130 528 1164
rect 320 1124 324 1130
rect 524 1124 528 1130
rect 72 1036 76 1042
rect 276 1036 280 1042
rect 72 1000 74 1036
rect 72 994 76 1000
rect 276 994 280 1000
rect 72 914 74 994
rect 62 912 74 914
rect 62 906 76 912
rect 276 906 280 912
rect 526 1042 528 1124
rect 320 1036 324 1042
rect 524 1036 528 1042
rect 526 1000 528 1036
rect 320 994 324 1000
rect 524 994 528 1000
rect 526 914 528 994
rect 536 914 538 1252
rect 526 912 538 914
rect 320 906 324 912
rect 524 906 538 912
rect 62 434 76 438
rect 62 86 64 434
rect 72 432 76 434
rect 276 432 280 438
rect 72 348 74 432
rect 320 432 324 438
rect 524 434 538 438
rect 524 432 528 434
rect 72 342 76 348
rect 276 342 280 348
rect 72 306 74 342
rect 72 300 76 306
rect 276 300 280 306
rect 72 218 74 300
rect 526 348 528 432
rect 320 342 324 348
rect 524 342 528 348
rect 526 306 528 342
rect 320 300 324 306
rect 524 300 528 306
rect 72 212 76 218
rect 276 212 280 218
rect 72 176 74 212
rect 72 170 76 176
rect 276 170 280 176
rect 72 88 74 170
rect 526 218 528 300
rect 320 212 324 218
rect 524 212 528 218
rect 526 176 528 212
rect 320 170 324 176
rect 524 170 528 176
rect 526 88 528 170
rect 72 86 76 88
rect 62 82 76 86
rect 276 82 280 88
rect 320 82 324 88
rect 524 86 528 88
rect 536 86 538 434
rect 524 82 538 86
<< polycontact >>
rect 64 914 72 1252
rect 528 914 536 1252
rect 64 86 72 434
rect 528 86 536 434
<< metal1 >>
rect 124 1460 476 1480
rect 144 1440 456 1460
rect 164 1420 436 1440
rect 184 1400 416 1420
rect 0 1338 198 1340
rect 0 840 2 1338
rect 190 1320 198 1338
rect 20 1318 198 1320
rect 20 846 22 1318
rect 204 1306 396 1400
rect 402 1338 600 1340
rect 402 1320 410 1338
rect 402 1318 580 1320
rect 40 1298 240 1300
rect 40 1290 42 1298
rect 50 1290 51 1298
rect 59 1290 62 1298
rect 70 1290 72 1298
rect 80 1294 240 1298
rect 40 1289 72 1290
rect 40 1288 62 1289
rect 40 1280 41 1288
rect 49 1287 62 1288
rect 49 1280 50 1287
rect 40 1279 50 1280
rect 58 1281 62 1287
rect 70 1282 72 1289
rect 80 1286 82 1290
rect 90 1286 92 1294
rect 100 1286 102 1294
rect 110 1286 112 1294
rect 120 1286 122 1294
rect 130 1286 132 1294
rect 140 1286 142 1294
rect 150 1286 152 1294
rect 160 1286 162 1294
rect 170 1286 172 1294
rect 180 1286 182 1294
rect 190 1286 192 1294
rect 200 1286 202 1294
rect 210 1286 212 1294
rect 220 1286 222 1294
rect 230 1286 232 1294
rect 80 1284 240 1286
rect 70 1281 82 1282
rect 58 1279 82 1281
rect 40 1278 82 1279
rect 40 1270 42 1278
rect 50 1270 51 1278
rect 59 1276 82 1278
rect 90 1276 92 1284
rect 100 1276 102 1284
rect 110 1276 112 1284
rect 120 1276 122 1284
rect 130 1276 132 1284
rect 140 1276 142 1284
rect 150 1276 152 1284
rect 160 1276 162 1284
rect 170 1276 172 1284
rect 180 1276 182 1284
rect 190 1276 192 1284
rect 200 1276 202 1284
rect 210 1276 212 1284
rect 220 1276 222 1284
rect 230 1276 232 1284
rect 59 1274 240 1276
rect 59 1270 82 1274
rect 40 1268 82 1270
rect 40 1260 41 1268
rect 49 1267 82 1268
rect 49 1260 50 1267
rect 40 1259 50 1260
rect 58 1266 82 1267
rect 58 1259 240 1266
rect 40 1258 240 1259
rect 40 1250 42 1258
rect 50 1250 51 1258
rect 59 1252 240 1258
rect 59 1250 64 1252
rect 40 1248 64 1250
rect 40 1240 41 1248
rect 49 1247 64 1248
rect 49 1240 50 1247
rect 40 1239 50 1240
rect 58 1239 64 1247
rect 40 1238 64 1239
rect 40 1230 42 1238
rect 50 1230 51 1238
rect 59 1230 64 1238
rect 40 1228 64 1230
rect 40 1220 41 1228
rect 49 1227 64 1228
rect 49 1220 50 1227
rect 40 1219 50 1220
rect 58 1219 64 1227
rect 40 1218 64 1219
rect 40 1210 42 1218
rect 50 1210 51 1218
rect 59 1210 64 1218
rect 40 1208 64 1210
rect 40 1200 41 1208
rect 49 1207 64 1208
rect 49 1200 50 1207
rect 40 1199 50 1200
rect 58 1199 64 1207
rect 40 1198 64 1199
rect 40 1190 42 1198
rect 50 1190 51 1198
rect 59 1190 64 1198
rect 40 1188 64 1190
rect 40 1180 41 1188
rect 49 1187 64 1188
rect 49 1180 50 1187
rect 40 1179 50 1180
rect 58 1179 64 1187
rect 40 1178 64 1179
rect 40 1170 42 1178
rect 50 1170 51 1178
rect 59 1170 64 1178
rect 40 1168 64 1170
rect 40 1160 41 1168
rect 49 1167 64 1168
rect 49 1160 50 1167
rect 40 1159 50 1160
rect 58 1159 64 1167
rect 40 1158 64 1159
rect 40 1150 42 1158
rect 50 1150 51 1158
rect 59 1150 64 1158
rect 40 1148 64 1150
rect 40 1140 41 1148
rect 49 1147 64 1148
rect 49 1140 50 1147
rect 40 1139 50 1140
rect 58 1139 64 1147
rect 40 1138 64 1139
rect 40 1130 42 1138
rect 50 1130 51 1138
rect 59 1130 64 1138
rect 40 1128 64 1130
rect 40 1120 41 1128
rect 49 1127 64 1128
rect 49 1120 50 1127
rect 40 1119 50 1120
rect 58 1119 64 1127
rect 40 1118 64 1119
rect 40 1110 42 1118
rect 50 1110 51 1118
rect 59 1110 64 1118
rect 40 1108 64 1110
rect 40 1100 41 1108
rect 49 1107 64 1108
rect 49 1100 50 1107
rect 40 1099 50 1100
rect 58 1099 64 1107
rect 40 1098 64 1099
rect 40 1090 42 1098
rect 50 1090 51 1098
rect 59 1090 64 1098
rect 40 1088 64 1090
rect 40 1080 41 1088
rect 49 1087 64 1088
rect 49 1080 50 1087
rect 40 1079 50 1080
rect 58 1079 64 1087
rect 40 1078 64 1079
rect 40 1070 42 1078
rect 50 1070 51 1078
rect 59 1070 64 1078
rect 40 1068 64 1070
rect 40 1060 41 1068
rect 49 1067 64 1068
rect 49 1060 50 1067
rect 40 1059 50 1060
rect 58 1059 64 1067
rect 40 1058 64 1059
rect 40 1050 42 1058
rect 50 1050 51 1058
rect 59 1050 64 1058
rect 40 1048 64 1050
rect 40 1040 41 1048
rect 49 1047 64 1048
rect 49 1040 50 1047
rect 40 1039 50 1040
rect 58 1039 64 1047
rect 40 1038 64 1039
rect 40 1030 42 1038
rect 50 1030 51 1038
rect 59 1030 64 1038
rect 40 1028 64 1030
rect 40 1020 41 1028
rect 49 1027 64 1028
rect 49 1020 50 1027
rect 40 1019 50 1020
rect 58 1019 64 1027
rect 40 1018 64 1019
rect 40 1010 42 1018
rect 50 1010 51 1018
rect 59 1010 64 1018
rect 40 1008 64 1010
rect 40 1000 41 1008
rect 49 1007 64 1008
rect 49 1000 50 1007
rect 40 999 50 1000
rect 58 999 64 1007
rect 40 998 64 999
rect 40 990 42 998
rect 50 990 51 998
rect 59 990 64 998
rect 40 988 64 990
rect 40 980 41 988
rect 49 987 64 988
rect 49 980 50 987
rect 40 979 50 980
rect 58 979 64 987
rect 40 978 64 979
rect 40 970 42 978
rect 50 970 51 978
rect 59 970 64 978
rect 40 968 64 970
rect 40 960 41 968
rect 49 967 64 968
rect 49 960 50 967
rect 40 959 50 960
rect 58 959 64 967
rect 40 958 64 959
rect 40 950 42 958
rect 50 950 51 958
rect 59 950 64 958
rect 40 948 64 950
rect 40 940 41 948
rect 49 947 64 948
rect 49 940 50 947
rect 40 939 50 940
rect 58 939 64 947
rect 40 938 64 939
rect 40 930 42 938
rect 50 930 51 938
rect 59 930 64 938
rect 40 928 64 930
rect 40 920 41 928
rect 49 927 64 928
rect 49 920 50 927
rect 40 919 50 920
rect 58 919 64 927
rect 40 918 64 919
rect 40 910 42 918
rect 50 910 51 918
rect 59 914 64 918
rect 72 1250 240 1252
rect 72 1172 78 1250
rect 236 1242 240 1250
rect 96 1180 102 1242
rect 246 1236 354 1306
rect 360 1298 528 1300
rect 360 1294 520 1298
rect 368 1286 370 1294
rect 378 1286 380 1294
rect 388 1286 390 1294
rect 398 1286 400 1294
rect 408 1286 410 1294
rect 418 1286 420 1294
rect 428 1286 430 1294
rect 438 1286 440 1294
rect 448 1286 450 1294
rect 458 1286 460 1294
rect 468 1286 470 1294
rect 478 1286 480 1294
rect 488 1286 490 1294
rect 498 1286 500 1294
rect 508 1286 510 1294
rect 528 1290 530 1298
rect 538 1290 541 1298
rect 549 1290 550 1298
rect 558 1290 560 1298
rect 518 1286 520 1290
rect 360 1284 520 1286
rect 528 1289 560 1290
rect 368 1276 370 1284
rect 378 1276 380 1284
rect 388 1276 390 1284
rect 398 1276 400 1284
rect 408 1276 410 1284
rect 418 1276 420 1284
rect 428 1276 430 1284
rect 438 1276 440 1284
rect 448 1276 450 1284
rect 458 1276 460 1284
rect 468 1276 470 1284
rect 478 1276 480 1284
rect 488 1276 490 1284
rect 498 1276 500 1284
rect 508 1276 510 1284
rect 528 1282 530 1289
rect 518 1281 530 1282
rect 538 1288 560 1289
rect 538 1287 551 1288
rect 538 1281 542 1287
rect 518 1279 542 1281
rect 550 1280 551 1287
rect 559 1280 560 1288
rect 550 1279 560 1280
rect 518 1278 560 1279
rect 518 1276 541 1278
rect 360 1274 541 1276
rect 518 1270 541 1274
rect 549 1270 550 1278
rect 558 1270 560 1278
rect 518 1268 560 1270
rect 518 1267 551 1268
rect 518 1266 542 1267
rect 360 1259 542 1266
rect 550 1260 551 1267
rect 559 1260 560 1268
rect 550 1259 560 1260
rect 360 1258 560 1259
rect 360 1252 541 1258
rect 360 1250 528 1252
rect 360 1242 364 1250
rect 112 1232 488 1236
rect 112 1220 285 1232
rect 240 1202 285 1220
rect 315 1220 488 1232
rect 315 1202 360 1220
rect 112 1196 285 1202
rect 315 1196 488 1202
rect 112 1186 488 1196
rect 236 1172 240 1180
rect 72 1156 240 1172
rect 72 1138 82 1156
rect 72 1122 240 1138
rect 72 1044 78 1122
rect 236 1114 240 1122
rect 96 1052 102 1114
rect 246 1108 354 1186
rect 498 1180 504 1242
rect 360 1172 364 1180
rect 522 1172 528 1250
rect 360 1156 528 1172
rect 518 1138 528 1156
rect 360 1122 528 1138
rect 360 1114 364 1122
rect 112 1104 488 1108
rect 112 1092 285 1104
rect 240 1074 285 1092
rect 315 1092 488 1104
rect 315 1074 360 1092
rect 112 1068 285 1074
rect 315 1068 488 1074
rect 112 1058 488 1068
rect 236 1044 240 1052
rect 72 1028 240 1044
rect 72 1020 82 1028
rect 72 1016 240 1020
rect 72 1008 82 1016
rect 72 992 240 1008
rect 72 914 78 992
rect 236 984 240 992
rect 96 922 102 984
rect 246 978 354 1058
rect 498 1052 504 1114
rect 360 1044 364 1052
rect 522 1044 528 1122
rect 360 1028 528 1044
rect 518 1020 528 1028
rect 360 1016 528 1020
rect 518 1008 528 1016
rect 360 992 528 1008
rect 360 984 364 992
rect 112 962 488 978
rect 240 944 360 962
rect 112 928 488 944
rect 196 914 198 922
rect 59 910 198 914
rect 40 908 198 910
rect 40 900 41 908
rect 49 907 198 908
rect 49 900 50 907
rect 40 899 50 900
rect 58 899 198 907
rect 40 898 198 899
rect 40 890 42 898
rect 50 890 51 898
rect 59 890 82 898
rect 190 890 198 898
rect 40 888 198 890
rect 40 880 41 888
rect 49 880 50 888
rect 58 883 198 888
rect 58 880 62 883
rect 40 873 62 880
rect 40 865 42 873
rect 190 865 198 883
rect 204 909 396 928
rect 498 922 504 984
rect 20 844 198 846
rect 20 840 24 844
rect 0 836 24 840
rect 0 828 4 836
rect 12 828 14 836
rect 22 828 24 836
rect 42 828 44 844
rect 52 828 54 844
rect 72 828 74 844
rect 82 828 84 844
rect 102 828 104 844
rect 112 828 114 844
rect 132 828 134 844
rect 142 828 144 844
rect 162 828 164 844
rect 172 828 174 844
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 184 828
rect 0 818 4 826
rect 12 818 14 826
rect 22 818 24 826
rect 32 818 34 826
rect 52 818 54 826
rect 62 818 64 826
rect 82 818 84 826
rect 92 818 94 826
rect 112 818 114 826
rect 122 818 124 826
rect 142 818 144 826
rect 152 818 154 826
rect 172 818 174 826
rect 182 818 184 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 184 818
rect 0 808 4 816
rect 12 808 14 816
rect 22 808 24 816
rect 42 808 44 816
rect 52 808 54 816
rect 72 808 74 816
rect 82 808 84 816
rect 102 808 104 816
rect 112 808 114 816
rect 132 808 134 816
rect 142 808 144 816
rect 162 808 164 816
rect 172 808 174 816
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 184 808
rect 0 798 4 806
rect 12 798 14 806
rect 22 798 24 806
rect 32 798 34 806
rect 52 798 54 806
rect 62 798 64 806
rect 82 798 84 806
rect 92 798 94 806
rect 112 798 114 806
rect 122 798 124 806
rect 142 798 144 806
rect 152 798 154 806
rect 172 798 174 806
rect 182 798 184 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 184 798
rect 0 788 4 796
rect 12 788 14 796
rect 22 788 24 796
rect 42 788 44 796
rect 52 788 54 796
rect 72 788 74 796
rect 82 788 84 796
rect 102 788 104 796
rect 112 788 114 796
rect 132 788 134 796
rect 142 788 144 796
rect 162 788 164 796
rect 172 788 174 796
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 184 788
rect 0 778 4 786
rect 12 778 14 786
rect 22 778 24 786
rect 32 778 34 786
rect 52 778 54 786
rect 62 778 64 786
rect 82 778 84 786
rect 92 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 778 114 786
rect 122 778 124 786
rect 112 776 124 778
rect 142 778 144 786
rect 152 778 154 786
rect 142 776 154 778
rect 172 778 174 786
rect 182 778 184 786
rect 172 776 184 778
rect 0 768 4 776
rect 12 768 14 776
rect 22 768 24 776
rect 42 768 44 776
rect 52 768 54 776
rect 72 768 74 776
rect 82 768 84 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 4 766
rect 12 758 14 766
rect 22 758 24 766
rect 32 758 34 766
rect 52 758 54 766
rect 62 758 64 766
rect 82 758 84 766
rect 92 758 94 766
rect 112 766 124 768
rect 112 758 114 766
rect 122 758 124 766
rect 142 766 154 768
rect 142 758 144 766
rect 152 758 154 766
rect 172 766 184 768
rect 172 758 174 766
rect 182 758 184 766
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 184 758
rect 0 748 4 756
rect 12 748 14 756
rect 22 748 24 756
rect 42 748 44 756
rect 52 748 54 756
rect 72 748 74 756
rect 82 748 84 756
rect 102 748 104 756
rect 112 748 114 756
rect 132 748 134 756
rect 142 748 144 756
rect 162 748 164 756
rect 172 748 174 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 184 748
rect 0 738 4 746
rect 12 738 14 746
rect 22 738 24 746
rect 32 738 34 746
rect 52 738 54 746
rect 62 738 64 746
rect 82 738 84 746
rect 92 738 94 746
rect 112 738 114 746
rect 122 738 124 746
rect 142 738 144 746
rect 152 738 154 746
rect 172 738 174 746
rect 182 738 184 746
rect 192 738 198 844
rect 0 737 198 738
rect 0 736 42 737
rect 0 728 4 736
rect 12 728 14 736
rect 22 728 24 736
rect 32 728 42 736
rect 0 727 42 728
rect 0 726 198 727
rect 0 718 4 726
rect 12 718 14 726
rect 22 718 24 726
rect 32 718 34 726
rect 52 718 54 726
rect 62 718 64 726
rect 82 718 84 726
rect 92 718 94 726
rect 112 718 114 726
rect 122 718 124 726
rect 142 718 144 726
rect 152 718 154 726
rect 172 718 174 726
rect 182 718 184 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 184 718
rect 0 708 4 716
rect 12 708 14 716
rect 22 708 24 716
rect 42 708 44 716
rect 52 708 54 716
rect 72 708 74 716
rect 82 708 84 716
rect 102 708 104 716
rect 112 708 114 716
rect 132 708 134 716
rect 142 708 144 716
rect 162 708 164 716
rect 172 708 174 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 184 708
rect 0 698 4 706
rect 12 698 14 706
rect 22 698 24 706
rect 32 698 34 706
rect 52 698 54 706
rect 62 698 64 706
rect 82 698 84 706
rect 92 698 94 706
rect 112 698 114 706
rect 122 698 124 706
rect 142 698 144 706
rect 152 698 154 706
rect 172 698 174 706
rect 182 698 184 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 184 698
rect 0 688 4 696
rect 12 688 14 696
rect 22 688 24 696
rect 42 688 44 696
rect 52 688 54 696
rect 72 688 74 696
rect 82 688 84 696
rect 102 688 104 696
rect 112 688 114 696
rect 132 688 134 696
rect 142 688 144 696
rect 162 688 164 696
rect 172 688 174 696
rect 192 688 198 726
rect 0 644 4 652
rect 12 644 14 652
rect 22 644 24 652
rect 42 644 44 652
rect 52 644 54 652
rect 72 644 74 652
rect 82 644 84 652
rect 102 644 104 652
rect 112 644 114 652
rect 132 644 134 652
rect 142 644 144 652
rect 162 644 164 652
rect 172 644 174 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 0 634 4 642
rect 12 634 14 642
rect 22 634 24 642
rect 32 634 34 642
rect 52 634 54 642
rect 62 634 64 642
rect 82 634 84 642
rect 92 634 94 642
rect 112 634 114 642
rect 122 634 124 642
rect 142 634 144 642
rect 152 634 154 642
rect 172 634 174 642
rect 182 634 184 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 0 624 4 632
rect 12 624 14 632
rect 22 624 24 632
rect 42 624 44 632
rect 52 624 54 632
rect 72 624 74 632
rect 82 624 84 632
rect 102 624 104 632
rect 112 624 114 632
rect 132 624 134 632
rect 142 624 144 632
rect 162 624 164 632
rect 172 624 174 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 0 614 4 622
rect 12 614 14 622
rect 22 614 24 622
rect 32 614 34 622
rect 52 614 54 622
rect 62 614 64 622
rect 82 614 84 622
rect 92 614 94 622
rect 112 614 114 622
rect 122 614 124 622
rect 142 614 144 622
rect 152 614 154 622
rect 172 614 174 622
rect 182 614 184 622
rect 192 614 198 652
rect 0 612 198 614
rect 0 604 4 612
rect 12 604 14 612
rect 22 604 24 612
rect 32 604 40 612
rect 0 602 40 604
rect 0 594 4 602
rect 12 594 14 602
rect 22 594 24 602
rect 32 594 34 602
rect 52 594 54 602
rect 62 594 64 602
rect 82 594 84 602
rect 92 594 94 602
rect 112 594 114 602
rect 122 594 124 602
rect 142 594 144 602
rect 152 594 154 602
rect 172 594 174 602
rect 182 594 184 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 0 584 4 592
rect 12 584 14 592
rect 22 584 24 592
rect 42 584 44 592
rect 52 584 54 592
rect 72 584 74 592
rect 82 584 84 592
rect 102 584 104 592
rect 112 584 114 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 584
rect 132 584 134 592
rect 142 584 144 592
rect 132 582 144 584
rect 162 584 164 592
rect 172 584 174 592
rect 162 582 174 584
rect 0 574 4 582
rect 12 574 14 582
rect 22 574 24 582
rect 32 574 34 582
rect 52 574 54 582
rect 62 574 64 582
rect 82 574 84 582
rect 92 574 94 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 102 572 114 574
rect 0 564 4 572
rect 12 564 14 572
rect 22 564 24 572
rect 42 564 44 572
rect 52 564 54 572
rect 72 564 74 572
rect 82 564 84 572
rect 102 564 104 572
rect 112 564 114 572
rect 132 572 144 574
rect 132 564 134 572
rect 142 564 144 572
rect 162 572 174 574
rect 162 564 164 572
rect 172 564 174 572
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 0 554 4 562
rect 12 554 14 562
rect 22 554 24 562
rect 32 554 34 562
rect 52 554 54 562
rect 62 554 64 562
rect 82 554 84 562
rect 92 554 94 562
rect 112 554 114 562
rect 122 554 124 562
rect 142 554 144 562
rect 152 554 154 562
rect 172 554 174 562
rect 182 554 184 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 0 544 4 552
rect 12 544 14 552
rect 22 544 24 552
rect 42 544 44 552
rect 52 544 54 552
rect 72 544 74 552
rect 82 544 84 552
rect 102 544 104 552
rect 112 544 114 552
rect 132 544 134 552
rect 142 544 144 552
rect 162 544 164 552
rect 172 544 174 552
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 0 534 4 542
rect 12 534 14 542
rect 22 534 24 542
rect 32 534 34 542
rect 52 534 54 542
rect 62 534 64 542
rect 82 534 84 542
rect 92 534 94 542
rect 112 534 114 542
rect 122 534 124 542
rect 142 534 144 542
rect 152 534 154 542
rect 172 534 174 542
rect 182 534 184 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 0 524 4 532
rect 12 524 14 532
rect 22 524 24 532
rect 42 524 44 532
rect 52 524 54 532
rect 72 524 74 532
rect 82 524 84 532
rect 102 524 104 532
rect 112 524 114 532
rect 132 524 134 532
rect 142 524 144 532
rect 162 524 164 532
rect 172 524 174 532
rect 192 524 198 602
rect 0 516 198 524
rect 0 512 14 516
rect 0 4 4 512
rect 12 508 14 512
rect 22 508 24 516
rect 32 508 34 516
rect 42 508 44 516
rect 52 508 54 516
rect 62 508 64 516
rect 72 508 74 516
rect 82 508 84 516
rect 92 508 94 516
rect 102 508 104 516
rect 112 508 114 516
rect 122 508 124 516
rect 132 508 134 516
rect 142 508 144 516
rect 152 508 154 516
rect 162 508 164 516
rect 172 508 174 516
rect 182 508 184 516
rect 192 508 198 516
rect 12 504 198 508
rect 12 16 16 504
rect 28 486 54 492
rect 28 484 198 486
rect 28 466 36 484
rect 74 466 82 484
rect 28 462 82 466
rect 28 454 36 462
rect 54 456 82 462
rect 190 456 198 484
rect 54 454 198 456
rect 28 452 82 454
rect 28 444 36 452
rect 54 446 82 452
rect 190 446 198 454
rect 54 444 198 446
rect 28 442 198 444
rect 28 434 36 442
rect 54 434 198 442
rect 28 432 64 434
rect 28 424 36 432
rect 54 424 64 432
rect 28 422 64 424
rect 28 414 36 422
rect 54 414 64 422
rect 28 412 64 414
rect 28 404 36 412
rect 54 404 64 412
rect 28 402 64 404
rect 28 394 36 402
rect 54 394 64 402
rect 28 392 64 394
rect 28 384 36 392
rect 54 384 64 392
rect 28 382 64 384
rect 28 374 36 382
rect 54 374 64 382
rect 28 372 64 374
rect 28 364 36 372
rect 54 364 64 372
rect 28 362 64 364
rect 28 354 36 362
rect 54 354 64 362
rect 28 352 64 354
rect 28 344 36 352
rect 54 344 64 352
rect 28 342 64 344
rect 28 334 36 342
rect 54 334 64 342
rect 28 332 64 334
rect 28 324 36 332
rect 54 324 64 332
rect 28 322 64 324
rect 28 314 36 322
rect 54 314 64 322
rect 28 312 64 314
rect 28 304 36 312
rect 54 304 64 312
rect 28 302 64 304
rect 28 294 36 302
rect 54 294 64 302
rect 28 292 64 294
rect 28 284 36 292
rect 54 284 64 292
rect 28 282 64 284
rect 28 274 36 282
rect 54 274 64 282
rect 28 272 64 274
rect 28 264 36 272
rect 54 264 64 272
rect 28 262 64 264
rect 28 254 36 262
rect 54 254 64 262
rect 28 252 64 254
rect 28 244 36 252
rect 54 244 64 252
rect 28 242 64 244
rect 28 234 36 242
rect 54 234 64 242
rect 28 232 64 234
rect 28 224 36 232
rect 54 224 64 232
rect 28 222 64 224
rect 28 214 36 222
rect 54 214 64 222
rect 28 212 64 214
rect 28 204 36 212
rect 54 204 64 212
rect 28 202 64 204
rect 28 194 36 202
rect 54 194 64 202
rect 28 192 64 194
rect 28 184 36 192
rect 54 184 64 192
rect 28 182 64 184
rect 28 174 36 182
rect 54 174 64 182
rect 28 172 64 174
rect 28 164 36 172
rect 54 164 64 172
rect 28 162 64 164
rect 28 154 36 162
rect 54 154 64 162
rect 28 152 64 154
rect 28 144 36 152
rect 54 144 64 152
rect 28 142 64 144
rect 28 134 36 142
rect 54 134 64 142
rect 28 132 64 134
rect 28 124 36 132
rect 54 124 64 132
rect 28 122 64 124
rect 28 114 36 122
rect 54 114 64 122
rect 28 112 64 114
rect 28 104 36 112
rect 54 104 64 112
rect 28 102 64 104
rect 28 94 36 102
rect 54 94 64 102
rect 28 92 64 94
rect 28 84 36 92
rect 54 86 64 92
rect 72 430 198 434
rect 72 392 78 430
rect 196 422 198 430
rect 204 432 280 909
rect 294 885 306 895
rect 286 883 314 885
rect 286 844 314 846
rect 286 836 290 844
rect 298 836 302 844
rect 310 836 314 844
rect 286 834 314 836
rect 286 824 314 826
rect 286 816 290 824
rect 298 816 302 824
rect 310 816 314 824
rect 286 814 314 816
rect 286 804 314 806
rect 286 796 290 804
rect 298 796 302 804
rect 310 796 314 804
rect 286 794 314 796
rect 286 778 290 786
rect 298 778 302 786
rect 310 778 314 786
rect 286 776 314 778
rect 286 756 314 758
rect 286 748 290 756
rect 298 748 302 756
rect 310 748 314 756
rect 286 746 314 748
rect 286 736 314 738
rect 286 728 290 736
rect 298 728 302 736
rect 310 728 314 736
rect 286 726 314 728
rect 286 716 314 718
rect 286 708 290 716
rect 298 708 302 716
rect 310 708 314 716
rect 286 706 314 708
rect 286 696 314 698
rect 286 688 290 696
rect 298 688 302 696
rect 310 688 314 696
rect 286 652 314 654
rect 286 642 314 644
rect 286 632 314 634
rect 286 622 314 624
rect 286 612 314 614
rect 286 602 314 604
rect 286 592 314 594
rect 286 574 314 584
rect 286 564 314 566
rect 286 554 314 556
rect 286 544 314 546
rect 286 534 314 536
rect 286 524 314 526
rect 286 514 314 516
rect 286 504 314 506
rect 286 486 314 492
rect 286 456 314 458
rect 320 432 396 909
rect 402 914 404 922
rect 522 914 528 992
rect 536 1250 541 1252
rect 549 1250 550 1258
rect 558 1250 560 1258
rect 536 1248 560 1250
rect 536 1247 551 1248
rect 536 1239 542 1247
rect 550 1240 551 1247
rect 559 1240 560 1248
rect 550 1239 560 1240
rect 536 1238 560 1239
rect 536 1230 541 1238
rect 549 1230 550 1238
rect 558 1230 560 1238
rect 536 1228 560 1230
rect 536 1227 551 1228
rect 536 1219 542 1227
rect 550 1220 551 1227
rect 559 1220 560 1228
rect 550 1219 560 1220
rect 536 1218 560 1219
rect 536 1210 541 1218
rect 549 1210 550 1218
rect 558 1210 560 1218
rect 536 1208 560 1210
rect 536 1207 551 1208
rect 536 1199 542 1207
rect 550 1200 551 1207
rect 559 1200 560 1208
rect 550 1199 560 1200
rect 536 1198 560 1199
rect 536 1190 541 1198
rect 549 1190 550 1198
rect 558 1190 560 1198
rect 536 1188 560 1190
rect 536 1187 551 1188
rect 536 1179 542 1187
rect 550 1180 551 1187
rect 559 1180 560 1188
rect 550 1179 560 1180
rect 536 1178 560 1179
rect 536 1170 541 1178
rect 549 1170 550 1178
rect 558 1170 560 1178
rect 536 1168 560 1170
rect 536 1167 551 1168
rect 536 1159 542 1167
rect 550 1160 551 1167
rect 559 1160 560 1168
rect 550 1159 560 1160
rect 536 1158 560 1159
rect 536 1150 541 1158
rect 549 1150 550 1158
rect 558 1150 560 1158
rect 536 1148 560 1150
rect 536 1147 551 1148
rect 536 1139 542 1147
rect 550 1140 551 1147
rect 559 1140 560 1148
rect 550 1139 560 1140
rect 536 1138 560 1139
rect 536 1130 541 1138
rect 549 1130 550 1138
rect 558 1130 560 1138
rect 536 1128 560 1130
rect 536 1127 551 1128
rect 536 1119 542 1127
rect 550 1120 551 1127
rect 559 1120 560 1128
rect 550 1119 560 1120
rect 536 1118 560 1119
rect 536 1110 541 1118
rect 549 1110 550 1118
rect 558 1110 560 1118
rect 536 1108 560 1110
rect 536 1107 551 1108
rect 536 1099 542 1107
rect 550 1100 551 1107
rect 559 1100 560 1108
rect 550 1099 560 1100
rect 536 1098 560 1099
rect 536 1090 541 1098
rect 549 1090 550 1098
rect 558 1090 560 1098
rect 536 1088 560 1090
rect 536 1087 551 1088
rect 536 1079 542 1087
rect 550 1080 551 1087
rect 559 1080 560 1088
rect 550 1079 560 1080
rect 536 1078 560 1079
rect 536 1070 541 1078
rect 549 1070 550 1078
rect 558 1070 560 1078
rect 536 1068 560 1070
rect 536 1067 551 1068
rect 536 1059 542 1067
rect 550 1060 551 1067
rect 559 1060 560 1068
rect 550 1059 560 1060
rect 536 1058 560 1059
rect 536 1050 541 1058
rect 549 1050 550 1058
rect 558 1050 560 1058
rect 536 1048 560 1050
rect 536 1047 551 1048
rect 536 1039 542 1047
rect 550 1040 551 1047
rect 559 1040 560 1048
rect 550 1039 560 1040
rect 536 1038 560 1039
rect 536 1030 541 1038
rect 549 1030 550 1038
rect 558 1030 560 1038
rect 536 1028 560 1030
rect 536 1027 551 1028
rect 536 1019 542 1027
rect 550 1020 551 1027
rect 559 1020 560 1028
rect 550 1019 560 1020
rect 536 1018 560 1019
rect 536 1010 541 1018
rect 549 1010 550 1018
rect 558 1010 560 1018
rect 536 1008 560 1010
rect 536 1007 551 1008
rect 536 999 542 1007
rect 550 1000 551 1007
rect 559 1000 560 1008
rect 550 999 560 1000
rect 536 998 560 999
rect 536 990 541 998
rect 549 990 550 998
rect 558 990 560 998
rect 536 988 560 990
rect 536 987 551 988
rect 536 979 542 987
rect 550 980 551 987
rect 559 980 560 988
rect 550 979 560 980
rect 536 978 560 979
rect 536 970 541 978
rect 549 970 550 978
rect 558 970 560 978
rect 536 968 560 970
rect 536 967 551 968
rect 536 959 542 967
rect 550 960 551 967
rect 559 960 560 968
rect 550 959 560 960
rect 536 958 560 959
rect 536 950 541 958
rect 549 950 550 958
rect 558 950 560 958
rect 536 948 560 950
rect 536 947 551 948
rect 536 939 542 947
rect 550 940 551 947
rect 559 940 560 948
rect 550 939 560 940
rect 536 938 560 939
rect 536 930 541 938
rect 549 930 550 938
rect 558 930 560 938
rect 536 928 560 930
rect 536 927 551 928
rect 536 919 542 927
rect 550 920 551 927
rect 559 920 560 928
rect 550 919 560 920
rect 536 918 560 919
rect 536 914 541 918
rect 402 910 541 914
rect 549 910 550 918
rect 558 910 560 918
rect 402 908 560 910
rect 402 907 551 908
rect 402 899 542 907
rect 550 900 551 907
rect 559 900 560 908
rect 550 899 560 900
rect 402 898 560 899
rect 402 890 410 898
rect 518 890 541 898
rect 549 890 550 898
rect 558 890 560 898
rect 402 888 560 890
rect 402 883 542 888
rect 402 865 410 883
rect 538 880 542 883
rect 550 880 551 888
rect 559 880 560 888
rect 538 873 560 880
rect 558 865 560 873
rect 578 846 580 1318
rect 402 844 580 846
rect 402 738 408 844
rect 426 828 428 844
rect 436 828 438 844
rect 456 828 458 844
rect 466 828 468 844
rect 486 828 488 844
rect 496 828 498 844
rect 516 828 518 844
rect 526 828 528 844
rect 546 828 548 844
rect 556 828 558 844
rect 576 840 580 844
rect 598 840 600 1338
rect 576 836 600 840
rect 576 828 578 836
rect 586 828 588 836
rect 596 828 600 836
rect 416 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 416 818 418 826
rect 426 818 428 826
rect 446 818 448 826
rect 456 818 458 826
rect 476 818 478 826
rect 486 818 488 826
rect 506 818 508 826
rect 516 818 518 826
rect 536 818 538 826
rect 546 818 548 826
rect 566 818 568 826
rect 576 818 578 826
rect 586 818 588 826
rect 596 818 600 826
rect 416 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 426 808 428 816
rect 436 808 438 816
rect 456 808 458 816
rect 466 808 468 816
rect 486 808 488 816
rect 496 808 498 816
rect 516 808 518 816
rect 526 808 528 816
rect 546 808 548 816
rect 556 808 558 816
rect 576 808 578 816
rect 586 808 588 816
rect 596 808 600 816
rect 416 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 416 798 418 806
rect 426 798 428 806
rect 446 798 448 806
rect 456 798 458 806
rect 476 798 478 806
rect 486 798 488 806
rect 506 798 508 806
rect 516 798 518 806
rect 536 798 538 806
rect 546 798 548 806
rect 566 798 568 806
rect 576 798 578 806
rect 586 798 588 806
rect 596 798 600 806
rect 416 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 426 788 428 796
rect 436 788 438 796
rect 456 788 458 796
rect 466 788 468 796
rect 486 788 488 796
rect 496 788 498 796
rect 516 788 518 796
rect 526 788 528 796
rect 546 788 548 796
rect 556 788 558 796
rect 576 788 578 796
rect 586 788 588 796
rect 596 788 600 796
rect 416 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 416 778 418 786
rect 426 778 428 786
rect 416 776 428 778
rect 446 778 448 786
rect 456 778 458 786
rect 446 776 458 778
rect 476 778 478 786
rect 486 778 488 786
rect 476 776 488 778
rect 506 778 508 786
rect 516 778 518 786
rect 536 778 538 786
rect 546 778 548 786
rect 566 778 568 786
rect 576 778 578 786
rect 586 778 588 786
rect 596 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 516 768 518 776
rect 526 768 528 776
rect 546 768 548 776
rect 556 768 558 776
rect 576 768 578 776
rect 586 768 588 776
rect 596 768 600 776
rect 416 766 428 768
rect 416 758 418 766
rect 426 758 428 766
rect 446 766 458 768
rect 446 758 448 766
rect 456 758 458 766
rect 476 766 488 768
rect 476 758 478 766
rect 486 758 488 766
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 508 766
rect 516 758 518 766
rect 536 758 538 766
rect 546 758 548 766
rect 566 758 568 766
rect 576 758 578 766
rect 586 758 588 766
rect 596 758 600 766
rect 416 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 426 748 428 756
rect 436 748 438 756
rect 456 748 458 756
rect 466 748 468 756
rect 486 748 488 756
rect 496 748 498 756
rect 516 748 518 756
rect 526 748 528 756
rect 546 748 548 756
rect 556 748 558 756
rect 576 748 578 756
rect 586 748 588 756
rect 596 748 600 756
rect 416 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 416 738 418 746
rect 426 738 428 746
rect 446 738 448 746
rect 456 738 458 746
rect 476 738 478 746
rect 486 738 488 746
rect 506 738 508 746
rect 516 738 518 746
rect 536 738 538 746
rect 546 738 548 746
rect 566 738 568 746
rect 576 738 578 746
rect 586 738 588 746
rect 596 738 600 746
rect 560 736 600 738
rect 560 728 568 736
rect 576 728 578 736
rect 586 728 588 736
rect 596 728 600 736
rect 402 726 600 728
rect 402 688 408 726
rect 416 718 418 726
rect 426 718 428 726
rect 446 718 448 726
rect 456 718 458 726
rect 476 718 478 726
rect 486 718 488 726
rect 506 718 508 726
rect 516 718 518 726
rect 536 718 538 726
rect 546 718 548 726
rect 566 718 568 726
rect 576 718 578 726
rect 586 718 588 726
rect 596 718 600 726
rect 416 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 426 708 428 716
rect 436 708 438 716
rect 456 708 458 716
rect 466 708 468 716
rect 486 708 488 716
rect 496 708 498 716
rect 516 708 518 716
rect 526 708 528 716
rect 546 708 548 716
rect 556 708 558 716
rect 576 708 578 716
rect 586 708 588 716
rect 596 708 600 716
rect 416 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 416 698 418 706
rect 426 698 428 706
rect 446 698 448 706
rect 456 698 458 706
rect 476 698 478 706
rect 486 698 488 706
rect 506 698 508 706
rect 516 698 518 706
rect 536 698 538 706
rect 546 698 548 706
rect 566 698 568 706
rect 576 698 578 706
rect 586 698 588 706
rect 596 698 600 706
rect 416 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 426 688 428 696
rect 436 688 438 696
rect 456 688 458 696
rect 466 688 468 696
rect 486 688 488 696
rect 496 688 498 696
rect 516 688 518 696
rect 526 688 528 696
rect 546 688 548 696
rect 556 688 558 696
rect 576 688 578 696
rect 586 688 588 696
rect 596 688 600 696
rect 402 614 408 652
rect 426 644 428 652
rect 436 644 438 652
rect 456 644 458 652
rect 466 644 468 652
rect 486 644 488 652
rect 496 644 498 652
rect 516 644 518 652
rect 526 644 528 652
rect 546 644 548 652
rect 556 644 558 652
rect 576 644 578 652
rect 586 644 588 652
rect 596 644 600 652
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 416 634 418 642
rect 426 634 428 642
rect 446 634 448 642
rect 456 634 458 642
rect 476 634 478 642
rect 486 634 488 642
rect 506 634 508 642
rect 516 634 518 642
rect 536 634 538 642
rect 546 634 548 642
rect 566 634 568 642
rect 576 634 578 642
rect 586 634 588 642
rect 596 634 600 642
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 426 624 428 632
rect 436 624 438 632
rect 456 624 458 632
rect 466 624 468 632
rect 486 624 488 632
rect 496 624 498 632
rect 516 624 518 632
rect 526 624 528 632
rect 546 624 548 632
rect 556 624 558 632
rect 576 624 578 632
rect 586 624 588 632
rect 596 624 600 632
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 416 614 418 622
rect 426 614 428 622
rect 446 614 448 622
rect 456 614 458 622
rect 476 614 478 622
rect 486 614 488 622
rect 506 614 508 622
rect 516 614 518 622
rect 536 614 538 622
rect 546 614 548 622
rect 566 614 568 622
rect 576 614 578 622
rect 586 614 588 622
rect 596 614 600 622
rect 402 612 600 614
rect 560 604 568 612
rect 576 604 578 612
rect 586 604 588 612
rect 596 604 600 612
rect 560 602 600 604
rect 402 524 408 602
rect 416 594 418 602
rect 426 594 428 602
rect 446 594 448 602
rect 456 594 458 602
rect 476 594 478 602
rect 486 594 488 602
rect 506 594 508 602
rect 516 594 518 602
rect 536 594 538 602
rect 546 594 548 602
rect 566 594 568 602
rect 576 594 578 602
rect 586 594 588 602
rect 596 594 600 602
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 426 584 428 592
rect 436 584 438 592
rect 426 582 438 584
rect 456 584 458 592
rect 466 584 468 592
rect 456 582 468 584
rect 486 584 488 592
rect 496 584 498 592
rect 516 584 518 592
rect 526 584 528 592
rect 546 584 548 592
rect 556 584 558 592
rect 576 584 578 592
rect 586 584 588 592
rect 596 584 600 592
rect 486 582 498 584
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 506 574 508 582
rect 516 574 518 582
rect 536 574 538 582
rect 546 574 548 582
rect 566 574 568 582
rect 576 574 578 582
rect 586 574 588 582
rect 596 574 600 582
rect 426 572 438 574
rect 426 564 428 572
rect 436 564 438 572
rect 456 572 468 574
rect 456 564 458 572
rect 466 564 468 572
rect 486 572 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 486 564 488 572
rect 496 564 498 572
rect 516 564 518 572
rect 526 564 528 572
rect 546 564 548 572
rect 556 564 558 572
rect 576 564 578 572
rect 586 564 588 572
rect 596 564 600 572
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 416 554 418 562
rect 426 554 428 562
rect 446 554 448 562
rect 456 554 458 562
rect 476 554 478 562
rect 486 554 488 562
rect 506 554 508 562
rect 516 554 518 562
rect 536 554 538 562
rect 546 554 548 562
rect 566 554 568 562
rect 576 554 578 562
rect 586 554 588 562
rect 596 554 600 562
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 426 544 428 552
rect 436 544 438 552
rect 456 544 458 552
rect 466 544 468 552
rect 486 544 488 552
rect 496 544 498 552
rect 516 544 518 552
rect 526 544 528 552
rect 546 544 548 552
rect 556 544 558 552
rect 576 544 578 552
rect 586 544 588 552
rect 596 544 600 552
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 416 534 418 542
rect 426 534 428 542
rect 446 534 448 542
rect 456 534 458 542
rect 476 534 478 542
rect 486 534 488 542
rect 506 534 508 542
rect 516 534 518 542
rect 536 534 538 542
rect 546 534 548 542
rect 566 534 568 542
rect 576 534 578 542
rect 586 534 588 542
rect 596 534 600 542
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 426 524 428 532
rect 436 524 438 532
rect 456 524 458 532
rect 466 524 468 532
rect 486 524 488 532
rect 496 524 498 532
rect 516 524 518 532
rect 526 524 528 532
rect 546 524 548 532
rect 556 524 558 532
rect 576 524 578 532
rect 586 524 588 532
rect 596 524 600 532
rect 402 516 600 524
rect 402 508 408 516
rect 416 508 418 516
rect 426 508 428 516
rect 436 508 438 516
rect 446 508 448 516
rect 456 508 458 516
rect 466 508 468 516
rect 476 508 478 516
rect 486 508 488 516
rect 496 508 498 516
rect 506 508 508 516
rect 516 508 518 516
rect 526 508 528 516
rect 536 508 538 516
rect 546 508 548 516
rect 556 508 558 516
rect 566 508 568 516
rect 576 508 578 516
rect 586 512 600 516
rect 586 508 588 512
rect 402 504 588 508
rect 546 486 572 492
rect 204 416 396 432
rect 402 474 572 486
rect 402 456 416 474
rect 564 466 572 474
rect 504 462 572 466
rect 504 456 546 462
rect 402 454 546 456
rect 564 454 572 462
rect 402 446 410 454
rect 518 452 572 454
rect 518 446 546 452
rect 402 444 546 446
rect 564 444 572 452
rect 402 442 572 444
rect 402 434 546 442
rect 564 434 572 442
rect 402 430 528 434
rect 402 422 404 430
rect 72 388 106 392
rect 72 350 78 388
rect 112 406 488 416
rect 112 400 285 406
rect 315 400 488 406
rect 240 392 285 400
rect 112 388 285 392
rect 240 380 285 388
rect 112 370 285 380
rect 315 392 360 400
rect 315 388 488 392
rect 315 380 360 388
rect 315 370 488 380
rect 112 364 488 370
rect 522 392 528 430
rect 494 388 528 392
rect 236 350 240 358
rect 72 334 240 350
rect 72 326 82 334
rect 72 322 240 326
rect 72 314 82 322
rect 72 298 240 314
rect 72 220 78 298
rect 236 290 240 298
rect 246 284 354 364
rect 360 350 364 358
rect 522 350 528 388
rect 360 334 528 350
rect 518 326 528 334
rect 360 322 528 326
rect 518 314 528 322
rect 360 298 528 314
rect 360 290 364 298
rect 112 278 488 284
rect 112 268 285 278
rect 240 250 285 268
rect 112 242 285 250
rect 315 268 488 278
rect 315 250 360 268
rect 315 242 488 250
rect 112 234 488 242
rect 236 220 240 228
rect 72 204 240 220
rect 72 196 82 204
rect 72 192 240 196
rect 72 184 82 192
rect 72 168 240 184
rect 72 90 78 168
rect 236 160 240 168
rect 246 154 354 234
rect 360 220 364 228
rect 522 220 528 298
rect 360 204 528 220
rect 518 196 528 204
rect 360 192 528 196
rect 518 184 528 192
rect 360 168 528 184
rect 360 160 364 168
rect 112 150 488 154
rect 112 138 285 150
rect 240 120 285 138
rect 112 104 285 120
rect 196 90 198 98
rect 72 86 198 90
rect 54 84 198 86
rect 28 82 198 84
rect 28 74 36 82
rect 54 74 198 82
rect 28 72 82 74
rect 28 64 36 72
rect 54 66 82 72
rect 190 66 198 74
rect 54 64 198 66
rect 28 62 198 64
rect 28 54 36 62
rect 54 54 88 62
rect 28 52 88 54
rect 28 44 36 52
rect 84 44 88 52
rect 28 42 88 44
rect 28 34 36 42
rect 84 34 88 42
rect 96 34 98 62
rect 106 34 108 62
rect 116 34 118 62
rect 126 34 128 62
rect 136 34 138 62
rect 146 34 148 62
rect 156 34 158 62
rect 166 34 168 62
rect 176 34 178 62
rect 186 34 188 62
rect 196 34 198 62
rect 28 28 198 34
rect 204 82 285 104
rect 315 138 488 150
rect 315 120 360 138
rect 315 104 488 120
rect 315 82 396 104
rect 204 58 396 82
rect 204 30 206 58
rect 394 30 396 58
rect 204 24 396 30
rect 402 90 404 98
rect 522 90 528 168
rect 402 86 528 90
rect 536 432 572 434
rect 536 424 546 432
rect 564 424 572 432
rect 536 422 572 424
rect 536 414 546 422
rect 564 414 572 422
rect 536 412 572 414
rect 536 404 546 412
rect 564 404 572 412
rect 536 402 572 404
rect 536 394 546 402
rect 564 394 572 402
rect 536 392 572 394
rect 536 384 546 392
rect 564 384 572 392
rect 536 382 572 384
rect 536 374 546 382
rect 564 374 572 382
rect 536 372 572 374
rect 536 364 546 372
rect 564 364 572 372
rect 536 362 572 364
rect 536 354 546 362
rect 564 354 572 362
rect 536 352 572 354
rect 536 344 546 352
rect 564 344 572 352
rect 536 342 572 344
rect 536 334 546 342
rect 564 334 572 342
rect 536 332 572 334
rect 536 324 546 332
rect 564 324 572 332
rect 536 322 572 324
rect 536 314 546 322
rect 564 314 572 322
rect 536 312 572 314
rect 536 304 546 312
rect 564 304 572 312
rect 536 302 572 304
rect 536 294 546 302
rect 564 294 572 302
rect 536 292 572 294
rect 536 284 546 292
rect 564 284 572 292
rect 536 282 572 284
rect 536 274 546 282
rect 564 274 572 282
rect 536 272 572 274
rect 536 264 546 272
rect 564 264 572 272
rect 536 262 572 264
rect 536 254 546 262
rect 564 254 572 262
rect 536 252 572 254
rect 536 244 546 252
rect 564 244 572 252
rect 536 242 572 244
rect 536 234 546 242
rect 564 234 572 242
rect 536 232 572 234
rect 536 224 546 232
rect 564 224 572 232
rect 536 222 572 224
rect 536 214 546 222
rect 564 214 572 222
rect 536 212 572 214
rect 536 204 546 212
rect 564 204 572 212
rect 536 202 572 204
rect 536 194 546 202
rect 564 194 572 202
rect 536 192 572 194
rect 536 184 546 192
rect 564 184 572 192
rect 536 182 572 184
rect 536 174 546 182
rect 564 174 572 182
rect 536 172 572 174
rect 536 164 546 172
rect 564 164 572 172
rect 536 162 572 164
rect 536 154 546 162
rect 564 154 572 162
rect 536 152 572 154
rect 536 144 546 152
rect 564 144 572 152
rect 536 142 572 144
rect 536 134 546 142
rect 564 134 572 142
rect 536 132 572 134
rect 536 124 546 132
rect 564 124 572 132
rect 536 122 572 124
rect 536 114 546 122
rect 564 114 572 122
rect 536 112 572 114
rect 536 104 546 112
rect 564 104 572 112
rect 536 102 572 104
rect 536 94 546 102
rect 564 94 572 102
rect 536 92 572 94
rect 536 86 546 92
rect 402 84 546 86
rect 564 84 572 92
rect 402 82 572 84
rect 402 74 546 82
rect 564 74 572 82
rect 402 66 410 74
rect 518 72 572 74
rect 518 66 546 72
rect 402 64 546 66
rect 564 64 572 72
rect 402 62 572 64
rect 402 34 404 62
rect 412 34 414 62
rect 422 34 424 62
rect 432 34 434 62
rect 442 34 444 62
rect 452 34 454 62
rect 462 34 464 62
rect 472 34 474 62
rect 482 34 484 62
rect 492 34 494 62
rect 502 34 504 62
rect 512 54 546 62
rect 564 54 572 62
rect 512 52 572 54
rect 512 44 516 52
rect 564 44 572 52
rect 512 42 572 44
rect 512 34 516 42
rect 564 34 572 42
rect 402 28 572 34
rect 584 16 588 504
rect 12 14 198 16
rect 402 14 588 16
rect 12 12 588 14
rect 192 4 196 12
rect 404 4 408 12
rect 596 4 600 512
rect 0 2 600 4
rect 0 0 198 2
rect 402 0 600 2
<< m2contact >>
rect 42 1290 50 1298
rect 62 1290 70 1298
rect 50 1279 58 1287
rect 72 1284 80 1290
rect 92 1286 100 1294
rect 112 1286 120 1294
rect 132 1286 140 1294
rect 152 1286 160 1294
rect 172 1286 180 1294
rect 192 1286 200 1294
rect 212 1286 220 1294
rect 232 1286 240 1294
rect 72 1282 90 1284
rect 42 1270 50 1278
rect 82 1276 90 1282
rect 102 1276 110 1284
rect 122 1276 130 1284
rect 142 1276 150 1284
rect 162 1276 170 1284
rect 182 1276 190 1284
rect 202 1276 210 1284
rect 222 1276 230 1284
rect 50 1259 58 1267
rect 42 1250 50 1258
rect 50 1239 58 1247
rect 42 1230 50 1238
rect 50 1219 58 1227
rect 42 1210 50 1218
rect 50 1199 58 1207
rect 42 1190 50 1198
rect 50 1179 58 1187
rect 42 1170 50 1178
rect 50 1159 58 1167
rect 42 1150 50 1158
rect 50 1139 58 1147
rect 42 1130 50 1138
rect 50 1119 58 1127
rect 42 1110 50 1118
rect 50 1099 58 1107
rect 42 1090 50 1098
rect 50 1079 58 1087
rect 42 1070 50 1078
rect 50 1059 58 1067
rect 42 1050 50 1058
rect 50 1039 58 1047
rect 42 1030 50 1038
rect 50 1019 58 1027
rect 42 1010 50 1018
rect 50 999 58 1007
rect 42 990 50 998
rect 50 979 58 987
rect 42 970 50 978
rect 50 959 58 967
rect 42 950 50 958
rect 50 939 58 947
rect 42 930 50 938
rect 50 919 58 927
rect 42 910 50 918
rect 78 1242 236 1250
rect 78 1180 96 1242
rect 360 1286 368 1294
rect 380 1286 388 1294
rect 400 1286 408 1294
rect 420 1286 428 1294
rect 440 1286 448 1294
rect 460 1286 468 1294
rect 480 1286 488 1294
rect 500 1286 508 1294
rect 530 1290 538 1298
rect 550 1290 558 1298
rect 520 1284 528 1290
rect 370 1276 378 1284
rect 390 1276 398 1284
rect 410 1276 418 1284
rect 430 1276 438 1284
rect 450 1276 458 1284
rect 470 1276 478 1284
rect 490 1276 498 1284
rect 510 1282 528 1284
rect 510 1276 518 1282
rect 542 1279 550 1287
rect 550 1270 558 1278
rect 542 1259 550 1267
rect 364 1242 522 1250
rect 291 1210 309 1218
rect 78 1172 236 1180
rect 78 1114 236 1122
rect 78 1052 96 1114
rect 504 1180 522 1242
rect 364 1172 522 1180
rect 364 1114 522 1122
rect 291 1082 309 1090
rect 78 1044 236 1052
rect 78 984 236 992
rect 78 922 96 984
rect 504 1052 522 1114
rect 364 1044 522 1052
rect 364 984 522 992
rect 78 914 196 922
rect 50 899 58 907
rect 42 890 50 898
rect 50 880 58 888
rect 504 922 522 984
rect 24 836 42 844
rect 14 828 22 836
rect 44 828 52 836
rect 54 836 72 844
rect 74 828 82 836
rect 84 836 102 844
rect 104 828 112 836
rect 114 836 132 844
rect 134 828 142 836
rect 144 836 162 844
rect 164 828 172 836
rect 174 836 192 844
rect 4 818 12 826
rect 24 818 32 826
rect 54 818 62 826
rect 84 818 92 826
rect 114 818 122 826
rect 144 818 152 826
rect 174 818 182 826
rect 14 808 22 816
rect 44 808 52 816
rect 74 808 82 816
rect 104 808 112 816
rect 134 808 142 816
rect 164 808 172 816
rect 4 798 12 806
rect 24 798 32 806
rect 54 798 62 806
rect 84 798 92 806
rect 114 798 122 806
rect 144 798 152 806
rect 174 798 182 806
rect 14 788 22 796
rect 44 788 52 796
rect 74 788 82 796
rect 104 788 112 796
rect 134 788 142 796
rect 164 788 172 796
rect 4 778 12 786
rect 24 778 32 786
rect 54 778 62 786
rect 84 778 92 786
rect 114 778 122 786
rect 144 778 152 786
rect 174 778 182 786
rect 14 768 22 776
rect 44 768 52 776
rect 74 768 82 776
rect 4 758 12 766
rect 24 758 32 766
rect 54 758 62 766
rect 84 758 92 766
rect 114 758 122 766
rect 144 758 152 766
rect 174 758 182 766
rect 14 748 22 756
rect 44 748 52 756
rect 74 748 82 756
rect 104 748 112 756
rect 134 748 142 756
rect 164 748 172 756
rect 4 738 12 746
rect 24 738 32 746
rect 54 738 62 746
rect 84 738 92 746
rect 114 738 122 746
rect 144 738 152 746
rect 174 738 182 746
rect 14 728 22 736
rect 4 718 12 726
rect 24 718 32 726
rect 54 718 62 726
rect 84 718 92 726
rect 114 718 122 726
rect 144 718 152 726
rect 174 718 182 726
rect 14 708 22 716
rect 44 708 52 716
rect 74 708 82 716
rect 104 708 112 716
rect 134 708 142 716
rect 164 708 172 716
rect 4 698 12 706
rect 24 698 32 706
rect 54 698 62 706
rect 84 698 92 706
rect 114 698 122 706
rect 144 698 152 706
rect 174 698 182 706
rect 14 688 22 696
rect 44 688 52 696
rect 74 688 82 696
rect 104 688 112 696
rect 134 688 142 696
rect 164 688 172 696
rect 14 644 22 652
rect 44 644 52 652
rect 74 644 82 652
rect 104 644 112 652
rect 134 644 142 652
rect 164 644 172 652
rect 4 634 12 642
rect 24 634 32 642
rect 54 634 62 642
rect 84 634 92 642
rect 114 634 122 642
rect 144 634 152 642
rect 174 634 182 642
rect 14 624 22 632
rect 44 624 52 632
rect 74 624 82 632
rect 104 624 112 632
rect 134 624 142 632
rect 164 624 172 632
rect 4 614 12 622
rect 24 614 32 622
rect 54 614 62 622
rect 84 614 92 622
rect 114 614 122 622
rect 144 614 152 622
rect 174 614 182 622
rect 14 604 22 612
rect 4 594 12 602
rect 24 594 32 602
rect 54 594 62 602
rect 84 594 92 602
rect 114 594 122 602
rect 144 594 152 602
rect 174 594 182 602
rect 14 584 22 592
rect 44 584 52 592
rect 74 584 82 592
rect 104 584 112 592
rect 134 584 142 592
rect 164 584 172 592
rect 4 574 12 582
rect 24 574 32 582
rect 54 574 62 582
rect 84 574 92 582
rect 14 564 22 572
rect 44 564 52 572
rect 74 564 82 572
rect 104 564 112 572
rect 134 564 142 572
rect 164 564 172 572
rect 4 554 12 562
rect 24 554 32 562
rect 54 554 62 562
rect 84 554 92 562
rect 114 554 122 562
rect 144 554 152 562
rect 174 554 182 562
rect 14 544 22 552
rect 44 544 52 552
rect 74 544 82 552
rect 104 544 112 552
rect 134 544 142 552
rect 164 544 172 552
rect 4 534 12 542
rect 24 534 32 542
rect 54 534 62 542
rect 84 534 92 542
rect 114 534 122 542
rect 144 534 152 542
rect 174 534 182 542
rect 14 524 22 532
rect 44 524 52 532
rect 74 524 82 532
rect 104 524 112 532
rect 134 524 142 532
rect 164 524 172 532
rect 14 508 22 516
rect 34 508 42 516
rect 54 508 62 516
rect 74 508 82 516
rect 94 508 102 516
rect 114 508 122 516
rect 134 508 142 516
rect 154 508 162 516
rect 174 508 182 516
rect 36 444 54 452
rect 36 424 54 432
rect 36 404 54 412
rect 36 384 54 392
rect 36 364 54 372
rect 36 344 54 352
rect 36 324 54 332
rect 36 304 54 312
rect 36 284 54 292
rect 36 264 54 272
rect 36 244 54 252
rect 36 224 54 232
rect 36 204 54 212
rect 36 184 54 192
rect 36 164 54 172
rect 36 144 54 152
rect 36 124 54 132
rect 36 104 54 112
rect 36 84 54 92
rect 78 422 196 430
rect 286 895 314 903
rect 286 885 294 895
rect 306 885 314 895
rect 290 836 298 844
rect 302 836 310 844
rect 290 816 298 824
rect 302 816 310 824
rect 290 796 298 804
rect 302 796 310 804
rect 290 778 298 786
rect 302 778 310 786
rect 290 748 298 756
rect 302 748 310 756
rect 290 728 298 736
rect 302 728 310 736
rect 290 708 298 716
rect 302 708 310 716
rect 290 688 298 696
rect 302 688 310 696
rect 286 644 314 652
rect 286 624 314 632
rect 286 604 314 612
rect 286 584 314 592
rect 286 556 314 564
rect 286 536 314 544
rect 286 516 314 524
rect 286 438 314 456
rect 404 914 522 922
rect 550 1250 558 1258
rect 542 1239 550 1247
rect 550 1230 558 1238
rect 542 1219 550 1227
rect 550 1210 558 1218
rect 542 1199 550 1207
rect 550 1190 558 1198
rect 542 1179 550 1187
rect 550 1170 558 1178
rect 542 1159 550 1167
rect 550 1150 558 1158
rect 542 1139 550 1147
rect 550 1130 558 1138
rect 542 1119 550 1127
rect 550 1110 558 1118
rect 542 1099 550 1107
rect 550 1090 558 1098
rect 542 1079 550 1087
rect 550 1070 558 1078
rect 542 1059 550 1067
rect 550 1050 558 1058
rect 542 1039 550 1047
rect 550 1030 558 1038
rect 542 1019 550 1027
rect 550 1010 558 1018
rect 542 999 550 1007
rect 550 990 558 998
rect 542 979 550 987
rect 550 970 558 978
rect 542 959 550 967
rect 550 950 558 958
rect 542 939 550 947
rect 550 930 558 938
rect 542 919 550 927
rect 550 910 558 918
rect 542 899 550 907
rect 550 890 558 898
rect 542 880 550 888
rect 408 836 426 844
rect 428 828 436 836
rect 438 836 456 844
rect 458 828 466 836
rect 468 836 486 844
rect 488 828 496 836
rect 498 836 516 844
rect 518 828 526 836
rect 528 836 546 844
rect 548 828 556 836
rect 558 836 576 844
rect 578 828 586 836
rect 418 818 426 826
rect 448 818 456 826
rect 478 818 486 826
rect 508 818 516 826
rect 538 818 546 826
rect 568 818 576 826
rect 588 818 596 826
rect 428 808 436 816
rect 458 808 466 816
rect 488 808 496 816
rect 518 808 526 816
rect 548 808 556 816
rect 578 808 586 816
rect 418 798 426 806
rect 448 798 456 806
rect 478 798 486 806
rect 508 798 516 806
rect 538 798 546 806
rect 568 798 576 806
rect 588 798 596 806
rect 428 788 436 796
rect 458 788 466 796
rect 488 788 496 796
rect 518 788 526 796
rect 548 788 556 796
rect 578 788 586 796
rect 418 778 426 786
rect 448 778 456 786
rect 478 778 486 786
rect 508 778 516 786
rect 538 778 546 786
rect 568 778 576 786
rect 588 778 596 786
rect 518 768 526 776
rect 548 768 556 776
rect 578 768 586 776
rect 418 758 426 766
rect 448 758 456 766
rect 478 758 486 766
rect 508 758 516 766
rect 538 758 546 766
rect 568 758 576 766
rect 588 758 596 766
rect 428 748 436 756
rect 458 748 466 756
rect 488 748 496 756
rect 518 748 526 756
rect 548 748 556 756
rect 578 748 586 756
rect 418 738 426 746
rect 448 738 456 746
rect 478 738 486 746
rect 508 738 516 746
rect 538 738 546 746
rect 568 738 576 746
rect 588 738 596 746
rect 578 728 586 736
rect 418 718 426 726
rect 448 718 456 726
rect 478 718 486 726
rect 508 718 516 726
rect 538 718 546 726
rect 568 718 576 726
rect 588 718 596 726
rect 428 708 436 716
rect 458 708 466 716
rect 488 708 496 716
rect 518 708 526 716
rect 548 708 556 716
rect 578 708 586 716
rect 418 698 426 706
rect 448 698 456 706
rect 478 698 486 706
rect 508 698 516 706
rect 538 698 546 706
rect 568 698 576 706
rect 588 698 596 706
rect 428 688 436 696
rect 458 688 466 696
rect 488 688 496 696
rect 518 688 526 696
rect 548 688 556 696
rect 578 688 586 696
rect 428 644 436 652
rect 458 644 466 652
rect 488 644 496 652
rect 518 644 526 652
rect 548 644 556 652
rect 578 644 586 652
rect 418 634 426 642
rect 448 634 456 642
rect 478 634 486 642
rect 508 634 516 642
rect 538 634 546 642
rect 568 634 576 642
rect 588 634 596 642
rect 428 624 436 632
rect 458 624 466 632
rect 488 624 496 632
rect 518 624 526 632
rect 548 624 556 632
rect 578 624 586 632
rect 418 614 426 622
rect 448 614 456 622
rect 478 614 486 622
rect 508 614 516 622
rect 538 614 546 622
rect 568 614 576 622
rect 588 614 596 622
rect 578 604 586 612
rect 418 594 426 602
rect 448 594 456 602
rect 478 594 486 602
rect 508 594 516 602
rect 538 594 546 602
rect 568 594 576 602
rect 588 594 596 602
rect 428 584 436 592
rect 458 584 466 592
rect 488 584 496 592
rect 518 584 526 592
rect 548 584 556 592
rect 578 584 586 592
rect 508 574 516 582
rect 538 574 546 582
rect 568 574 576 582
rect 588 574 596 582
rect 428 564 436 572
rect 458 564 466 572
rect 488 564 496 572
rect 518 564 526 572
rect 548 564 556 572
rect 578 564 586 572
rect 418 554 426 562
rect 448 554 456 562
rect 478 554 486 562
rect 508 554 516 562
rect 538 554 546 562
rect 568 554 576 562
rect 588 554 596 562
rect 428 544 436 552
rect 458 544 466 552
rect 488 544 496 552
rect 518 544 526 552
rect 548 544 556 552
rect 578 544 586 552
rect 418 534 426 542
rect 448 534 456 542
rect 478 534 486 542
rect 508 534 516 542
rect 538 534 546 542
rect 568 534 576 542
rect 588 534 596 542
rect 428 524 436 532
rect 458 524 466 532
rect 488 524 496 532
rect 518 524 526 532
rect 548 524 556 532
rect 578 524 586 532
rect 418 508 426 516
rect 438 508 446 516
rect 458 508 466 516
rect 478 508 486 516
rect 498 508 506 516
rect 518 508 526 516
rect 538 508 546 516
rect 558 508 566 516
rect 578 508 586 516
rect 78 392 106 422
rect 546 444 564 452
rect 404 422 522 430
rect 78 358 106 388
rect 291 384 309 392
rect 494 392 522 422
rect 78 350 236 358
rect 78 290 236 298
rect 78 228 106 290
rect 494 358 522 388
rect 364 350 522 358
rect 364 290 522 298
rect 291 256 309 264
rect 78 220 236 228
rect 78 160 236 168
rect 78 98 106 160
rect 494 228 522 290
rect 364 220 522 228
rect 364 160 522 168
rect 78 90 196 98
rect 36 64 54 72
rect 36 44 84 52
rect 98 34 106 62
rect 118 34 126 62
rect 138 34 146 62
rect 158 34 166 62
rect 178 34 186 62
rect 291 128 309 136
rect 291 112 309 120
rect 291 96 309 104
rect 494 98 522 160
rect 206 30 394 58
rect 404 90 522 98
rect 546 424 564 432
rect 546 404 564 412
rect 546 384 564 392
rect 546 364 564 372
rect 546 344 564 352
rect 546 324 564 332
rect 546 304 564 312
rect 546 284 564 292
rect 546 264 564 272
rect 546 244 564 252
rect 546 224 564 232
rect 546 204 564 212
rect 546 184 564 192
rect 546 164 564 172
rect 546 144 564 152
rect 546 124 564 132
rect 546 104 564 112
rect 546 84 564 92
rect 546 64 564 72
rect 414 34 422 62
rect 434 34 442 62
rect 454 34 462 62
rect 474 34 482 62
rect 494 34 502 62
rect 516 44 564 52
<< metal2 >>
rect 0 1298 600 1340
rect 0 1290 42 1298
rect 50 1290 62 1298
rect 70 1294 530 1298
rect 70 1290 92 1294
rect 0 1287 72 1290
rect 0 1279 50 1287
rect 58 1282 72 1287
rect 80 1286 92 1290
rect 100 1286 112 1294
rect 120 1286 132 1294
rect 140 1286 152 1294
rect 160 1286 172 1294
rect 180 1286 192 1294
rect 200 1286 212 1294
rect 220 1286 232 1294
rect 240 1286 360 1294
rect 368 1286 380 1294
rect 388 1286 400 1294
rect 408 1286 420 1294
rect 428 1286 440 1294
rect 448 1286 460 1294
rect 468 1286 480 1294
rect 488 1286 500 1294
rect 508 1290 530 1294
rect 538 1290 550 1298
rect 558 1290 600 1298
rect 508 1286 520 1290
rect 80 1284 520 1286
rect 528 1287 600 1290
rect 58 1279 82 1282
rect 0 1278 82 1279
rect 0 1270 42 1278
rect 50 1276 82 1278
rect 90 1276 102 1284
rect 110 1276 122 1284
rect 130 1276 142 1284
rect 150 1276 162 1284
rect 170 1276 182 1284
rect 190 1276 202 1284
rect 210 1276 222 1284
rect 230 1276 370 1284
rect 378 1276 390 1284
rect 398 1276 410 1284
rect 418 1276 430 1284
rect 438 1276 450 1284
rect 458 1276 470 1284
rect 478 1276 490 1284
rect 498 1276 510 1284
rect 528 1282 542 1287
rect 518 1279 542 1282
rect 550 1279 600 1287
rect 518 1278 600 1279
rect 518 1276 550 1278
rect 50 1270 550 1276
rect 558 1270 600 1278
rect 0 1267 600 1270
rect 0 1259 50 1267
rect 58 1259 542 1267
rect 550 1259 600 1267
rect 0 1258 600 1259
rect 0 1250 42 1258
rect 50 1250 550 1258
rect 558 1250 600 1258
rect 0 1247 78 1250
rect 0 1239 50 1247
rect 58 1239 78 1247
rect 236 1242 364 1250
rect 522 1247 600 1250
rect 0 1238 78 1239
rect 0 1230 42 1238
rect 50 1230 78 1238
rect 0 1227 78 1230
rect 0 1219 50 1227
rect 58 1219 78 1227
rect 0 1218 78 1219
rect 0 1210 42 1218
rect 50 1210 78 1218
rect 0 1207 78 1210
rect 0 1199 50 1207
rect 58 1199 78 1207
rect 0 1198 78 1199
rect 0 1190 42 1198
rect 50 1190 78 1198
rect 0 1187 78 1190
rect 0 1179 50 1187
rect 58 1179 78 1187
rect 96 1218 504 1242
rect 96 1210 291 1218
rect 309 1210 504 1218
rect 96 1190 504 1210
rect 96 1180 100 1190
rect 500 1180 504 1190
rect 522 1239 542 1247
rect 550 1239 600 1247
rect 522 1238 600 1239
rect 522 1230 550 1238
rect 558 1230 600 1238
rect 522 1227 600 1230
rect 522 1219 542 1227
rect 550 1219 600 1227
rect 522 1218 600 1219
rect 522 1210 550 1218
rect 558 1210 600 1218
rect 522 1207 600 1210
rect 522 1199 542 1207
rect 550 1199 600 1207
rect 522 1198 600 1199
rect 522 1190 550 1198
rect 558 1190 600 1198
rect 522 1187 600 1190
rect 0 1178 78 1179
rect 0 1170 42 1178
rect 50 1172 78 1178
rect 236 1172 364 1180
rect 522 1179 542 1187
rect 550 1179 600 1187
rect 522 1178 600 1179
rect 522 1172 550 1178
rect 50 1170 550 1172
rect 558 1170 600 1178
rect 0 1167 600 1170
rect 0 1159 50 1167
rect 58 1159 542 1167
rect 550 1159 600 1167
rect 0 1158 600 1159
rect 0 1150 42 1158
rect 50 1150 550 1158
rect 558 1150 600 1158
rect 0 1147 600 1150
rect 0 1139 50 1147
rect 58 1139 542 1147
rect 550 1139 600 1147
rect 0 1138 600 1139
rect 0 1130 42 1138
rect 50 1130 550 1138
rect 558 1130 600 1138
rect 0 1127 600 1130
rect 0 1119 50 1127
rect 58 1122 542 1127
rect 58 1119 78 1122
rect 0 1118 78 1119
rect 0 1110 42 1118
rect 50 1110 78 1118
rect 236 1114 364 1122
rect 522 1119 542 1122
rect 550 1119 600 1127
rect 522 1118 600 1119
rect 0 1107 78 1110
rect 0 1099 50 1107
rect 58 1099 78 1107
rect 0 1098 78 1099
rect 0 1090 42 1098
rect 50 1090 78 1098
rect 0 1087 78 1090
rect 0 1079 50 1087
rect 58 1079 78 1087
rect 0 1078 78 1079
rect 0 1070 42 1078
rect 50 1070 78 1078
rect 0 1067 78 1070
rect 0 1059 50 1067
rect 58 1059 78 1067
rect 0 1058 78 1059
rect 0 1050 42 1058
rect 50 1050 78 1058
rect 96 1090 504 1114
rect 96 1082 291 1090
rect 309 1082 504 1090
rect 96 1052 504 1082
rect 522 1110 550 1118
rect 558 1110 600 1118
rect 522 1107 600 1110
rect 522 1099 542 1107
rect 550 1099 600 1107
rect 522 1098 600 1099
rect 522 1090 550 1098
rect 558 1090 600 1098
rect 522 1087 600 1090
rect 522 1079 542 1087
rect 550 1079 600 1087
rect 522 1078 600 1079
rect 522 1070 550 1078
rect 558 1070 600 1078
rect 522 1067 600 1070
rect 522 1059 542 1067
rect 550 1059 600 1067
rect 522 1058 600 1059
rect 0 1047 78 1050
rect 0 1039 50 1047
rect 58 1044 78 1047
rect 236 1044 364 1052
rect 522 1050 550 1058
rect 558 1050 600 1058
rect 522 1047 600 1050
rect 522 1044 542 1047
rect 58 1040 542 1044
rect 58 1039 100 1040
rect 0 1038 100 1039
rect 0 1030 42 1038
rect 50 1030 100 1038
rect 500 1039 542 1040
rect 550 1039 600 1047
rect 500 1038 600 1039
rect 500 1030 550 1038
rect 558 1030 600 1038
rect 0 1027 600 1030
rect 0 1019 50 1027
rect 58 1019 542 1027
rect 550 1019 600 1027
rect 0 1018 600 1019
rect 0 1010 42 1018
rect 50 1010 550 1018
rect 558 1010 600 1018
rect 0 1007 600 1010
rect 0 999 50 1007
rect 58 999 542 1007
rect 550 999 600 1007
rect 0 998 600 999
rect 0 990 42 998
rect 50 992 550 998
rect 50 990 78 992
rect 0 987 78 990
rect 0 979 50 987
rect 58 979 78 987
rect 236 984 364 992
rect 522 990 550 992
rect 558 990 600 998
rect 522 987 600 990
rect 0 978 78 979
rect 0 970 42 978
rect 50 970 78 978
rect 0 967 78 970
rect 0 959 50 967
rect 58 959 78 967
rect 0 958 78 959
rect 0 950 42 958
rect 50 950 78 958
rect 0 947 78 950
rect 0 939 50 947
rect 58 939 78 947
rect 0 938 78 939
rect 0 930 42 938
rect 50 930 78 938
rect 0 927 78 930
rect 0 919 50 927
rect 58 919 78 927
rect 96 922 504 984
rect 522 979 542 987
rect 550 979 600 987
rect 522 978 600 979
rect 522 970 550 978
rect 558 970 600 978
rect 522 967 600 970
rect 522 959 542 967
rect 550 959 600 967
rect 522 958 600 959
rect 522 950 550 958
rect 558 950 600 958
rect 522 947 600 950
rect 522 939 542 947
rect 550 939 600 947
rect 522 938 600 939
rect 522 930 550 938
rect 558 930 600 938
rect 522 927 600 930
rect 0 918 78 919
rect 0 910 42 918
rect 50 914 78 918
rect 196 914 404 922
rect 522 919 542 927
rect 550 919 600 927
rect 522 918 600 919
rect 522 914 550 918
rect 50 910 550 914
rect 558 910 600 918
rect 0 907 600 910
rect 0 899 50 907
rect 58 903 542 907
rect 58 899 286 903
rect 0 898 286 899
rect 0 890 42 898
rect 50 890 286 898
rect 314 899 542 903
rect 550 899 600 907
rect 314 898 600 899
rect 0 888 286 890
rect 0 880 50 888
rect 58 885 286 888
rect 294 885 306 895
rect 314 890 550 898
rect 558 890 600 898
rect 314 888 600 890
rect 314 885 542 888
rect 58 880 542 885
rect 550 880 600 888
rect 0 844 600 848
rect 0 836 24 844
rect 42 836 54 844
rect 72 836 84 844
rect 102 836 114 844
rect 132 836 144 844
rect 162 836 174 844
rect 192 836 290 844
rect 298 836 302 844
rect 310 836 408 844
rect 426 836 438 844
rect 456 836 468 844
rect 486 836 498 844
rect 516 836 528 844
rect 546 836 558 844
rect 576 836 600 844
rect 0 828 14 836
rect 22 828 44 836
rect 52 828 74 836
rect 82 828 104 836
rect 112 828 134 836
rect 142 828 164 836
rect 172 828 428 836
rect 436 828 458 836
rect 466 828 488 836
rect 496 828 518 836
rect 526 828 548 836
rect 556 828 578 836
rect 586 828 600 836
rect 0 826 600 828
rect 0 818 4 826
rect 12 818 24 826
rect 32 818 54 826
rect 62 818 84 826
rect 92 818 114 826
rect 122 818 144 826
rect 152 818 174 826
rect 182 824 418 826
rect 182 818 290 824
rect 0 816 290 818
rect 298 816 302 824
rect 310 818 418 824
rect 426 818 448 826
rect 456 818 478 826
rect 486 818 508 826
rect 516 818 538 826
rect 546 818 568 826
rect 576 818 588 826
rect 596 818 600 826
rect 310 816 600 818
rect 0 808 14 816
rect 22 808 44 816
rect 52 808 74 816
rect 82 808 104 816
rect 112 808 134 816
rect 142 808 164 816
rect 172 808 428 816
rect 436 808 458 816
rect 466 808 488 816
rect 496 808 518 816
rect 526 808 548 816
rect 556 808 578 816
rect 586 808 600 816
rect 0 806 600 808
rect 0 798 4 806
rect 12 798 24 806
rect 32 798 54 806
rect 62 798 84 806
rect 92 798 114 806
rect 122 798 144 806
rect 152 798 174 806
rect 182 804 418 806
rect 182 798 290 804
rect 0 796 290 798
rect 298 796 302 804
rect 310 798 418 804
rect 426 798 448 806
rect 456 798 478 806
rect 486 798 508 806
rect 516 798 538 806
rect 546 798 568 806
rect 576 798 588 806
rect 596 798 600 806
rect 310 796 600 798
rect 0 788 14 796
rect 22 788 44 796
rect 52 788 74 796
rect 82 788 104 796
rect 112 788 134 796
rect 142 788 164 796
rect 172 788 428 796
rect 436 788 458 796
rect 466 788 488 796
rect 496 788 518 796
rect 526 788 548 796
rect 556 788 578 796
rect 586 788 600 796
rect 0 786 600 788
rect 0 778 4 786
rect 12 778 24 786
rect 32 778 54 786
rect 62 778 84 786
rect 92 778 114 786
rect 122 778 144 786
rect 152 778 174 786
rect 182 778 290 786
rect 298 778 302 786
rect 310 778 418 786
rect 426 778 448 786
rect 456 778 478 786
rect 486 778 508 786
rect 516 778 538 786
rect 546 778 568 786
rect 576 778 588 786
rect 596 778 600 786
rect 0 776 100 778
rect 0 768 14 776
rect 22 768 44 776
rect 52 768 74 776
rect 82 768 100 776
rect 500 776 600 778
rect 500 768 518 776
rect 526 768 548 776
rect 556 768 578 776
rect 586 768 600 776
rect 0 766 600 768
rect 0 758 4 766
rect 12 758 24 766
rect 32 758 54 766
rect 62 758 84 766
rect 92 758 114 766
rect 122 758 144 766
rect 152 758 174 766
rect 182 758 418 766
rect 426 758 448 766
rect 456 758 478 766
rect 486 758 508 766
rect 516 758 538 766
rect 546 758 568 766
rect 576 758 588 766
rect 596 758 600 766
rect 0 756 600 758
rect 0 748 14 756
rect 22 748 44 756
rect 52 748 74 756
rect 82 748 104 756
rect 112 748 134 756
rect 142 748 164 756
rect 172 748 290 756
rect 298 748 302 756
rect 310 748 428 756
rect 436 748 458 756
rect 466 748 488 756
rect 496 748 518 756
rect 526 748 548 756
rect 556 748 578 756
rect 586 748 600 756
rect 0 746 600 748
rect 0 738 4 746
rect 12 738 24 746
rect 32 738 54 746
rect 62 738 84 746
rect 92 738 114 746
rect 122 738 144 746
rect 152 738 174 746
rect 182 738 418 746
rect 426 738 448 746
rect 456 738 478 746
rect 486 738 508 746
rect 516 738 538 746
rect 546 738 568 746
rect 576 738 588 746
rect 596 738 600 746
rect 0 736 600 738
rect 0 728 14 736
rect 22 728 290 736
rect 298 728 302 736
rect 310 728 578 736
rect 586 728 600 736
rect 0 726 600 728
rect 0 718 4 726
rect 12 718 24 726
rect 32 718 54 726
rect 62 718 84 726
rect 92 718 114 726
rect 122 718 144 726
rect 152 718 174 726
rect 182 718 418 726
rect 426 718 448 726
rect 456 718 478 726
rect 486 718 508 726
rect 516 718 538 726
rect 546 718 568 726
rect 576 718 588 726
rect 596 718 600 726
rect 0 716 600 718
rect 0 708 14 716
rect 22 708 44 716
rect 52 708 74 716
rect 82 708 104 716
rect 112 708 134 716
rect 142 708 164 716
rect 172 708 290 716
rect 298 708 302 716
rect 310 708 428 716
rect 436 708 458 716
rect 466 708 488 716
rect 496 708 518 716
rect 526 708 548 716
rect 556 708 578 716
rect 586 708 600 716
rect 0 706 600 708
rect 0 698 4 706
rect 12 698 24 706
rect 32 698 54 706
rect 62 698 84 706
rect 92 698 114 706
rect 122 698 144 706
rect 152 698 174 706
rect 182 698 418 706
rect 426 698 448 706
rect 456 698 478 706
rect 486 698 508 706
rect 516 698 538 706
rect 546 698 568 706
rect 576 698 588 706
rect 596 698 600 706
rect 0 696 600 698
rect 0 688 14 696
rect 22 688 44 696
rect 52 688 74 696
rect 82 688 104 696
rect 112 688 134 696
rect 142 688 164 696
rect 172 688 290 696
rect 298 688 302 696
rect 310 688 428 696
rect 436 688 458 696
rect 466 688 488 696
rect 496 688 518 696
rect 526 688 548 696
rect 556 688 578 696
rect 586 688 600 696
rect 0 644 14 652
rect 22 644 44 652
rect 52 644 74 652
rect 82 644 104 652
rect 112 644 134 652
rect 142 644 164 652
rect 172 644 286 652
rect 314 644 428 652
rect 436 644 458 652
rect 466 644 488 652
rect 496 644 518 652
rect 526 644 548 652
rect 556 644 578 652
rect 586 644 600 652
rect 0 642 600 644
rect 0 634 4 642
rect 12 634 24 642
rect 32 634 54 642
rect 62 634 84 642
rect 92 634 114 642
rect 122 634 144 642
rect 152 634 174 642
rect 182 634 418 642
rect 426 634 448 642
rect 456 634 478 642
rect 486 634 508 642
rect 516 634 538 642
rect 546 634 568 642
rect 576 634 588 642
rect 596 634 600 642
rect 0 632 600 634
rect 0 624 14 632
rect 22 624 44 632
rect 52 624 74 632
rect 82 624 104 632
rect 112 624 134 632
rect 142 624 164 632
rect 172 624 286 632
rect 314 624 428 632
rect 436 624 458 632
rect 466 624 488 632
rect 496 624 518 632
rect 526 624 548 632
rect 556 624 578 632
rect 586 624 600 632
rect 0 622 600 624
rect 0 614 4 622
rect 12 614 24 622
rect 32 614 54 622
rect 62 614 84 622
rect 92 614 114 622
rect 122 614 144 622
rect 152 614 174 622
rect 182 614 418 622
rect 426 614 448 622
rect 456 614 478 622
rect 486 614 508 622
rect 516 614 538 622
rect 546 614 568 622
rect 576 614 588 622
rect 596 614 600 622
rect 0 612 600 614
rect 0 604 14 612
rect 22 604 286 612
rect 314 604 578 612
rect 586 604 600 612
rect 0 602 600 604
rect 0 594 4 602
rect 12 594 24 602
rect 32 594 54 602
rect 62 594 84 602
rect 92 594 114 602
rect 122 594 144 602
rect 152 594 174 602
rect 182 594 418 602
rect 426 594 448 602
rect 456 594 478 602
rect 486 594 508 602
rect 516 594 538 602
rect 546 594 568 602
rect 576 594 588 602
rect 596 594 600 602
rect 0 592 600 594
rect 0 584 14 592
rect 22 584 44 592
rect 52 584 74 592
rect 82 584 104 592
rect 112 584 134 592
rect 142 584 164 592
rect 172 584 286 592
rect 314 584 428 592
rect 436 584 458 592
rect 466 584 488 592
rect 496 584 518 592
rect 526 584 548 592
rect 556 584 578 592
rect 586 584 600 592
rect 0 582 600 584
rect 0 574 4 582
rect 12 574 24 582
rect 32 574 54 582
rect 62 574 84 582
rect 92 574 100 582
rect 0 572 100 574
rect 500 574 508 582
rect 516 574 538 582
rect 546 574 568 582
rect 576 574 588 582
rect 596 574 600 582
rect 500 572 600 574
rect 0 564 14 572
rect 22 564 44 572
rect 52 564 74 572
rect 82 564 104 572
rect 112 564 134 572
rect 142 564 164 572
rect 172 564 428 572
rect 436 564 458 572
rect 466 564 488 572
rect 496 564 518 572
rect 526 564 548 572
rect 556 564 578 572
rect 586 564 600 572
rect 0 562 286 564
rect 0 554 4 562
rect 12 554 24 562
rect 32 554 54 562
rect 62 554 84 562
rect 92 554 114 562
rect 122 554 144 562
rect 152 554 174 562
rect 182 556 286 562
rect 314 562 600 564
rect 314 556 418 562
rect 182 554 418 556
rect 426 554 448 562
rect 456 554 478 562
rect 486 554 508 562
rect 516 554 538 562
rect 546 554 568 562
rect 576 554 588 562
rect 596 554 600 562
rect 0 552 600 554
rect 0 544 14 552
rect 22 544 44 552
rect 52 544 74 552
rect 82 544 104 552
rect 112 544 134 552
rect 142 544 164 552
rect 172 544 428 552
rect 436 544 458 552
rect 466 544 488 552
rect 496 544 518 552
rect 526 544 548 552
rect 556 544 578 552
rect 586 544 600 552
rect 0 542 286 544
rect 0 534 4 542
rect 12 534 24 542
rect 32 534 54 542
rect 62 534 84 542
rect 92 534 114 542
rect 122 534 144 542
rect 152 534 174 542
rect 182 536 286 542
rect 314 542 600 544
rect 314 536 418 542
rect 182 534 418 536
rect 426 534 448 542
rect 456 534 478 542
rect 486 534 508 542
rect 516 534 538 542
rect 546 534 568 542
rect 576 534 588 542
rect 596 534 600 542
rect 0 532 600 534
rect 0 524 14 532
rect 22 524 44 532
rect 52 524 74 532
rect 82 524 104 532
rect 112 524 134 532
rect 142 524 164 532
rect 172 524 428 532
rect 436 524 458 532
rect 466 524 488 532
rect 496 524 518 532
rect 526 524 548 532
rect 556 524 578 532
rect 586 524 600 532
rect 0 516 286 524
rect 314 516 600 524
rect 0 508 14 516
rect 22 508 34 516
rect 42 508 54 516
rect 62 508 74 516
rect 82 508 94 516
rect 102 508 114 516
rect 122 508 134 516
rect 142 508 154 516
rect 162 508 174 516
rect 182 508 418 516
rect 426 508 438 516
rect 446 508 458 516
rect 466 508 478 516
rect 486 508 498 516
rect 506 508 518 516
rect 526 508 538 516
rect 546 508 558 516
rect 566 508 578 516
rect 586 508 600 516
rect 0 492 600 508
rect 0 456 600 460
rect 0 452 286 456
rect 0 444 36 452
rect 54 444 286 452
rect 0 438 286 444
rect 314 452 600 456
rect 314 444 546 452
rect 564 444 600 452
rect 314 438 600 444
rect 0 432 600 438
rect 0 424 36 432
rect 54 430 546 432
rect 54 424 78 430
rect 0 412 78 424
rect 196 422 404 430
rect 522 424 546 430
rect 564 424 600 432
rect 0 404 36 412
rect 54 404 78 412
rect 0 392 78 404
rect 106 392 494 422
rect 522 412 600 424
rect 522 404 546 412
rect 564 404 600 412
rect 522 392 600 404
rect 0 384 36 392
rect 54 388 291 392
rect 54 384 78 388
rect 0 372 78 384
rect 0 364 36 372
rect 54 364 78 372
rect 0 352 78 364
rect 106 384 291 388
rect 309 388 546 392
rect 309 384 494 388
rect 106 358 494 384
rect 522 384 546 388
rect 564 384 600 392
rect 522 372 600 384
rect 522 364 546 372
rect 564 364 600 372
rect 0 344 36 352
rect 54 350 78 352
rect 236 350 364 358
rect 522 352 600 364
rect 522 350 546 352
rect 54 344 546 350
rect 564 344 600 352
rect 0 332 600 344
rect 0 324 36 332
rect 54 324 546 332
rect 564 324 600 332
rect 0 312 600 324
rect 0 304 36 312
rect 54 310 546 312
rect 54 304 100 310
rect 0 300 100 304
rect 500 304 546 310
rect 564 304 600 312
rect 500 300 600 304
rect 0 298 600 300
rect 0 292 78 298
rect 0 284 36 292
rect 54 284 78 292
rect 236 290 364 298
rect 522 292 600 298
rect 0 272 78 284
rect 0 264 36 272
rect 54 264 78 272
rect 0 252 78 264
rect 0 244 36 252
rect 54 244 78 252
rect 0 232 78 244
rect 0 224 36 232
rect 54 224 78 232
rect 106 264 494 290
rect 106 256 291 264
rect 309 256 494 264
rect 106 228 494 256
rect 522 284 546 292
rect 564 284 600 292
rect 522 272 600 284
rect 522 264 546 272
rect 564 264 600 272
rect 522 252 600 264
rect 522 244 546 252
rect 564 244 600 252
rect 522 232 600 244
rect 0 220 78 224
rect 236 220 364 228
rect 522 224 546 232
rect 564 224 600 232
rect 522 220 600 224
rect 0 212 600 220
rect 0 204 36 212
rect 54 204 546 212
rect 564 204 600 212
rect 0 192 600 204
rect 0 184 36 192
rect 54 184 546 192
rect 564 184 600 192
rect 0 172 600 184
rect 0 164 36 172
rect 54 168 546 172
rect 54 164 78 168
rect 0 152 78 164
rect 236 160 364 168
rect 522 164 546 168
rect 564 164 600 172
rect 0 144 36 152
rect 54 144 78 152
rect 0 132 78 144
rect 0 124 36 132
rect 54 124 78 132
rect 0 112 78 124
rect 0 104 36 112
rect 54 104 78 112
rect 0 92 78 104
rect 106 136 494 150
rect 106 128 291 136
rect 309 128 494 136
rect 106 120 494 128
rect 106 112 291 120
rect 309 112 494 120
rect 106 104 494 112
rect 106 98 291 104
rect 0 84 36 92
rect 54 90 78 92
rect 196 96 291 98
rect 309 98 494 104
rect 522 152 600 164
rect 522 144 546 152
rect 564 144 600 152
rect 522 132 600 144
rect 522 124 546 132
rect 564 124 600 132
rect 522 112 600 124
rect 522 104 546 112
rect 564 104 600 112
rect 309 96 404 98
rect 196 90 404 96
rect 522 92 600 104
rect 522 90 546 92
rect 54 84 546 90
rect 564 84 600 92
rect 0 72 600 84
rect 0 64 36 72
rect 54 66 546 72
rect 54 64 195 66
rect 0 62 195 64
rect 0 52 98 62
rect 0 44 36 52
rect 84 44 98 52
rect 0 34 98 44
rect 106 34 118 62
rect 126 34 138 62
rect 146 34 158 62
rect 166 34 178 62
rect 186 34 195 62
rect 405 64 546 66
rect 564 64 600 72
rect 405 62 600 64
rect 0 0 195 34
rect 204 30 206 58
rect 394 30 396 58
rect 204 0 396 30
rect 405 34 414 62
rect 422 34 434 62
rect 442 34 454 62
rect 462 34 474 62
rect 482 34 494 62
rect 502 52 600 62
rect 502 44 516 52
rect 564 44 600 52
rect 502 34 600 44
rect 405 0 600 34
use PadBox  PadBox_0
timestamp 1570494029
transform 1 0 40 0 1 1480
box 0 0 520 520
<< labels >>
flabel nwell 600 -6 600 -6 6 FreeSans 16 0 0 0 VddNW
flabel nwell 0 -6 0 -6 4 FreeSans 16 0 0 0 VddNW
flabel nwell 600 -6 600 -6 6 FreeSans 16 0 0 0 VddNW
flabel nwell 0 -6 0 -6 4 FreeSans 16 0 0 0 VddNW
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 VddAct
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 VddAct
flabel psubstratepdiff 0 686 0 686 4 FreeSans 16 0 0 0 GndAct
flabel psubstratepdiff 600 686 600 686 6 FreeSans 16 0 0 0 GndAct
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 VddAct
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 VddAct
flabel psubstratepdiff 0 686 0 686 4 FreeSans 16 0 0 0 GndAct
flabel psubstratepdiff 600 686 600 686 6 FreeSans 16 0 0 0 GndAct
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 688 600 688 6 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 688 0 688 4 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 880 0 880 4 FreeSans 16 0 0 0 VddM2A
flabel metal2 600 880 600 880 6 FreeSans 16 0 0 0 VddM2A
flabel metal2 0 492 0 492 4 FreeSans 16 0 0 0 VddM2B
flabel metal2 600 492 600 492 6 FreeSans 16 0 0 0 VddM2B
flabel metal2 204 0 204 0 4 FreeSans 64 0 0 0 DATA
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 688 600 688 6 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 688 0 688 4 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 880 0 880 4 FreeSans 16 0 0 0 VddM2A
flabel metal2 600 880 600 880 6 FreeSans 16 0 0 0 VddM2A
flabel metal2 0 492 0 492 4 FreeSans 16 0 0 0 VddM2B
flabel metal2 600 492 600 492 6 FreeSans 16 0 0 0 VddM2B
<< properties >>
string path 459.000 0.000 891.000 0.000 891.000 130.500 459.000 130.500 459.000 0.000 
<< end >>
