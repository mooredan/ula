magic
tech amic5n
timestamp 1622386505
<< metal1 >>
rect -120 1555 -30 1660
rect 30 1555 120 1660
rect 180 1555 270 1660
rect 330 1555 420 1660
rect 480 1555 570 1660
rect 630 1555 720 1660
rect 780 1555 870 1660
rect 930 1555 1020 1660
rect 1080 1555 1170 1660
rect -120 -250 -30 -115
rect 30 -250 120 -115
rect 180 -250 270 -115
rect 330 -250 420 -115
rect 480 -250 570 -115
rect 630 -250 720 -115
rect 780 -250 870 -115
rect 930 -250 1020 -115
rect 1080 -250 1170 -115
rect 1230 -250 1320 -115
<< metal2 >>
rect -125 1555 1350 1645
rect -125 1395 1350 1485
rect -125 1235 1350 1325
rect -125 1075 1350 1165
rect -125 915 1350 1005
rect -125 755 1350 845
rect -125 595 1350 685
rect -125 435 1350 525
rect -125 275 1350 365
rect -125 115 1350 205
rect -125 -45 1350 45
rect -125 -205 1350 -115
<< bb >>
rect 0 1550 450 1660
rect 600 1550 1050 1660
rect 0 0 1200 1440
rect 0 -255 450 -115
<< end >>
