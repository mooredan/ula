magic
tech amic5n
timestamp 1608317705
<< nwell >>
rect -120 810 1650 1950
<< ntransistor >>
rect 630 120 690 630
<< ptransistor >>
rect 600 990 660 1770
rect 870 990 930 1770
<< ndiffusion >>
rect 510 120 630 630
rect 690 120 810 630
<< pdiffusion >>
rect 420 990 600 1770
rect 660 990 870 1770
rect 930 990 1140 1770
<< polysilicon >>
rect 600 1770 660 1830
rect 870 1770 930 1830
rect 600 930 660 990
rect 870 930 930 990
rect 630 630 690 810
rect 630 60 690 120
<< metal1 >>
rect 0 1800 1530 1890
rect 0 1620 510 1710
rect 1110 1620 1530 1710
rect 0 1440 420 1530
rect 1110 1440 1530 1530
rect 0 1260 420 1350
rect 1110 1260 1530 1350
rect 0 1080 1530 1170
rect 0 900 1530 990
rect 0 720 300 810
rect 1230 720 1530 810
rect 0 540 510 630
rect 930 540 1530 630
rect 0 360 1530 450
rect 0 180 1530 270
rect 0 0 1530 90
<< labels >>
flabel metal1  0 0 0 0 2 FreeSans 400 0 0 0 Gnd
port 3 ne
flabel nwell  0 810 0 810 2 FreeSans 400 0 0 0 Vdd
flabel metal1  0 1800 0 1800 2 FreeSans 400 0 0 0 Vdd
port 2 ne
<< checkpaint >>
rect -130 -10 1660 1960
<< end >>
