magic
tech amic5n
timestamp 1621863012
<< nwell >>
rect -105 805 495 2455
<< ntransistor >>
rect 165 95 225 655
<< ptransistor >>
rect 165 955 225 2305
<< nselect >>
rect 0 0 390 685
<< pselect >>
rect 0 925 390 2400
<< ndiffusion >>
rect 45 625 165 655
rect 45 575 75 625
rect 125 575 165 625
rect 45 475 165 575
rect 45 425 75 475
rect 125 425 165 475
rect 45 375 165 425
rect 45 325 75 375
rect 125 325 165 375
rect 45 275 165 325
rect 45 225 75 275
rect 125 225 165 275
rect 45 175 165 225
rect 45 125 75 175
rect 125 125 165 175
rect 45 95 165 125
rect 225 625 345 655
rect 225 575 265 625
rect 315 575 345 625
rect 225 475 345 575
rect 225 425 265 475
rect 315 425 345 475
rect 225 375 345 425
rect 225 325 265 375
rect 315 325 345 375
rect 225 275 345 325
rect 225 225 265 275
rect 315 225 345 275
rect 225 175 345 225
rect 225 125 265 175
rect 315 125 345 175
rect 225 95 345 125
<< pdiffusion >>
rect 45 2275 165 2305
rect 45 2225 75 2275
rect 125 2225 165 2275
rect 45 2135 165 2225
rect 45 2085 75 2135
rect 125 2085 165 2135
rect 45 2035 165 2085
rect 45 1985 75 2035
rect 125 1985 165 2035
rect 45 1935 165 1985
rect 45 1885 75 1935
rect 125 1885 165 1935
rect 45 1835 165 1885
rect 45 1785 75 1835
rect 125 1785 165 1835
rect 45 1735 165 1785
rect 45 1685 75 1735
rect 125 1685 165 1735
rect 45 1635 165 1685
rect 45 1585 75 1635
rect 125 1585 165 1635
rect 45 1535 165 1585
rect 45 1485 75 1535
rect 125 1485 165 1535
rect 45 1435 165 1485
rect 45 1385 75 1435
rect 125 1385 165 1435
rect 45 1335 165 1385
rect 45 1285 75 1335
rect 125 1285 165 1335
rect 45 1235 165 1285
rect 45 1185 75 1235
rect 125 1185 165 1235
rect 45 1135 165 1185
rect 45 1085 75 1135
rect 125 1085 165 1135
rect 45 1035 165 1085
rect 45 985 75 1035
rect 125 985 165 1035
rect 45 955 165 985
rect 225 2275 345 2305
rect 225 2225 265 2275
rect 315 2225 345 2275
rect 225 2135 345 2225
rect 225 2085 265 2135
rect 315 2085 345 2135
rect 225 2035 345 2085
rect 225 1985 265 2035
rect 315 1985 345 2035
rect 225 1935 345 1985
rect 225 1885 265 1935
rect 315 1885 345 1935
rect 225 1835 345 1885
rect 225 1785 265 1835
rect 315 1785 345 1835
rect 225 1735 345 1785
rect 225 1685 265 1735
rect 315 1685 345 1735
rect 225 1635 345 1685
rect 225 1585 265 1635
rect 315 1585 345 1635
rect 225 1535 345 1585
rect 225 1485 265 1535
rect 315 1485 345 1535
rect 225 1435 345 1485
rect 225 1385 265 1435
rect 315 1385 345 1435
rect 225 1335 345 1385
rect 225 1285 265 1335
rect 315 1285 345 1335
rect 225 1235 345 1285
rect 225 1185 265 1235
rect 315 1185 345 1235
rect 225 1135 345 1185
rect 225 1085 265 1135
rect 315 1085 345 1135
rect 225 1035 345 1085
rect 225 985 265 1035
rect 315 985 345 1035
rect 225 955 345 985
<< ndcontact >>
rect 75 575 125 625
rect 75 425 125 475
rect 75 325 125 375
rect 75 225 125 275
rect 75 125 125 175
rect 265 575 315 625
rect 265 425 315 475
rect 265 325 315 375
rect 265 225 315 275
rect 265 125 315 175
<< pdcontact >>
rect 75 2225 125 2275
rect 75 2085 125 2135
rect 75 1985 125 2035
rect 75 1885 125 1935
rect 75 1785 125 1835
rect 75 1685 125 1735
rect 75 1585 125 1635
rect 75 1485 125 1535
rect 75 1385 125 1435
rect 75 1285 125 1335
rect 75 1185 125 1235
rect 75 1085 125 1135
rect 75 985 125 1035
rect 265 2225 315 2275
rect 265 2085 315 2135
rect 265 1985 315 2035
rect 265 1885 315 1935
rect 265 1785 315 1835
rect 265 1685 315 1735
rect 265 1585 315 1635
rect 265 1485 315 1535
rect 265 1385 315 1435
rect 265 1285 315 1335
rect 265 1185 315 1235
rect 265 1085 315 1135
rect 265 985 315 1035
<< polysilicon >>
rect 165 2305 225 2370
rect 165 845 225 955
rect 55 825 225 845
rect 55 775 75 825
rect 125 775 225 825
rect 55 755 225 775
rect 165 655 225 755
rect 165 30 225 95
<< polycontact >>
rect 75 775 125 825
<< metal1 >>
rect 0 2355 390 2445
rect 55 2275 145 2355
rect 55 2225 75 2275
rect 125 2225 145 2275
rect 55 2135 145 2225
rect 55 2085 75 2135
rect 125 2085 145 2135
rect 55 2035 145 2085
rect 55 1985 75 2035
rect 125 1985 145 2035
rect 55 1935 145 1985
rect 55 1885 75 1935
rect 125 1885 145 1935
rect 55 1835 145 1885
rect 55 1785 75 1835
rect 125 1785 145 1835
rect 55 1735 145 1785
rect 55 1685 75 1735
rect 125 1685 145 1735
rect 55 1635 145 1685
rect 55 1585 75 1635
rect 125 1585 145 1635
rect 55 1535 145 1585
rect 55 1485 75 1535
rect 125 1485 145 1535
rect 55 1435 145 1485
rect 55 1385 75 1435
rect 125 1385 145 1435
rect 55 1335 145 1385
rect 55 1285 75 1335
rect 125 1285 145 1335
rect 55 1235 145 1285
rect 55 1185 75 1235
rect 125 1185 145 1235
rect 55 1135 145 1185
rect 55 1085 75 1135
rect 125 1085 145 1135
rect 55 1035 145 1085
rect 55 985 75 1035
rect 125 985 145 1035
rect 55 965 145 985
rect 245 2275 335 2295
rect 245 2225 265 2275
rect 315 2225 335 2275
rect 245 2135 335 2225
rect 245 2085 265 2135
rect 315 2085 335 2135
rect 245 2035 335 2085
rect 245 1985 265 2035
rect 315 1985 335 2035
rect 245 1935 335 1985
rect 245 1885 265 1935
rect 315 1885 335 1935
rect 245 1835 335 1885
rect 245 1785 265 1835
rect 315 1785 335 1835
rect 245 1735 335 1785
rect 245 1685 265 1735
rect 315 1685 335 1735
rect 245 1635 335 1685
rect 245 1585 265 1635
rect 315 1585 335 1635
rect 245 1535 335 1585
rect 245 1485 265 1535
rect 315 1485 335 1535
rect 245 1435 335 1485
rect 245 1385 265 1435
rect 315 1385 335 1435
rect 245 1335 335 1385
rect 245 1285 265 1335
rect 315 1285 335 1335
rect 245 1235 335 1285
rect 245 1185 265 1235
rect 315 1185 335 1235
rect 245 1135 335 1185
rect 245 1085 265 1135
rect 315 1085 335 1135
rect 245 1035 335 1085
rect 245 985 265 1035
rect 315 985 335 1035
rect 55 825 145 845
rect 55 775 75 825
rect 125 775 145 825
rect 55 755 145 775
rect 55 625 145 645
rect 55 575 75 625
rect 125 575 145 625
rect 55 475 145 575
rect 55 425 75 475
rect 125 425 145 475
rect 55 375 145 425
rect 55 325 75 375
rect 125 325 145 375
rect 55 275 145 325
rect 55 225 75 275
rect 125 225 145 275
rect 55 175 145 225
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 245 625 335 985
rect 245 575 265 625
rect 315 575 335 625
rect 245 475 335 575
rect 245 425 265 475
rect 315 425 335 475
rect 245 375 335 425
rect 245 325 265 375
rect 315 325 335 375
rect 245 275 335 325
rect 245 225 265 275
rect 315 225 335 275
rect 245 175 335 225
rect 245 125 265 175
rect 315 125 335 175
rect 245 105 335 125
rect 0 -45 390 45
<< labels >>
flabel metal1 s 275 725 275 725 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 75 -25 75 -25 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 65 2375 65 2375 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 75 765 75 765 2 FreeSans 400 0 0 0 a
port 2 ne
flabel nwell 365 855 365 855 2 FreeSans 400 0 0 0 vdd
<< end >>
