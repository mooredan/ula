magic
tech scmos
timestamp 1606793110
<< nwell >>
rect -120 870 600 2430
<< ntransistor >>
rect 210 120 270 690
<< ptransistor >>
rect 210 1050 270 2250
<< nselect >>
rect 0 60 480 750
<< pselect >>
rect 0 990 480 2310
<< ndiffusion >>
rect 60 655 210 690
rect 60 605 95 655
rect 145 605 210 655
rect 60 505 210 605
rect 60 455 95 505
rect 145 455 210 505
rect 60 355 210 455
rect 60 305 95 355
rect 145 305 210 355
rect 60 205 210 305
rect 60 155 95 205
rect 145 155 210 205
rect 60 120 210 155
rect 270 655 420 690
rect 270 605 335 655
rect 385 605 420 655
rect 270 445 420 605
rect 270 395 335 445
rect 385 395 420 445
rect 270 265 420 395
rect 270 215 335 265
rect 385 215 420 265
rect 270 120 420 215
<< pdiffusion >>
rect 60 2215 210 2250
rect 60 2165 95 2215
rect 145 2165 210 2215
rect 60 2035 210 2165
rect 60 1985 95 2035
rect 145 1985 210 2035
rect 60 1885 210 1985
rect 60 1835 95 1885
rect 145 1835 210 1885
rect 60 1735 210 1835
rect 60 1685 95 1735
rect 145 1685 210 1735
rect 60 1585 210 1685
rect 60 1535 95 1585
rect 145 1535 210 1585
rect 60 1435 210 1535
rect 60 1385 95 1435
rect 145 1385 210 1435
rect 60 1285 210 1385
rect 60 1235 95 1285
rect 145 1235 210 1285
rect 60 1135 210 1235
rect 60 1085 95 1135
rect 145 1085 210 1135
rect 60 1050 210 1085
rect 270 2155 420 2250
rect 270 2105 335 2155
rect 385 2105 420 2155
rect 270 2005 420 2105
rect 270 1955 335 2005
rect 385 1955 420 2005
rect 270 1825 420 1955
rect 270 1775 335 1825
rect 385 1775 420 1825
rect 270 1645 420 1775
rect 270 1595 335 1645
rect 385 1595 420 1645
rect 270 1465 420 1595
rect 270 1415 335 1465
rect 385 1415 420 1465
rect 270 1285 420 1415
rect 270 1235 335 1285
rect 385 1235 420 1285
rect 270 1135 420 1235
rect 270 1085 335 1135
rect 385 1085 420 1135
rect 270 1050 420 1085
<< ndcontact >>
rect 95 605 145 655
rect 95 455 145 505
rect 95 305 145 355
rect 95 155 145 205
rect 335 605 385 655
rect 335 395 385 445
rect 335 215 385 265
<< pdcontact >>
rect 95 2165 145 2215
rect 95 1985 145 2035
rect 95 1835 145 1885
rect 95 1685 145 1735
rect 95 1535 145 1585
rect 95 1385 145 1435
rect 95 1235 145 1285
rect 95 1085 145 1135
rect 335 2105 385 2155
rect 335 1955 385 2005
rect 335 1775 385 1825
rect 335 1595 385 1645
rect 335 1415 385 1465
rect 335 1235 385 1285
rect 335 1085 385 1135
<< polysilicon >>
rect 210 2250 270 2320
rect 210 960 270 1050
rect 60 895 270 960
rect 60 845 125 895
rect 175 845 270 895
rect 60 780 270 845
rect 210 690 270 780
rect 210 50 270 120
<< polycontact >>
rect 125 845 175 895
<< metal1 >>
rect 0 2280 480 2370
rect 60 2215 180 2280
rect 60 2165 95 2215
rect 145 2165 180 2215
rect 60 2035 180 2165
rect 60 1985 95 2035
rect 145 1985 180 2035
rect 60 1885 180 1985
rect 60 1835 95 1885
rect 145 1835 180 1885
rect 60 1735 180 1835
rect 60 1685 95 1735
rect 145 1685 180 1735
rect 60 1585 180 1685
rect 60 1535 95 1585
rect 145 1535 180 1585
rect 60 1435 180 1535
rect 60 1385 95 1435
rect 145 1385 180 1435
rect 60 1285 180 1385
rect 60 1235 95 1285
rect 145 1235 180 1285
rect 60 1135 180 1235
rect 60 1085 95 1135
rect 145 1085 180 1135
rect 60 1050 180 1085
rect 300 2155 420 2190
rect 300 2105 335 2155
rect 385 2105 420 2155
rect 300 2005 420 2105
rect 300 1955 335 2005
rect 385 1955 420 2005
rect 300 1825 420 1955
rect 300 1775 335 1825
rect 385 1775 420 1825
rect 300 1645 420 1775
rect 300 1595 335 1645
rect 385 1595 420 1645
rect 300 1465 420 1595
rect 300 1415 335 1465
rect 385 1415 420 1465
rect 300 1285 420 1415
rect 300 1235 335 1285
rect 385 1235 420 1285
rect 300 1135 420 1235
rect 300 1085 335 1135
rect 385 1085 420 1135
rect 90 895 210 930
rect 90 845 125 895
rect 175 845 210 895
rect 90 810 210 845
rect 60 655 180 690
rect 60 605 95 655
rect 145 605 180 655
rect 60 505 180 605
rect 60 455 95 505
rect 145 455 180 505
rect 60 355 180 455
rect 60 305 95 355
rect 145 305 180 355
rect 60 205 180 305
rect 60 155 95 205
rect 145 155 180 205
rect 300 655 420 1085
rect 300 605 335 655
rect 385 605 420 655
rect 300 445 420 605
rect 300 395 335 445
rect 385 395 420 445
rect 300 265 420 395
rect 300 215 335 265
rect 385 215 420 265
rect 300 180 420 215
rect 60 90 180 155
rect 0 0 480 90
<< labels >>
flabel nwell 0 930 0 930 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 30 30 30 30 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 30 2310 30 2310 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 360 810 360 810 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 150 870 150 870 2 FreeSans 400 0 0 0 a
port 2 ne
<< end >>
