magic
tech amic5n
timestamp 1624310457
<< nwell >>
rect -130 550 1330 1495
<< ntransistor >>
rect 225 95 285 400
rect 615 125 675 400
rect 805 125 865 400
rect 995 125 1055 400
<< ptransistor >>
rect 225 705 285 1345
rect 615 705 675 1290
rect 805 705 865 1290
rect 995 705 1055 1290
<< nselect >>
rect -10 0 1210 430
<< pselect >>
rect -10 670 1210 1440
<< ndiffusion >>
rect 105 370 225 400
rect 105 320 135 370
rect 185 320 225 370
rect 105 175 225 320
rect 105 125 135 175
rect 185 125 225 175
rect 105 95 225 125
rect 285 370 405 400
rect 285 320 325 370
rect 375 320 405 370
rect 285 175 405 320
rect 285 125 325 175
rect 375 125 405 175
rect 495 370 615 400
rect 495 320 525 370
rect 575 320 615 370
rect 495 205 615 320
rect 495 155 525 205
rect 575 155 615 205
rect 495 125 615 155
rect 675 370 805 400
rect 675 320 715 370
rect 765 320 805 370
rect 675 205 805 320
rect 675 155 715 205
rect 765 155 805 205
rect 675 125 805 155
rect 865 345 995 400
rect 865 295 905 345
rect 955 295 995 345
rect 865 205 995 295
rect 865 155 905 205
rect 955 155 995 205
rect 865 125 995 155
rect 1055 370 1175 400
rect 1055 320 1095 370
rect 1145 320 1175 370
rect 1055 205 1175 320
rect 1055 155 1095 205
rect 1145 155 1175 205
rect 1055 125 1175 155
rect 285 95 405 125
<< pdiffusion >>
rect 105 1315 225 1345
rect 105 1265 135 1315
rect 185 1265 225 1315
rect 105 1215 225 1265
rect 105 1165 135 1215
rect 185 1165 225 1215
rect 105 1115 225 1165
rect 105 1065 135 1115
rect 185 1065 225 1115
rect 105 1015 225 1065
rect 105 965 135 1015
rect 185 965 225 1015
rect 105 915 225 965
rect 105 865 135 915
rect 185 865 225 915
rect 105 815 225 865
rect 105 765 135 815
rect 185 765 225 815
rect 105 705 225 765
rect 285 1315 405 1345
rect 285 1265 325 1315
rect 375 1265 405 1315
rect 285 1185 405 1265
rect 285 1135 325 1185
rect 375 1135 405 1185
rect 285 1085 405 1135
rect 285 1035 325 1085
rect 375 1035 405 1085
rect 285 985 405 1035
rect 285 935 325 985
rect 375 935 405 985
rect 285 885 405 935
rect 285 835 325 885
rect 375 835 405 885
rect 285 785 405 835
rect 285 735 325 785
rect 375 735 405 785
rect 285 705 405 735
rect 495 1260 615 1290
rect 495 1210 525 1260
rect 575 1210 615 1260
rect 495 1115 615 1210
rect 495 1065 525 1115
rect 575 1065 615 1115
rect 495 1015 615 1065
rect 495 965 525 1015
rect 575 965 615 1015
rect 495 915 615 965
rect 495 865 525 915
rect 575 865 615 915
rect 495 815 615 865
rect 495 765 525 815
rect 575 765 615 815
rect 495 705 615 765
rect 675 1260 805 1290
rect 675 1210 715 1260
rect 765 1210 805 1260
rect 675 1080 805 1210
rect 675 1030 715 1080
rect 765 1030 805 1080
rect 675 980 805 1030
rect 675 930 715 980
rect 765 930 805 980
rect 675 825 805 930
rect 675 775 715 825
rect 765 775 805 825
rect 675 705 805 775
rect 865 1260 995 1290
rect 865 1210 905 1260
rect 955 1210 995 1260
rect 865 1115 995 1210
rect 865 1065 905 1115
rect 955 1065 995 1115
rect 865 975 995 1065
rect 865 925 905 975
rect 955 925 995 975
rect 865 705 995 925
rect 1055 1260 1175 1290
rect 1055 1210 1095 1260
rect 1145 1210 1175 1260
rect 1055 1085 1175 1210
rect 1055 1035 1095 1085
rect 1145 1035 1175 1085
rect 1055 985 1175 1035
rect 1055 935 1095 985
rect 1145 935 1175 985
rect 1055 885 1175 935
rect 1055 835 1095 885
rect 1145 835 1175 885
rect 1055 785 1175 835
rect 1055 735 1095 785
rect 1145 735 1175 785
rect 1055 705 1175 735
<< ndcontact >>
rect 135 320 185 370
rect 135 125 185 175
rect 325 320 375 370
rect 325 125 375 175
rect 525 320 575 370
rect 525 155 575 205
rect 715 320 765 370
rect 715 155 765 205
rect 905 295 955 345
rect 905 155 955 205
rect 1095 320 1145 370
rect 1095 155 1145 205
<< pdcontact >>
rect 135 1265 185 1315
rect 135 1165 185 1215
rect 135 1065 185 1115
rect 135 965 185 1015
rect 135 865 185 915
rect 135 765 185 815
rect 325 1265 375 1315
rect 325 1135 375 1185
rect 325 1035 375 1085
rect 325 935 375 985
rect 325 835 375 885
rect 325 735 375 785
rect 525 1210 575 1260
rect 525 1065 575 1115
rect 525 965 575 1015
rect 525 865 575 915
rect 525 765 575 815
rect 715 1210 765 1260
rect 715 1030 765 1080
rect 715 930 765 980
rect 715 775 765 825
rect 905 1210 955 1260
rect 905 1065 955 1115
rect 905 925 955 975
rect 1095 1210 1145 1260
rect 1095 1035 1145 1085
rect 1095 935 1145 985
rect 1095 835 1145 885
rect 1095 735 1145 785
<< polysilicon >>
rect 225 1345 285 1410
rect 615 1290 675 1355
rect 805 1290 865 1355
rect 995 1290 1055 1355
rect 225 685 285 705
rect 615 685 675 705
rect 805 685 865 705
rect 995 685 1055 705
rect 115 665 285 685
rect 115 615 135 665
rect 185 615 285 665
rect 115 595 285 615
rect 505 665 1055 685
rect 505 615 525 665
rect 575 615 625 665
rect 675 615 725 665
rect 775 615 825 665
rect 875 615 925 665
rect 975 615 1055 665
rect 505 595 1055 615
rect 225 400 285 595
rect 615 400 675 595
rect 805 400 865 595
rect 995 400 1055 595
rect 225 30 285 95
rect 615 60 675 125
rect 805 60 865 125
rect 995 60 1055 125
<< polycontact >>
rect 135 615 185 665
rect 525 615 575 665
rect 625 615 675 665
rect 725 615 775 665
rect 825 615 875 665
rect 925 615 975 665
<< metal1 >>
rect 0 1395 1200 1485
rect 115 1315 205 1395
rect 115 1265 135 1315
rect 185 1265 205 1315
rect 115 1215 205 1265
rect 115 1165 135 1215
rect 185 1165 205 1215
rect 115 1115 205 1165
rect 115 1065 135 1115
rect 185 1065 205 1115
rect 115 1015 205 1065
rect 115 965 135 1015
rect 185 965 205 1015
rect 115 915 205 965
rect 115 865 135 915
rect 185 865 205 915
rect 115 815 205 865
rect 115 765 135 815
rect 185 765 205 815
rect 115 745 205 765
rect 305 1315 395 1335
rect 305 1265 325 1315
rect 375 1265 395 1315
rect 305 1185 395 1265
rect 305 1135 325 1185
rect 375 1135 395 1185
rect 305 1085 395 1135
rect 305 1035 325 1085
rect 375 1035 395 1085
rect 305 985 395 1035
rect 305 935 325 985
rect 375 935 395 985
rect 305 885 395 935
rect 305 835 325 885
rect 375 835 395 885
rect 305 785 395 835
rect 305 735 325 785
rect 375 735 395 785
rect 505 1260 595 1395
rect 505 1210 525 1260
rect 575 1210 595 1260
rect 505 1115 595 1210
rect 505 1065 525 1115
rect 575 1065 595 1115
rect 505 1015 595 1065
rect 505 965 525 1015
rect 575 965 595 1015
rect 505 915 595 965
rect 505 865 525 915
rect 575 865 595 915
rect 505 815 595 865
rect 505 765 525 815
rect 575 765 595 815
rect 505 745 595 765
rect 695 1260 785 1280
rect 695 1210 715 1260
rect 765 1210 785 1260
rect 695 1080 785 1210
rect 695 1030 715 1080
rect 765 1030 785 1080
rect 695 980 785 1030
rect 695 930 715 980
rect 765 930 785 980
rect 695 845 785 930
rect 885 1260 975 1395
rect 885 1210 905 1260
rect 955 1210 975 1260
rect 885 1115 975 1210
rect 885 1065 905 1115
rect 955 1065 975 1115
rect 885 975 975 1065
rect 885 925 905 975
rect 955 925 975 975
rect 885 905 975 925
rect 1075 1260 1165 1280
rect 1075 1210 1095 1260
rect 1145 1210 1165 1260
rect 1075 1085 1165 1210
rect 1075 1035 1095 1085
rect 1145 1035 1165 1085
rect 1075 985 1165 1035
rect 1075 935 1095 985
rect 1145 935 1165 985
rect 1075 885 1165 935
rect 1075 845 1095 885
rect 695 835 1095 845
rect 1145 835 1165 885
rect 695 825 1165 835
rect 695 775 715 825
rect 765 785 1165 825
rect 765 775 1095 785
rect 695 755 1095 775
rect 305 685 395 735
rect 1075 735 1095 755
rect 1145 735 1165 785
rect 115 665 205 685
rect 115 615 135 665
rect 185 615 205 665
rect 115 595 205 615
rect 305 665 995 685
rect 305 615 525 665
rect 575 615 625 665
rect 675 615 725 665
rect 775 615 825 665
rect 875 615 925 665
rect 975 615 995 665
rect 305 595 995 615
rect 115 370 205 390
rect 115 320 135 370
rect 185 320 205 370
rect 115 175 205 320
rect 115 125 135 175
rect 185 125 205 175
rect 115 45 205 125
rect 305 370 395 595
rect 1075 525 1165 735
rect 695 435 1165 525
rect 305 320 325 370
rect 375 320 395 370
rect 305 175 395 320
rect 305 125 325 175
rect 375 125 395 175
rect 305 105 395 125
rect 505 370 595 390
rect 505 320 525 370
rect 575 320 595 370
rect 505 205 595 320
rect 505 155 525 205
rect 575 155 595 205
rect 505 45 595 155
rect 695 370 785 435
rect 695 320 715 370
rect 765 320 785 370
rect 1075 370 1165 435
rect 695 205 785 320
rect 695 155 715 205
rect 765 155 785 205
rect 695 135 785 155
rect 885 345 975 365
rect 885 295 905 345
rect 955 295 975 345
rect 885 205 975 295
rect 885 155 905 205
rect 955 155 975 205
rect 885 45 975 155
rect 1075 320 1095 370
rect 1145 320 1165 370
rect 1075 205 1165 320
rect 1075 155 1095 205
rect 1145 155 1165 205
rect 1075 135 1165 155
rect 0 -45 1200 45
<< labels >>
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 2 ne
flabel metal1 s 5 5 5 5 2 FreeSans 200 0 0 0 vss
port 3 ne
flabel metal1 s 1115 485 1115 485 2 FreeSans 400 0 0 0 z
port 0 ne
flabel nwell 405 560 405 560 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 135 605 135 605 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 330 470 330 470 2 FreeSans 200 0 0 0 x1
<< properties >>
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
<< end >>
