magic
tech amic5n
timestamp 1625244951
<< nwell >>
rect -130 550 1180 1495
rect 105 150 945 550
<< polysilicon >>
rect 105 1240 945 1290
rect 105 1220 225 1240
rect 105 1170 125 1220
rect 175 1170 225 1220
rect 825 1220 945 1240
rect 105 1120 225 1170
rect 825 1170 875 1220
rect 925 1170 945 1220
rect 105 1070 125 1120
rect 175 1070 225 1120
rect 825 1120 945 1170
rect 825 1070 875 1120
rect 925 1070 945 1120
rect 105 1020 225 1070
rect 825 1020 945 1070
rect 105 970 125 1020
rect 175 970 225 1020
rect 105 920 225 970
rect 825 970 875 1020
rect 925 970 945 1020
rect 105 870 125 920
rect 175 870 225 920
rect 825 920 945 970
rect 105 820 225 870
rect 825 870 875 920
rect 925 870 945 920
rect 105 770 125 820
rect 175 770 225 820
rect 825 820 945 870
rect 105 720 225 770
rect 825 770 875 820
rect 925 770 945 820
rect 105 670 125 720
rect 175 670 225 720
rect 825 720 945 770
rect 105 620 225 670
rect 825 670 875 720
rect 925 670 945 720
rect 105 570 125 620
rect 175 570 225 620
rect 825 620 945 670
rect 105 520 225 570
rect 825 570 875 620
rect 925 570 945 620
rect 825 520 945 570
rect 105 470 125 520
rect 175 470 225 520
rect 825 470 875 520
rect 925 470 945 520
rect 105 420 225 470
rect 105 370 125 420
rect 175 370 225 420
rect 825 420 945 470
rect 105 320 225 370
rect 825 370 875 420
rect 925 370 945 420
rect 105 270 125 320
rect 175 270 225 320
rect 825 320 945 370
rect 105 220 225 270
rect 825 270 875 320
rect 925 270 945 320
rect 105 170 125 220
rect 175 200 225 220
rect 825 220 945 270
rect 825 200 875 220
rect 175 170 875 200
rect 925 170 945 220
rect 105 150 945 170
<< polycontact >>
rect 125 1170 175 1220
rect 875 1170 925 1220
rect 125 1070 175 1120
rect 875 1070 925 1120
rect 125 970 175 1020
rect 875 970 925 1020
rect 125 870 175 920
rect 875 870 925 920
rect 125 770 175 820
rect 875 770 925 820
rect 125 670 175 720
rect 875 670 925 720
rect 125 570 175 620
rect 875 570 925 620
rect 125 470 175 520
rect 875 470 925 520
rect 125 370 175 420
rect 875 370 925 420
rect 125 270 175 320
rect 875 270 925 320
rect 125 170 175 220
rect 875 170 925 220
<< poly2cap >>
rect 225 1180 825 1240
rect 225 1130 275 1180
rect 325 1130 385 1180
rect 435 1130 495 1180
rect 545 1130 610 1180
rect 660 1130 725 1180
rect 775 1130 825 1180
rect 225 1070 825 1130
rect 225 1020 275 1070
rect 325 1020 385 1070
rect 435 1020 495 1070
rect 545 1020 610 1070
rect 660 1020 725 1070
rect 775 1020 825 1070
rect 225 960 825 1020
rect 225 910 275 960
rect 325 910 385 960
rect 435 910 495 960
rect 545 910 610 960
rect 660 910 725 960
rect 775 910 825 960
rect 225 850 825 910
rect 225 800 275 850
rect 325 800 385 850
rect 435 800 495 850
rect 545 800 610 850
rect 660 800 725 850
rect 775 800 825 850
rect 225 740 825 800
rect 225 690 275 740
rect 325 690 385 740
rect 435 690 495 740
rect 545 690 610 740
rect 660 690 725 740
rect 775 690 825 740
rect 225 630 825 690
rect 225 580 275 630
rect 325 580 385 630
rect 435 580 495 630
rect 545 580 610 630
rect 660 580 725 630
rect 775 580 825 630
rect 225 520 825 580
rect 225 470 275 520
rect 325 470 385 520
rect 435 470 495 520
rect 545 470 610 520
rect 660 470 725 520
rect 775 470 825 520
rect 225 410 825 470
rect 225 360 275 410
rect 325 360 385 410
rect 435 360 495 410
rect 545 360 610 410
rect 660 360 725 410
rect 775 360 825 410
rect 225 300 825 360
rect 225 250 275 300
rect 325 250 385 300
rect 435 250 495 300
rect 545 250 610 300
rect 660 250 725 300
rect 775 250 825 300
rect 225 200 825 250
<< poly2capcontact >>
rect 275 1130 325 1180
rect 385 1130 435 1180
rect 495 1130 545 1180
rect 610 1130 660 1180
rect 725 1130 775 1180
rect 275 1020 325 1070
rect 385 1020 435 1070
rect 495 1020 545 1070
rect 610 1020 660 1070
rect 725 1020 775 1070
rect 275 910 325 960
rect 385 910 435 960
rect 495 910 545 960
rect 610 910 660 960
rect 725 910 775 960
rect 275 800 325 850
rect 385 800 435 850
rect 495 800 545 850
rect 610 800 660 850
rect 725 800 775 850
rect 275 690 325 740
rect 385 690 435 740
rect 495 690 545 740
rect 610 690 660 740
rect 725 690 775 740
rect 275 580 325 630
rect 385 580 435 630
rect 495 580 545 630
rect 610 580 660 630
rect 725 580 775 630
rect 275 470 325 520
rect 385 470 435 520
rect 495 470 545 520
rect 610 470 660 520
rect 725 470 775 520
rect 275 360 325 410
rect 385 360 435 410
rect 495 360 545 410
rect 610 360 660 410
rect 725 360 775 410
rect 275 250 325 300
rect 385 250 435 300
rect 495 250 545 300
rect 610 250 660 300
rect 725 250 775 300
<< metal1 >>
rect 0 1395 1050 1485
rect 165 1305 885 1395
rect 105 1220 195 1240
rect 105 1170 125 1220
rect 175 1170 195 1220
rect 105 1120 195 1170
rect 105 1070 125 1120
rect 175 1070 195 1120
rect 105 1020 195 1070
rect 105 970 125 1020
rect 175 970 195 1020
rect 105 920 195 970
rect 105 870 125 920
rect 175 870 195 920
rect 105 820 195 870
rect 105 770 125 820
rect 175 770 195 820
rect 105 720 195 770
rect 105 670 125 720
rect 175 670 195 720
rect 105 620 195 670
rect 105 570 125 620
rect 175 570 195 620
rect 105 520 195 570
rect 105 470 125 520
rect 175 470 195 520
rect 105 420 195 470
rect 105 370 125 420
rect 175 370 195 420
rect 105 320 195 370
rect 105 270 125 320
rect 175 270 195 320
rect 105 220 195 270
rect 255 1180 795 1305
rect 255 1130 275 1180
rect 325 1130 385 1180
rect 435 1130 495 1180
rect 545 1130 610 1180
rect 660 1130 725 1180
rect 775 1130 795 1180
rect 255 1070 795 1130
rect 255 1020 275 1070
rect 325 1020 385 1070
rect 435 1020 495 1070
rect 545 1020 610 1070
rect 660 1020 725 1070
rect 775 1020 795 1070
rect 255 960 795 1020
rect 255 910 275 960
rect 325 910 385 960
rect 435 910 495 960
rect 545 910 610 960
rect 660 910 725 960
rect 775 910 795 960
rect 255 850 795 910
rect 255 800 275 850
rect 325 800 385 850
rect 435 800 495 850
rect 545 800 610 850
rect 660 800 725 850
rect 775 800 795 850
rect 255 740 795 800
rect 255 690 275 740
rect 325 690 385 740
rect 435 690 495 740
rect 545 690 610 740
rect 660 690 725 740
rect 775 690 795 740
rect 255 630 795 690
rect 255 580 275 630
rect 325 580 385 630
rect 435 580 495 630
rect 545 580 610 630
rect 660 580 725 630
rect 775 580 795 630
rect 255 520 795 580
rect 255 470 275 520
rect 325 470 385 520
rect 435 470 495 520
rect 545 470 610 520
rect 660 470 725 520
rect 775 470 795 520
rect 255 410 795 470
rect 255 360 275 410
rect 325 360 385 410
rect 435 360 495 410
rect 545 360 610 410
rect 660 360 725 410
rect 775 360 795 410
rect 255 300 795 360
rect 255 250 275 300
rect 325 250 385 300
rect 435 250 495 300
rect 545 250 610 300
rect 660 250 725 300
rect 775 250 795 300
rect 255 230 795 250
rect 855 1220 945 1240
rect 855 1170 875 1220
rect 925 1170 945 1220
rect 855 1120 945 1170
rect 855 1070 875 1120
rect 925 1070 945 1120
rect 855 1020 945 1070
rect 855 970 875 1020
rect 925 970 945 1020
rect 855 920 945 970
rect 855 870 875 920
rect 925 870 945 920
rect 855 820 945 870
rect 855 770 875 820
rect 925 770 945 820
rect 855 720 945 770
rect 855 670 875 720
rect 925 670 945 720
rect 855 620 945 670
rect 855 570 875 620
rect 925 570 945 620
rect 855 520 945 570
rect 855 470 875 520
rect 925 470 945 520
rect 855 420 945 470
rect 855 370 875 420
rect 925 370 945 420
rect 855 320 945 370
rect 855 270 875 320
rect 925 270 945 320
rect 105 170 125 220
rect 175 170 195 220
rect 105 150 195 170
rect 855 220 945 270
rect 855 170 875 220
rect 925 170 945 220
rect 855 150 945 170
rect 105 45 945 150
rect 0 -45 1050 45
<< labels >>
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 0 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 1 ne
flabel nwell 5 580 5 580 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFsite core
string LEFclass CORE
string FIXED_BBOX 0 0 1050 1440
string LEFsymmetry X Y
<< end >>
