magic
tech scmos
timestamp 1606679270
<< nwell >>
rect 420 13560 10380 20430
rect -90 12540 10890 13050
rect -90 11190 10890 11700
rect -90 4320 420 11190
rect 10380 4320 10890 11190
rect -90 3810 10890 4320
<< nselect >>
rect 510 19920 10290 20340
rect 510 14070 1020 19920
rect 5100 14070 5700 19920
rect 9780 14070 10290 19920
rect 510 13650 10290 14070
rect -90 12540 10890 13050
rect -60 11220 10860 11700
rect -60 4290 390 11220
rect 1020 4830 4890 10680
rect 5910 4830 9780 10680
rect 10410 4290 10860 11220
rect -60 3840 10860 4290
rect 660 390 2220 2820
rect 8580 390 10140 2820
<< pselect >>
rect -90 20430 10890 20940
rect -90 13560 420 20430
rect 1020 14070 5100 19920
rect 5700 14070 9780 19920
rect 10380 13560 10890 20430
rect -90 13050 10890 13560
rect -90 11700 10890 12210
rect 510 10680 10290 11100
rect 510 4830 1020 10680
rect 4890 4830 5910 10680
rect 9780 4830 10290 10680
rect 510 4410 10290 4830
rect -60 3330 10860 3780
rect -60 390 390 3330
rect 10410 390 10860 3330
rect -60 -60 10860 390
<< ntransistor >>
rect 1140 10320 4770 10410
rect 1140 9000 4770 9090
rect 1140 8370 4770 8460
rect 1140 7050 4770 7140
rect 1140 6420 4770 6510
rect 1140 5100 4770 5190
rect 6030 10320 9660 10410
rect 6030 9000 9660 9090
rect 6030 8370 9660 8460
rect 6030 7050 9660 7140
rect 6030 6420 9660 6510
rect 6030 5100 9660 5190
rect 870 2520 2160 2580
rect 8640 2520 9930 2580
rect 870 2280 2160 2340
rect 8640 2280 9930 2340
rect 870 2040 2160 2100
rect 870 1800 2160 1860
rect 870 1560 2160 1620
rect 8640 2040 9930 2100
rect 8640 1800 9930 1860
rect 8640 1560 9930 1620
rect 870 1320 2160 1380
rect 870 1080 2160 1140
rect 8640 1320 9930 1380
rect 8640 1080 9930 1140
rect 870 840 2160 900
rect 870 600 2160 660
rect 8640 840 9930 900
rect 8640 600 9930 660
<< ptransistor >>
rect 1140 19560 4980 19650
rect 1140 18240 4980 18330
rect 1140 17610 4980 17700
rect 1140 16290 4980 16380
rect 1140 15660 4980 15750
rect 1140 14340 4980 14430
rect 5820 19560 9660 19650
rect 5820 18240 9660 18330
rect 5820 17610 9660 17700
rect 5820 16290 9660 16380
rect 5820 15660 9660 15750
rect 5820 14340 9660 14430
<< ndiffusion >>
rect 1020 10500 4890 10680
rect 5910 10500 9780 10680
rect 1140 10410 4770 10500
rect 1140 9090 4770 10320
rect 1140 8460 4770 9000
rect 1140 7140 4770 8370
rect 1140 6510 4770 7050
rect 1140 5190 4770 6420
rect 1140 5010 4770 5100
rect 6030 10410 9660 10500
rect 6030 9090 9660 10320
rect 6030 8460 9660 9000
rect 6030 7140 9660 8370
rect 6030 6510 9660 7050
rect 6030 5190 9660 6420
rect 6030 5010 9660 5100
rect 1020 4830 4890 5010
rect 5910 4830 9780 5010
rect 870 2580 2160 2760
rect 8640 2580 9930 2760
rect 870 2340 2160 2520
rect 870 2100 2160 2280
rect 8640 2340 9930 2520
rect 870 1860 2160 2040
rect 870 1620 2160 1800
rect 870 1380 2160 1560
rect 8640 2100 9930 2280
rect 8640 1860 9930 2040
rect 8640 1620 9930 1800
rect 870 1140 2160 1320
rect 8640 1380 9930 1560
rect 8640 1140 9930 1320
rect 870 900 2160 1080
rect 870 660 2160 840
rect 8640 900 9930 1080
rect 8640 660 9930 840
rect 870 450 2160 600
rect 8640 450 9930 600
<< pdiffusion >>
rect 1020 19740 5100 19920
rect 5700 19740 9780 19920
rect 1140 19650 4980 19740
rect 1140 18330 4980 19560
rect 1140 17700 4980 18240
rect 1140 16380 4980 17610
rect 1140 15750 4980 16290
rect 1140 14430 4980 15660
rect 1140 14250 4980 14340
rect 5820 19650 9660 19740
rect 5820 18330 9660 19560
rect 5820 17700 9660 18240
rect 5820 16380 9660 17610
rect 5820 15750 9660 16290
rect 5820 14430 9660 15660
rect 5820 14250 9660 14340
rect 1020 14070 5100 14250
rect 5700 14070 9780 14250
<< psubstratepdiff >>
rect 0 20520 10800 20850
rect 0 13470 330 20520
rect 10470 13470 10800 20520
rect 0 13140 10800 13470
rect 0 11790 10800 12120
rect 570 10680 10230 11040
rect 570 10500 1020 10680
rect 4890 10500 5910 10680
rect 9780 10500 10230 10680
rect 570 5010 900 10500
rect 5010 5010 5790 10500
rect 9900 5010 10230 10500
rect 570 4830 1020 5010
rect 4890 4830 5910 5010
rect 9780 4830 10230 5010
rect 570 4470 10230 4830
rect 0 3390 10800 3720
rect 0 330 330 3390
rect 10470 330 10800 3390
rect 0 0 10800 330
<< nsubstratendiff >>
rect 570 19920 10230 20280
rect 570 19740 1020 19920
rect 5100 19740 5700 19920
rect 9780 19740 10230 19920
rect 570 14250 900 19740
rect 5220 14250 5580 19740
rect 9900 14250 10230 19740
rect 570 14070 1020 14250
rect 5100 14070 5700 14250
rect 9780 14070 10230 14250
rect 570 13710 10230 14070
rect 0 12630 10800 12960
rect 0 11280 10800 11610
rect 0 4230 330 11280
rect 10470 4230 10800 11280
rect 0 3900 10800 4230
rect 2430 2130 8370 2460
rect 2430 1080 8370 1410
<< polysilicon >>
rect 930 19560 1140 19650
rect 4980 19560 5190 19650
rect 930 18330 1110 19560
rect 5010 18330 5190 19560
rect 930 18240 1140 18330
rect 4980 18240 5190 18330
rect 930 17700 1110 18240
rect 5010 17700 5190 18240
rect 930 17610 1140 17700
rect 4980 17610 5190 17700
rect 930 16380 1110 17610
rect 5010 16380 5190 17610
rect 930 16290 1140 16380
rect 4980 16290 5190 16380
rect 930 15750 1110 16290
rect 5010 15750 5190 16290
rect 930 15660 1140 15750
rect 4980 15660 5190 15750
rect 930 14430 1110 15660
rect 5010 14430 5190 15660
rect 930 14340 1140 14430
rect 4980 14340 5190 14430
rect 5610 19560 5820 19650
rect 9660 19560 9870 19650
rect 5610 18330 5790 19560
rect 9690 18330 9870 19560
rect 5610 18240 5820 18330
rect 9660 18240 9870 18330
rect 5610 17700 5790 18240
rect 9690 17700 9870 18240
rect 5610 17610 5820 17700
rect 9660 17610 9870 17700
rect 5610 16380 5790 17610
rect 9690 16380 9870 17610
rect 5610 16290 5820 16380
rect 9660 16290 9870 16380
rect 5610 15750 5790 16290
rect 9690 15750 9870 16290
rect 5610 15660 5820 15750
rect 9660 15660 9870 15750
rect 5610 14430 5790 15660
rect 9690 14430 9870 15660
rect 5610 14340 5820 14430
rect 9660 14340 9870 14430
rect 930 10320 1140 10410
rect 4770 10320 4980 10410
rect 930 9090 1110 10320
rect 4800 9090 4980 10320
rect 930 9000 1140 9090
rect 4770 9000 4980 9090
rect 930 8460 1110 9000
rect 4800 8460 4980 9000
rect 930 8370 1140 8460
rect 4770 8370 4980 8460
rect 930 7140 1110 8370
rect 4800 7140 4980 8370
rect 930 7050 1140 7140
rect 4770 7050 4980 7140
rect 930 6510 1110 7050
rect 4800 6510 4980 7050
rect 930 6420 1140 6510
rect 4770 6420 4980 6510
rect 930 5190 1110 6420
rect 4800 5190 4980 6420
rect 930 5100 1140 5190
rect 4770 5100 4980 5190
rect 5820 10320 6030 10410
rect 9660 10320 9870 10410
rect 5820 9090 6000 10320
rect 9690 9090 9870 10320
rect 5820 9000 6030 9090
rect 9660 9000 9870 9090
rect 5820 8460 6000 9000
rect 9690 8460 9870 9000
rect 5820 8370 6030 8460
rect 9660 8370 9870 8460
rect 5820 7140 6000 8370
rect 9690 7140 9870 8370
rect 5820 7050 6030 7140
rect 9660 7050 9870 7140
rect 5820 6510 6000 7050
rect 9690 6510 9870 7050
rect 5820 6420 6030 6510
rect 9660 6420 9870 6510
rect 5820 5190 6000 6420
rect 9690 5190 9870 6420
rect 5820 5100 6030 5190
rect 9660 5100 9870 5190
rect 660 2520 870 2580
rect 2160 2520 2280 2580
rect 660 2340 840 2520
rect 2220 2340 2280 2520
rect 8520 2520 8640 2580
rect 9930 2520 10140 2580
rect 660 2280 870 2340
rect 2160 2280 2280 2340
rect 660 2100 840 2280
rect 2220 2100 2280 2280
rect 8520 2340 8580 2520
rect 9960 2340 10140 2520
rect 8520 2280 8640 2340
rect 9930 2280 10140 2340
rect 660 2040 870 2100
rect 2160 2040 2280 2100
rect 660 1860 840 2040
rect 2220 1860 2280 2040
rect 660 1800 870 1860
rect 2160 1800 2280 1860
rect 660 1620 840 1800
rect 2220 1620 2280 1800
rect 660 1560 870 1620
rect 2160 1560 2280 1620
rect 660 1380 840 1560
rect 2220 1380 2280 1560
rect 8520 2100 8580 2280
rect 9960 2100 10140 2280
rect 8520 2040 8640 2100
rect 9930 2040 10140 2100
rect 8520 1860 8580 2040
rect 9960 1860 10140 2040
rect 8520 1800 8640 1860
rect 9930 1800 10140 1860
rect 8520 1620 8580 1800
rect 9960 1620 10140 1800
rect 8520 1560 8640 1620
rect 9930 1560 10140 1620
rect 660 1320 870 1380
rect 2160 1320 2280 1380
rect 660 1140 840 1320
rect 2220 1140 2280 1320
rect 660 1080 870 1140
rect 2160 1080 2280 1140
rect 8520 1380 8580 1560
rect 9960 1380 10140 1560
rect 8520 1320 8640 1380
rect 9930 1320 10140 1380
rect 8520 1140 8580 1320
rect 9960 1140 10140 1320
rect 8520 1080 8640 1140
rect 9930 1080 10140 1140
rect 660 900 840 1080
rect 2220 900 2280 1080
rect 660 840 870 900
rect 2160 840 2280 900
rect 660 660 840 840
rect 2220 660 2280 840
rect 660 600 870 660
rect 2160 600 2280 660
rect 8520 900 8580 1080
rect 9960 900 10140 1080
rect 8520 840 8640 900
rect 9930 840 10140 900
rect 8520 660 8580 840
rect 9960 660 10140 840
rect 8520 600 8640 660
rect 9930 600 10140 660
rect 660 450 840 600
rect 9960 450 10140 600
<< psubstratepcontact >>
rect 275 20735 325 20785
<< psubstratepcontact >>
rect 515 20735 565 20785
<< psubstratepcontact >>
rect 755 20735 805 20785
<< psubstratepcontact >>
rect 995 20735 1045 20785
<< psubstratepcontact >>
rect 1235 20735 1285 20785
<< psubstratepcontact >>
rect 1475 20735 1525 20785
<< psubstratepcontact >>
rect 1715 20735 1765 20785
<< psubstratepcontact >>
rect 1955 20735 2005 20785
<< psubstratepcontact >>
rect 2195 20735 2245 20785
<< psubstratepcontact >>
rect 2435 20735 2485 20785
<< psubstratepcontact >>
rect 2675 20735 2725 20785
<< psubstratepcontact >>
rect 2915 20735 2965 20785
<< psubstratepcontact >>
rect 3155 20735 3205 20785
<< psubstratepcontact >>
rect 3395 20735 3445 20785
<< psubstratepcontact >>
rect 4535 20735 4585 20785
<< psubstratepcontact >>
rect 4775 20735 4825 20785
<< psubstratepcontact >>
rect 5015 20735 5065 20785
<< psubstratepcontact >>
rect 5255 20735 5305 20785
<< psubstratepcontact >>
rect 5495 20735 5545 20785
<< psubstratepcontact >>
rect 5735 20735 5785 20785
<< psubstratepcontact >>
rect 5975 20735 6025 20785
<< psubstratepcontact >>
rect 6215 20735 6265 20785
<< psubstratepcontact >>
rect 7355 20735 7405 20785
<< psubstratepcontact >>
rect 7595 20735 7645 20785
<< psubstratepcontact >>
rect 7835 20735 7885 20785
<< psubstratepcontact >>
rect 8075 20735 8125 20785
<< psubstratepcontact >>
rect 8315 20735 8365 20785
<< psubstratepcontact >>
rect 8555 20735 8605 20785
<< psubstratepcontact >>
rect 8795 20735 8845 20785
<< psubstratepcontact >>
rect 9035 20735 9085 20785
<< psubstratepcontact >>
rect 9275 20735 9325 20785
<< psubstratepcontact >>
rect 9515 20735 9565 20785
<< psubstratepcontact >>
rect 9755 20735 9805 20785
<< psubstratepcontact >>
rect 9995 20735 10045 20785
<< psubstratepcontact >>
rect 10235 20735 10285 20785
<< psubstratepcontact >>
rect 10475 20735 10525 20785
<< psubstratepcontact >>
rect 275 20585 325 20635
<< psubstratepcontact >>
rect 515 20585 565 20635
<< psubstratepcontact >>
rect 755 20585 805 20635
<< psubstratepcontact >>
rect 995 20585 1045 20635
<< psubstratepcontact >>
rect 1235 20585 1285 20635
<< psubstratepcontact >>
rect 1475 20585 1525 20635
<< psubstratepcontact >>
rect 1715 20585 1765 20635
<< psubstratepcontact >>
rect 1955 20585 2005 20635
<< psubstratepcontact >>
rect 2195 20585 2245 20635
<< psubstratepcontact >>
rect 2435 20585 2485 20635
<< psubstratepcontact >>
rect 2675 20585 2725 20635
<< psubstratepcontact >>
rect 2915 20585 2965 20635
<< psubstratepcontact >>
rect 3155 20585 3205 20635
<< psubstratepcontact >>
rect 3395 20585 3445 20635
<< psubstratepcontact >>
rect 4535 20585 4585 20635
<< psubstratepcontact >>
rect 4775 20585 4825 20635
<< psubstratepcontact >>
rect 5015 20585 5065 20635
<< psubstratepcontact >>
rect 5255 20585 5305 20635
<< psubstratepcontact >>
rect 5495 20585 5545 20635
<< psubstratepcontact >>
rect 5735 20585 5785 20635
<< psubstratepcontact >>
rect 5975 20585 6025 20635
<< psubstratepcontact >>
rect 6215 20585 6265 20635
<< psubstratepcontact >>
rect 7355 20585 7405 20635
<< psubstratepcontact >>
rect 7595 20585 7645 20635
<< psubstratepcontact >>
rect 7835 20585 7885 20635
<< psubstratepcontact >>
rect 8075 20585 8125 20635
<< psubstratepcontact >>
rect 8315 20585 8365 20635
<< psubstratepcontact >>
rect 8555 20585 8605 20635
<< psubstratepcontact >>
rect 8795 20585 8845 20635
<< psubstratepcontact >>
rect 9035 20585 9085 20635
<< psubstratepcontact >>
rect 9275 20585 9325 20635
<< psubstratepcontact >>
rect 9515 20585 9565 20635
<< psubstratepcontact >>
rect 9755 20585 9805 20635
<< psubstratepcontact >>
rect 9995 20585 10045 20635
<< psubstratepcontact >>
rect 10235 20585 10285 20635
<< psubstratepcontact >>
rect 10475 20585 10525 20635
<< psubstratepcontact >>
rect 65 20345 115 20395
<< psubstratepcontact >>
rect 215 20345 265 20395
<< psubstratepcontact >>
rect 10535 20345 10585 20395
<< psubstratepcontact >>
rect 10685 20345 10735 20395
<< psubstratepcontact >>
rect 65 20105 115 20155
<< psubstratepcontact >>
rect 215 20105 265 20155
<< psubstratepcontact >>
rect 10535 20105 10585 20155
<< psubstratepcontact >>
rect 10685 20105 10735 20155
<< nsubstratencontact >>
rect 905 20045 955 20095
<< nsubstratencontact >>
rect 1235 20045 1285 20095
<< nsubstratencontact >>
rect 1535 20045 1585 20095
<< nsubstratencontact >>
rect 1835 20045 1885 20095
<< nsubstratencontact >>
rect 2135 20045 2185 20095
<< nsubstratencontact >>
rect 2435 20045 2485 20095
<< nsubstratencontact >>
rect 2735 20045 2785 20095
<< nsubstratencontact >>
rect 3035 20045 3085 20095
<< nsubstratencontact >>
rect 3335 20045 3385 20095
<< nsubstratencontact >>
rect 4505 20045 4555 20095
<< nsubstratencontact >>
rect 4805 20045 4855 20095
<< nsubstratencontact >>
rect 5945 20045 5995 20095
<< nsubstratencontact >>
rect 6245 20045 6295 20095
<< nsubstratencontact >>
rect 7415 20045 7465 20095
<< nsubstratencontact >>
rect 7715 20045 7765 20095
<< nsubstratencontact >>
rect 8015 20045 8065 20095
<< nsubstratencontact >>
rect 8315 20045 8365 20095
<< nsubstratencontact >>
rect 8615 20045 8665 20095
<< nsubstratencontact >>
rect 8915 20045 8965 20095
<< nsubstratencontact >>
rect 9215 20045 9265 20095
<< nsubstratencontact >>
rect 9515 20045 9565 20095
<< nsubstratencontact >>
rect 9815 20045 9865 20095
<< psubstratepcontact >>
rect 65 19865 115 19915
<< psubstratepcontact >>
rect 215 19865 265 19915
<< nsubstratencontact >>
rect 905 19895 955 19945
<< pdcontact >>
rect 1235 19895 1285 19945
<< pdcontact >>
rect 1535 19895 1585 19945
<< pdcontact >>
rect 1835 19895 1885 19945
<< pdcontact >>
rect 2135 19895 2185 19945
<< pdcontact >>
rect 2435 19895 2485 19945
<< pdcontact >>
rect 2735 19895 2785 19945
<< pdcontact >>
rect 3035 19895 3085 19945
<< pdcontact >>
rect 3335 19895 3385 19945
<< pdcontact >>
rect 4505 19895 4555 19945
<< pdcontact >>
rect 4805 19895 4855 19945
<< pdcontact >>
rect 5945 19895 5995 19945
<< pdcontact >>
rect 6245 19895 6295 19945
<< pdcontact >>
rect 7415 19895 7465 19945
<< pdcontact >>
rect 7715 19895 7765 19945
<< pdcontact >>
rect 8015 19895 8065 19945
<< pdcontact >>
rect 8315 19895 8365 19945
<< pdcontact >>
rect 8615 19895 8665 19945
<< pdcontact >>
rect 8915 19895 8965 19945
<< pdcontact >>
rect 9215 19895 9265 19945
<< pdcontact >>
rect 9515 19895 9565 19945
<< nsubstratencontact >>
rect 9815 19895 9865 19945
<< psubstratepcontact >>
rect 10535 19865 10585 19915
<< psubstratepcontact >>
rect 10685 19865 10735 19915
<< pdcontact >>
rect 1235 19745 1285 19795
<< pdcontact >>
rect 1535 19745 1585 19795
<< pdcontact >>
rect 1835 19745 1885 19795
<< pdcontact >>
rect 2135 19745 2185 19795
<< pdcontact >>
rect 2435 19745 2485 19795
<< pdcontact >>
rect 2735 19745 2785 19795
<< pdcontact >>
rect 3035 19745 3085 19795
<< pdcontact >>
rect 3335 19745 3385 19795
<< pdcontact >>
rect 4505 19745 4555 19795
<< pdcontact >>
rect 4805 19745 4855 19795
<< pdcontact >>
rect 5945 19745 5995 19795
<< pdcontact >>
rect 6245 19745 6295 19795
<< pdcontact >>
rect 7415 19745 7465 19795
<< pdcontact >>
rect 7715 19745 7765 19795
<< pdcontact >>
rect 8015 19745 8065 19795
<< pdcontact >>
rect 8315 19745 8365 19795
<< pdcontact >>
rect 8615 19745 8665 19795
<< pdcontact >>
rect 8915 19745 8965 19795
<< pdcontact >>
rect 9215 19745 9265 19795
<< pdcontact >>
rect 9515 19745 9565 19795
<< psubstratepcontact >>
rect 65 19625 115 19675
<< psubstratepcontact >>
rect 215 19625 265 19675
<< nsubstratencontact >>
rect 605 19595 655 19645
<< nsubstratencontact >>
rect 755 19595 805 19645
<< nsubstratencontact >>
rect 5315 19595 5365 19645
<< nsubstratencontact >>
rect 5465 19595 5515 19645
<< nsubstratencontact >>
rect 9995 19595 10045 19645
<< nsubstratencontact >>
rect 10145 19595 10195 19645
<< psubstratepcontact >>
rect 10535 19625 10585 19675
<< psubstratepcontact >>
rect 10685 19625 10735 19675
<< polycontact >>
rect 995 19505 1045 19555
<< polycontact >>
rect 5075 19505 5125 19555
<< polycontact >>
rect 5675 19505 5725 19555
<< polycontact >>
rect 9755 19505 9805 19555
<< nsubstratencontact >>
rect 605 19445 655 19495
<< nsubstratencontact >>
rect 755 19445 805 19495
<< pdcontact >>
rect 1265 19445 1315 19495
<< pdcontact >>
rect 1415 19445 1465 19495
<< pdcontact >>
rect 1565 19445 1615 19495
<< pdcontact >>
rect 1715 19445 1765 19495
<< pdcontact >>
rect 1865 19445 1915 19495
<< pdcontact >>
rect 2015 19445 2065 19495
<< pdcontact >>
rect 2165 19445 2215 19495
<< pdcontact >>
rect 2315 19445 2365 19495
<< pdcontact >>
rect 2465 19445 2515 19495
<< pdcontact >>
rect 2615 19445 2665 19495
<< pdcontact >>
rect 2765 19445 2815 19495
<< pdcontact >>
rect 2915 19445 2965 19495
<< pdcontact >>
rect 3065 19445 3115 19495
<< pdcontact >>
rect 3215 19445 3265 19495
<< pdcontact >>
rect 3365 19445 3415 19495
<< pdcontact >>
rect 3515 19445 3565 19495
<< pdcontact >>
rect 3665 19445 3715 19495
<< pdcontact >>
rect 3815 19445 3865 19495
<< pdcontact >>
rect 3965 19445 4015 19495
<< pdcontact >>
rect 4115 19445 4165 19495
<< pdcontact >>
rect 4265 19445 4315 19495
<< pdcontact >>
rect 4415 19445 4465 19495
<< pdcontact >>
rect 4565 19445 4615 19495
<< pdcontact >>
rect 4715 19445 4765 19495
<< pdcontact >>
rect 4865 19445 4915 19495
<< nsubstratencontact >>
rect 5315 19445 5365 19495
<< nsubstratencontact >>
rect 5465 19445 5515 19495
<< pdcontact >>
rect 5885 19445 5935 19495
<< pdcontact >>
rect 6035 19445 6085 19495
<< pdcontact >>
rect 6185 19445 6235 19495
<< pdcontact >>
rect 6335 19445 6385 19495
<< pdcontact >>
rect 6485 19445 6535 19495
<< pdcontact >>
rect 6635 19445 6685 19495
<< pdcontact >>
rect 6785 19445 6835 19495
<< pdcontact >>
rect 6935 19445 6985 19495
<< pdcontact >>
rect 7085 19445 7135 19495
<< pdcontact >>
rect 7235 19445 7285 19495
<< pdcontact >>
rect 7385 19445 7435 19495
<< pdcontact >>
rect 7535 19445 7585 19495
<< pdcontact >>
rect 7685 19445 7735 19495
<< pdcontact >>
rect 7835 19445 7885 19495
<< pdcontact >>
rect 7985 19445 8035 19495
<< pdcontact >>
rect 8135 19445 8185 19495
<< pdcontact >>
rect 8285 19445 8335 19495
<< pdcontact >>
rect 8435 19445 8485 19495
<< pdcontact >>
rect 8585 19445 8635 19495
<< pdcontact >>
rect 8735 19445 8785 19495
<< pdcontact >>
rect 8885 19445 8935 19495
<< pdcontact >>
rect 9035 19445 9085 19495
<< pdcontact >>
rect 9185 19445 9235 19495
<< pdcontact >>
rect 9335 19445 9385 19495
<< pdcontact >>
rect 9485 19445 9535 19495
<< nsubstratencontact >>
rect 9995 19445 10045 19495
<< nsubstratencontact >>
rect 10145 19445 10195 19495
<< psubstratepcontact >>
rect 65 19385 115 19435
<< psubstratepcontact >>
rect 215 19385 265 19435
<< polycontact >>
rect 995 19355 1045 19405
<< polycontact >>
rect 5075 19355 5125 19405
<< polycontact >>
rect 5675 19355 5725 19405
<< polycontact >>
rect 9755 19355 9805 19405
<< psubstratepcontact >>
rect 10535 19385 10585 19435
<< psubstratepcontact >>
rect 10685 19385 10735 19435
<< nsubstratencontact >>
rect 605 19295 655 19345
<< nsubstratencontact >>
rect 755 19295 805 19345
<< pdcontact >>
rect 1265 19295 1315 19345
<< pdcontact >>
rect 1415 19295 1465 19345
<< pdcontact >>
rect 1565 19295 1615 19345
<< pdcontact >>
rect 1715 19295 1765 19345
<< pdcontact >>
rect 1865 19295 1915 19345
<< pdcontact >>
rect 2015 19295 2065 19345
<< pdcontact >>
rect 2165 19295 2215 19345
<< pdcontact >>
rect 2315 19295 2365 19345
<< pdcontact >>
rect 2465 19295 2515 19345
<< pdcontact >>
rect 2615 19295 2665 19345
<< pdcontact >>
rect 2765 19295 2815 19345
<< pdcontact >>
rect 2915 19295 2965 19345
<< pdcontact >>
rect 3065 19295 3115 19345
<< pdcontact >>
rect 3215 19295 3265 19345
<< pdcontact >>
rect 3365 19295 3415 19345
<< pdcontact >>
rect 3515 19295 3565 19345
<< pdcontact >>
rect 3665 19295 3715 19345
<< pdcontact >>
rect 3815 19295 3865 19345
<< pdcontact >>
rect 3965 19295 4015 19345
<< pdcontact >>
rect 4115 19295 4165 19345
<< pdcontact >>
rect 4265 19295 4315 19345
<< pdcontact >>
rect 4415 19295 4465 19345
<< pdcontact >>
rect 4565 19295 4615 19345
<< pdcontact >>
rect 4715 19295 4765 19345
<< pdcontact >>
rect 4865 19295 4915 19345
<< nsubstratencontact >>
rect 5315 19295 5365 19345
<< nsubstratencontact >>
rect 5465 19295 5515 19345
<< pdcontact >>
rect 5885 19295 5935 19345
<< pdcontact >>
rect 6035 19295 6085 19345
<< pdcontact >>
rect 6185 19295 6235 19345
<< pdcontact >>
rect 6335 19295 6385 19345
<< pdcontact >>
rect 6485 19295 6535 19345
<< pdcontact >>
rect 6635 19295 6685 19345
<< pdcontact >>
rect 6785 19295 6835 19345
<< pdcontact >>
rect 6935 19295 6985 19345
<< pdcontact >>
rect 7085 19295 7135 19345
<< pdcontact >>
rect 7235 19295 7285 19345
<< pdcontact >>
rect 7385 19295 7435 19345
<< pdcontact >>
rect 7535 19295 7585 19345
<< pdcontact >>
rect 7685 19295 7735 19345
<< pdcontact >>
rect 7835 19295 7885 19345
<< pdcontact >>
rect 7985 19295 8035 19345
<< pdcontact >>
rect 8135 19295 8185 19345
<< pdcontact >>
rect 8285 19295 8335 19345
<< pdcontact >>
rect 8435 19295 8485 19345
<< pdcontact >>
rect 8585 19295 8635 19345
<< pdcontact >>
rect 8735 19295 8785 19345
<< pdcontact >>
rect 8885 19295 8935 19345
<< pdcontact >>
rect 9035 19295 9085 19345
<< pdcontact >>
rect 9185 19295 9235 19345
<< pdcontact >>
rect 9335 19295 9385 19345
<< pdcontact >>
rect 9485 19295 9535 19345
<< nsubstratencontact >>
rect 9995 19295 10045 19345
<< nsubstratencontact >>
rect 10145 19295 10195 19345
<< polycontact >>
rect 995 19205 1045 19255
<< polycontact >>
rect 5075 19205 5125 19255
<< polycontact >>
rect 5675 19205 5725 19255
<< polycontact >>
rect 9755 19205 9805 19255
<< psubstratepcontact >>
rect 65 19145 115 19195
<< psubstratepcontact >>
rect 215 19145 265 19195
<< nsubstratencontact >>
rect 605 19145 655 19195
<< nsubstratencontact >>
rect 755 19145 805 19195
<< pdcontact >>
rect 1265 19145 1315 19195
<< pdcontact >>
rect 1415 19145 1465 19195
<< pdcontact >>
rect 1565 19145 1615 19195
<< pdcontact >>
rect 1715 19145 1765 19195
<< pdcontact >>
rect 1865 19145 1915 19195
<< pdcontact >>
rect 2015 19145 2065 19195
<< pdcontact >>
rect 2165 19145 2215 19195
<< pdcontact >>
rect 2315 19145 2365 19195
<< pdcontact >>
rect 2465 19145 2515 19195
<< pdcontact >>
rect 2615 19145 2665 19195
<< pdcontact >>
rect 2765 19145 2815 19195
<< pdcontact >>
rect 2915 19145 2965 19195
<< pdcontact >>
rect 3065 19145 3115 19195
<< pdcontact >>
rect 3215 19145 3265 19195
<< pdcontact >>
rect 3365 19145 3415 19195
<< pdcontact >>
rect 3515 19145 3565 19195
<< pdcontact >>
rect 3665 19145 3715 19195
<< pdcontact >>
rect 3815 19145 3865 19195
<< pdcontact >>
rect 3965 19145 4015 19195
<< pdcontact >>
rect 4115 19145 4165 19195
<< pdcontact >>
rect 4265 19145 4315 19195
<< pdcontact >>
rect 4415 19145 4465 19195
<< pdcontact >>
rect 4565 19145 4615 19195
<< pdcontact >>
rect 4715 19145 4765 19195
<< pdcontact >>
rect 4865 19145 4915 19195
<< nsubstratencontact >>
rect 5315 19145 5365 19195
<< nsubstratencontact >>
rect 5465 19145 5515 19195
<< pdcontact >>
rect 5885 19145 5935 19195
<< pdcontact >>
rect 6035 19145 6085 19195
<< pdcontact >>
rect 6185 19145 6235 19195
<< pdcontact >>
rect 6335 19145 6385 19195
<< pdcontact >>
rect 6485 19145 6535 19195
<< pdcontact >>
rect 6635 19145 6685 19195
<< pdcontact >>
rect 6785 19145 6835 19195
<< pdcontact >>
rect 6935 19145 6985 19195
<< pdcontact >>
rect 7085 19145 7135 19195
<< pdcontact >>
rect 7235 19145 7285 19195
<< pdcontact >>
rect 7385 19145 7435 19195
<< pdcontact >>
rect 7535 19145 7585 19195
<< pdcontact >>
rect 7685 19145 7735 19195
<< pdcontact >>
rect 7835 19145 7885 19195
<< pdcontact >>
rect 7985 19145 8035 19195
<< pdcontact >>
rect 8135 19145 8185 19195
<< pdcontact >>
rect 8285 19145 8335 19195
<< pdcontact >>
rect 8435 19145 8485 19195
<< pdcontact >>
rect 8585 19145 8635 19195
<< pdcontact >>
rect 8735 19145 8785 19195
<< pdcontact >>
rect 8885 19145 8935 19195
<< pdcontact >>
rect 9035 19145 9085 19195
<< pdcontact >>
rect 9185 19145 9235 19195
<< pdcontact >>
rect 9335 19145 9385 19195
<< pdcontact >>
rect 9485 19145 9535 19195
<< nsubstratencontact >>
rect 9995 19145 10045 19195
<< nsubstratencontact >>
rect 10145 19145 10195 19195
<< psubstratepcontact >>
rect 10535 19145 10585 19195
<< psubstratepcontact >>
rect 10685 19145 10735 19195
<< polycontact >>
rect 995 19055 1045 19105
<< polycontact >>
rect 5075 19055 5125 19105
<< polycontact >>
rect 5675 19055 5725 19105
<< polycontact >>
rect 9755 19055 9805 19105
<< nsubstratencontact >>
rect 605 18995 655 19045
<< nsubstratencontact >>
rect 755 18995 805 19045
<< pdcontact >>
rect 1265 18995 1315 19045
<< pdcontact >>
rect 1415 18995 1465 19045
<< pdcontact >>
rect 1565 18995 1615 19045
<< pdcontact >>
rect 1715 18995 1765 19045
<< pdcontact >>
rect 1865 18995 1915 19045
<< pdcontact >>
rect 2015 18995 2065 19045
<< pdcontact >>
rect 2165 18995 2215 19045
<< pdcontact >>
rect 2315 18995 2365 19045
<< pdcontact >>
rect 2465 18995 2515 19045
<< pdcontact >>
rect 2615 18995 2665 19045
<< pdcontact >>
rect 2765 18995 2815 19045
<< pdcontact >>
rect 2915 18995 2965 19045
<< pdcontact >>
rect 3065 18995 3115 19045
<< pdcontact >>
rect 3215 18995 3265 19045
<< pdcontact >>
rect 3365 18995 3415 19045
<< pdcontact >>
rect 3515 18995 3565 19045
<< pdcontact >>
rect 3665 18995 3715 19045
<< pdcontact >>
rect 3815 18995 3865 19045
<< pdcontact >>
rect 3965 18995 4015 19045
<< pdcontact >>
rect 4115 18995 4165 19045
<< pdcontact >>
rect 4265 18995 4315 19045
<< pdcontact >>
rect 4415 18995 4465 19045
<< pdcontact >>
rect 4565 18995 4615 19045
<< pdcontact >>
rect 4715 18995 4765 19045
<< pdcontact >>
rect 4865 18995 4915 19045
<< nsubstratencontact >>
rect 5315 18995 5365 19045
<< nsubstratencontact >>
rect 5465 18995 5515 19045
<< pdcontact >>
rect 5885 18995 5935 19045
<< pdcontact >>
rect 6035 18995 6085 19045
<< pdcontact >>
rect 6185 18995 6235 19045
<< pdcontact >>
rect 6335 18995 6385 19045
<< pdcontact >>
rect 6485 18995 6535 19045
<< pdcontact >>
rect 6635 18995 6685 19045
<< pdcontact >>
rect 6785 18995 6835 19045
<< pdcontact >>
rect 6935 18995 6985 19045
<< pdcontact >>
rect 7085 18995 7135 19045
<< pdcontact >>
rect 7235 18995 7285 19045
<< pdcontact >>
rect 7385 18995 7435 19045
<< pdcontact >>
rect 7535 18995 7585 19045
<< pdcontact >>
rect 7685 18995 7735 19045
<< pdcontact >>
rect 7835 18995 7885 19045
<< pdcontact >>
rect 7985 18995 8035 19045
<< pdcontact >>
rect 8135 18995 8185 19045
<< pdcontact >>
rect 8285 18995 8335 19045
<< pdcontact >>
rect 8435 18995 8485 19045
<< pdcontact >>
rect 8585 18995 8635 19045
<< pdcontact >>
rect 8735 18995 8785 19045
<< pdcontact >>
rect 8885 18995 8935 19045
<< pdcontact >>
rect 9035 18995 9085 19045
<< pdcontact >>
rect 9185 18995 9235 19045
<< pdcontact >>
rect 9335 18995 9385 19045
<< pdcontact >>
rect 9485 18995 9535 19045
<< nsubstratencontact >>
rect 9995 18995 10045 19045
<< nsubstratencontact >>
rect 10145 18995 10195 19045
<< psubstratepcontact >>
rect 65 18905 115 18955
<< psubstratepcontact >>
rect 215 18905 265 18955
<< polycontact >>
rect 995 18905 1045 18955
<< polycontact >>
rect 5075 18905 5125 18955
<< polycontact >>
rect 5675 18905 5725 18955
<< polycontact >>
rect 9755 18905 9805 18955
<< psubstratepcontact >>
rect 10535 18905 10585 18955
<< psubstratepcontact >>
rect 10685 18905 10735 18955
<< nsubstratencontact >>
rect 605 18845 655 18895
<< nsubstratencontact >>
rect 755 18845 805 18895
<< pdcontact >>
rect 1265 18845 1315 18895
<< pdcontact >>
rect 1415 18845 1465 18895
<< pdcontact >>
rect 1565 18845 1615 18895
<< pdcontact >>
rect 1715 18845 1765 18895
<< pdcontact >>
rect 1865 18845 1915 18895
<< pdcontact >>
rect 2015 18845 2065 18895
<< pdcontact >>
rect 2165 18845 2215 18895
<< pdcontact >>
rect 2315 18845 2365 18895
<< pdcontact >>
rect 2465 18845 2515 18895
<< pdcontact >>
rect 2615 18845 2665 18895
<< pdcontact >>
rect 2765 18845 2815 18895
<< pdcontact >>
rect 2915 18845 2965 18895
<< pdcontact >>
rect 3065 18845 3115 18895
<< pdcontact >>
rect 3215 18845 3265 18895
<< pdcontact >>
rect 3365 18845 3415 18895
<< pdcontact >>
rect 3515 18845 3565 18895
<< pdcontact >>
rect 3665 18845 3715 18895
<< pdcontact >>
rect 3815 18845 3865 18895
<< pdcontact >>
rect 3965 18845 4015 18895
<< pdcontact >>
rect 4115 18845 4165 18895
<< pdcontact >>
rect 4265 18845 4315 18895
<< pdcontact >>
rect 4415 18845 4465 18895
<< pdcontact >>
rect 4565 18845 4615 18895
<< pdcontact >>
rect 4715 18845 4765 18895
<< pdcontact >>
rect 4865 18845 4915 18895
<< nsubstratencontact >>
rect 5315 18845 5365 18895
<< nsubstratencontact >>
rect 5465 18845 5515 18895
<< pdcontact >>
rect 5885 18845 5935 18895
<< pdcontact >>
rect 6035 18845 6085 18895
<< pdcontact >>
rect 6185 18845 6235 18895
<< pdcontact >>
rect 6335 18845 6385 18895
<< pdcontact >>
rect 6485 18845 6535 18895
<< pdcontact >>
rect 6635 18845 6685 18895
<< pdcontact >>
rect 6785 18845 6835 18895
<< pdcontact >>
rect 6935 18845 6985 18895
<< pdcontact >>
rect 7085 18845 7135 18895
<< pdcontact >>
rect 7235 18845 7285 18895
<< pdcontact >>
rect 7385 18845 7435 18895
<< pdcontact >>
rect 7535 18845 7585 18895
<< pdcontact >>
rect 7685 18845 7735 18895
<< pdcontact >>
rect 7835 18845 7885 18895
<< pdcontact >>
rect 7985 18845 8035 18895
<< pdcontact >>
rect 8135 18845 8185 18895
<< pdcontact >>
rect 8285 18845 8335 18895
<< pdcontact >>
rect 8435 18845 8485 18895
<< pdcontact >>
rect 8585 18845 8635 18895
<< pdcontact >>
rect 8735 18845 8785 18895
<< pdcontact >>
rect 8885 18845 8935 18895
<< pdcontact >>
rect 9035 18845 9085 18895
<< pdcontact >>
rect 9185 18845 9235 18895
<< pdcontact >>
rect 9335 18845 9385 18895
<< pdcontact >>
rect 9485 18845 9535 18895
<< nsubstratencontact >>
rect 9995 18845 10045 18895
<< nsubstratencontact >>
rect 10145 18845 10195 18895
<< polycontact >>
rect 995 18755 1045 18805
<< polycontact >>
rect 5075 18755 5125 18805
<< polycontact >>
rect 5675 18755 5725 18805
<< polycontact >>
rect 9755 18755 9805 18805
<< psubstratepcontact >>
rect 65 18665 115 18715
<< psubstratepcontact >>
rect 215 18665 265 18715
<< nsubstratencontact >>
rect 605 18695 655 18745
<< nsubstratencontact >>
rect 755 18695 805 18745
<< pdcontact >>
rect 1265 18695 1315 18745
<< pdcontact >>
rect 1415 18695 1465 18745
<< pdcontact >>
rect 1565 18695 1615 18745
<< pdcontact >>
rect 1715 18695 1765 18745
<< pdcontact >>
rect 1865 18695 1915 18745
<< pdcontact >>
rect 2015 18695 2065 18745
<< pdcontact >>
rect 2165 18695 2215 18745
<< pdcontact >>
rect 2315 18695 2365 18745
<< pdcontact >>
rect 2465 18695 2515 18745
<< pdcontact >>
rect 2615 18695 2665 18745
<< pdcontact >>
rect 2765 18695 2815 18745
<< pdcontact >>
rect 2915 18695 2965 18745
<< pdcontact >>
rect 3065 18695 3115 18745
<< pdcontact >>
rect 3215 18695 3265 18745
<< pdcontact >>
rect 3365 18695 3415 18745
<< pdcontact >>
rect 3515 18695 3565 18745
<< pdcontact >>
rect 3665 18695 3715 18745
<< pdcontact >>
rect 3815 18695 3865 18745
<< pdcontact >>
rect 3965 18695 4015 18745
<< pdcontact >>
rect 4115 18695 4165 18745
<< pdcontact >>
rect 4265 18695 4315 18745
<< pdcontact >>
rect 4415 18695 4465 18745
<< pdcontact >>
rect 4565 18695 4615 18745
<< pdcontact >>
rect 4715 18695 4765 18745
<< pdcontact >>
rect 4865 18695 4915 18745
<< nsubstratencontact >>
rect 5315 18695 5365 18745
<< nsubstratencontact >>
rect 5465 18695 5515 18745
<< pdcontact >>
rect 5885 18695 5935 18745
<< pdcontact >>
rect 6035 18695 6085 18745
<< pdcontact >>
rect 6185 18695 6235 18745
<< pdcontact >>
rect 6335 18695 6385 18745
<< pdcontact >>
rect 6485 18695 6535 18745
<< pdcontact >>
rect 6635 18695 6685 18745
<< pdcontact >>
rect 6785 18695 6835 18745
<< pdcontact >>
rect 6935 18695 6985 18745
<< pdcontact >>
rect 7085 18695 7135 18745
<< pdcontact >>
rect 7235 18695 7285 18745
<< pdcontact >>
rect 7385 18695 7435 18745
<< pdcontact >>
rect 7535 18695 7585 18745
<< pdcontact >>
rect 7685 18695 7735 18745
<< pdcontact >>
rect 7835 18695 7885 18745
<< pdcontact >>
rect 7985 18695 8035 18745
<< pdcontact >>
rect 8135 18695 8185 18745
<< pdcontact >>
rect 8285 18695 8335 18745
<< pdcontact >>
rect 8435 18695 8485 18745
<< pdcontact >>
rect 8585 18695 8635 18745
<< pdcontact >>
rect 8735 18695 8785 18745
<< pdcontact >>
rect 8885 18695 8935 18745
<< pdcontact >>
rect 9035 18695 9085 18745
<< pdcontact >>
rect 9185 18695 9235 18745
<< pdcontact >>
rect 9335 18695 9385 18745
<< pdcontact >>
rect 9485 18695 9535 18745
<< nsubstratencontact >>
rect 9995 18695 10045 18745
<< nsubstratencontact >>
rect 10145 18695 10195 18745
<< psubstratepcontact >>
rect 10535 18665 10585 18715
<< psubstratepcontact >>
rect 10685 18665 10735 18715
<< polycontact >>
rect 995 18605 1045 18655
<< polycontact >>
rect 5075 18605 5125 18655
<< polycontact >>
rect 5675 18605 5725 18655
<< polycontact >>
rect 9755 18605 9805 18655
<< nsubstratencontact >>
rect 605 18545 655 18595
<< nsubstratencontact >>
rect 755 18545 805 18595
<< pdcontact >>
rect 1265 18545 1315 18595
<< pdcontact >>
rect 1415 18545 1465 18595
<< pdcontact >>
rect 1565 18545 1615 18595
<< pdcontact >>
rect 1715 18545 1765 18595
<< pdcontact >>
rect 1865 18545 1915 18595
<< pdcontact >>
rect 2015 18545 2065 18595
<< pdcontact >>
rect 2165 18545 2215 18595
<< pdcontact >>
rect 2315 18545 2365 18595
<< pdcontact >>
rect 2465 18545 2515 18595
<< pdcontact >>
rect 2615 18545 2665 18595
<< pdcontact >>
rect 2765 18545 2815 18595
<< pdcontact >>
rect 2915 18545 2965 18595
<< pdcontact >>
rect 3065 18545 3115 18595
<< pdcontact >>
rect 3215 18545 3265 18595
<< pdcontact >>
rect 3365 18545 3415 18595
<< pdcontact >>
rect 3515 18545 3565 18595
<< pdcontact >>
rect 3665 18545 3715 18595
<< pdcontact >>
rect 3815 18545 3865 18595
<< pdcontact >>
rect 3965 18545 4015 18595
<< pdcontact >>
rect 4115 18545 4165 18595
<< pdcontact >>
rect 4265 18545 4315 18595
<< pdcontact >>
rect 4415 18545 4465 18595
<< pdcontact >>
rect 4565 18545 4615 18595
<< pdcontact >>
rect 4715 18545 4765 18595
<< pdcontact >>
rect 4865 18545 4915 18595
<< nsubstratencontact >>
rect 5315 18545 5365 18595
<< nsubstratencontact >>
rect 5465 18545 5515 18595
<< pdcontact >>
rect 5885 18545 5935 18595
<< pdcontact >>
rect 6035 18545 6085 18595
<< pdcontact >>
rect 6185 18545 6235 18595
<< pdcontact >>
rect 6335 18545 6385 18595
<< pdcontact >>
rect 6485 18545 6535 18595
<< pdcontact >>
rect 6635 18545 6685 18595
<< pdcontact >>
rect 6785 18545 6835 18595
<< pdcontact >>
rect 6935 18545 6985 18595
<< pdcontact >>
rect 7085 18545 7135 18595
<< pdcontact >>
rect 7235 18545 7285 18595
<< pdcontact >>
rect 7385 18545 7435 18595
<< pdcontact >>
rect 7535 18545 7585 18595
<< pdcontact >>
rect 7685 18545 7735 18595
<< pdcontact >>
rect 7835 18545 7885 18595
<< pdcontact >>
rect 7985 18545 8035 18595
<< pdcontact >>
rect 8135 18545 8185 18595
<< pdcontact >>
rect 8285 18545 8335 18595
<< pdcontact >>
rect 8435 18545 8485 18595
<< pdcontact >>
rect 8585 18545 8635 18595
<< pdcontact >>
rect 8735 18545 8785 18595
<< pdcontact >>
rect 8885 18545 8935 18595
<< pdcontact >>
rect 9035 18545 9085 18595
<< pdcontact >>
rect 9185 18545 9235 18595
<< pdcontact >>
rect 9335 18545 9385 18595
<< pdcontact >>
rect 9485 18545 9535 18595
<< nsubstratencontact >>
rect 9995 18545 10045 18595
<< nsubstratencontact >>
rect 10145 18545 10195 18595
<< psubstratepcontact >>
rect 65 18425 115 18475
<< psubstratepcontact >>
rect 215 18425 265 18475
<< polycontact >>
rect 995 18455 1045 18505
<< polycontact >>
rect 5075 18455 5125 18505
<< polycontact >>
rect 5675 18455 5725 18505
<< polycontact >>
rect 9755 18455 9805 18505
<< nsubstratencontact >>
rect 605 18395 655 18445
<< nsubstratencontact >>
rect 755 18395 805 18445
<< pdcontact >>
rect 1265 18395 1315 18445
<< pdcontact >>
rect 1415 18395 1465 18445
<< pdcontact >>
rect 1565 18395 1615 18445
<< pdcontact >>
rect 1715 18395 1765 18445
<< pdcontact >>
rect 1865 18395 1915 18445
<< pdcontact >>
rect 2015 18395 2065 18445
<< pdcontact >>
rect 2165 18395 2215 18445
<< pdcontact >>
rect 2315 18395 2365 18445
<< pdcontact >>
rect 2465 18395 2515 18445
<< pdcontact >>
rect 2615 18395 2665 18445
<< pdcontact >>
rect 2765 18395 2815 18445
<< pdcontact >>
rect 2915 18395 2965 18445
<< pdcontact >>
rect 3065 18395 3115 18445
<< pdcontact >>
rect 3215 18395 3265 18445
<< pdcontact >>
rect 3365 18395 3415 18445
<< pdcontact >>
rect 3515 18395 3565 18445
<< pdcontact >>
rect 3665 18395 3715 18445
<< pdcontact >>
rect 3815 18395 3865 18445
<< pdcontact >>
rect 3965 18395 4015 18445
<< pdcontact >>
rect 4115 18395 4165 18445
<< pdcontact >>
rect 4265 18395 4315 18445
<< pdcontact >>
rect 4415 18395 4465 18445
<< pdcontact >>
rect 4565 18395 4615 18445
<< pdcontact >>
rect 4715 18395 4765 18445
<< pdcontact >>
rect 4865 18395 4915 18445
<< nsubstratencontact >>
rect 5315 18395 5365 18445
<< nsubstratencontact >>
rect 5465 18395 5515 18445
<< pdcontact >>
rect 5885 18395 5935 18445
<< pdcontact >>
rect 6035 18395 6085 18445
<< pdcontact >>
rect 6185 18395 6235 18445
<< pdcontact >>
rect 6335 18395 6385 18445
<< pdcontact >>
rect 6485 18395 6535 18445
<< pdcontact >>
rect 6635 18395 6685 18445
<< pdcontact >>
rect 6785 18395 6835 18445
<< pdcontact >>
rect 6935 18395 6985 18445
<< pdcontact >>
rect 7085 18395 7135 18445
<< pdcontact >>
rect 7235 18395 7285 18445
<< pdcontact >>
rect 7385 18395 7435 18445
<< pdcontact >>
rect 7535 18395 7585 18445
<< pdcontact >>
rect 7685 18395 7735 18445
<< pdcontact >>
rect 7835 18395 7885 18445
<< pdcontact >>
rect 7985 18395 8035 18445
<< pdcontact >>
rect 8135 18395 8185 18445
<< pdcontact >>
rect 8285 18395 8335 18445
<< pdcontact >>
rect 8435 18395 8485 18445
<< pdcontact >>
rect 8585 18395 8635 18445
<< pdcontact >>
rect 8735 18395 8785 18445
<< pdcontact >>
rect 8885 18395 8935 18445
<< pdcontact >>
rect 9035 18395 9085 18445
<< pdcontact >>
rect 9185 18395 9235 18445
<< pdcontact >>
rect 9335 18395 9385 18445
<< pdcontact >>
rect 9485 18395 9535 18445
<< nsubstratencontact >>
rect 9995 18395 10045 18445
<< nsubstratencontact >>
rect 10145 18395 10195 18445
<< psubstratepcontact >>
rect 10535 18425 10585 18475
<< psubstratepcontact >>
rect 10685 18425 10735 18475
<< polycontact >>
rect 995 18305 1045 18355
<< polycontact >>
rect 5075 18305 5125 18355
<< polycontact >>
rect 5675 18305 5725 18355
<< polycontact >>
rect 9755 18305 9805 18355
<< nsubstratencontact >>
rect 605 18245 655 18295
<< nsubstratencontact >>
rect 755 18245 805 18295
<< nsubstratencontact >>
rect 5315 18245 5365 18295
<< nsubstratencontact >>
rect 5465 18245 5515 18295
<< nsubstratencontact >>
rect 9995 18245 10045 18295
<< nsubstratencontact >>
rect 10145 18245 10195 18295
<< psubstratepcontact >>
rect 65 18185 115 18235
<< psubstratepcontact >>
rect 215 18185 265 18235
<< polycontact >>
rect 995 18155 1045 18205
<< polycontact >>
rect 5075 18155 5125 18205
<< polycontact >>
rect 5675 18155 5725 18205
<< polycontact >>
rect 9755 18155 9805 18205
<< psubstratepcontact >>
rect 10535 18185 10585 18235
<< psubstratepcontact >>
rect 10685 18185 10735 18235
<< pdcontact >>
rect 1235 18095 1285 18145
<< pdcontact >>
rect 1535 18095 1585 18145
<< pdcontact >>
rect 1835 18095 1885 18145
<< pdcontact >>
rect 2135 18095 2185 18145
<< pdcontact >>
rect 2435 18095 2485 18145
<< pdcontact >>
rect 2735 18095 2785 18145
<< pdcontact >>
rect 3035 18095 3085 18145
<< pdcontact >>
rect 3335 18095 3385 18145
<< pdcontact >>
rect 4505 18095 4555 18145
<< pdcontact >>
rect 4805 18095 4855 18145
<< pdcontact >>
rect 5945 18095 5995 18145
<< pdcontact >>
rect 6245 18095 6295 18145
<< pdcontact >>
rect 7415 18095 7465 18145
<< pdcontact >>
rect 7715 18095 7765 18145
<< pdcontact >>
rect 8015 18095 8065 18145
<< pdcontact >>
rect 8315 18095 8365 18145
<< pdcontact >>
rect 8615 18095 8665 18145
<< pdcontact >>
rect 8915 18095 8965 18145
<< pdcontact >>
rect 9215 18095 9265 18145
<< pdcontact >>
rect 9515 18095 9565 18145
<< polycontact >>
rect 995 18005 1045 18055
<< polycontact >>
rect 5075 18005 5125 18055
<< polycontact >>
rect 5675 18005 5725 18055
<< polycontact >>
rect 9755 18005 9805 18055
<< psubstratepcontact >>
rect 65 17945 115 17995
<< psubstratepcontact >>
rect 215 17945 265 17995
<< pdcontact >>
rect 1235 17945 1285 17995
<< pdcontact >>
rect 1535 17945 1585 17995
<< pdcontact >>
rect 1835 17945 1885 17995
<< pdcontact >>
rect 2135 17945 2185 17995
<< pdcontact >>
rect 2435 17945 2485 17995
<< pdcontact >>
rect 2735 17945 2785 17995
<< pdcontact >>
rect 3035 17945 3085 17995
<< pdcontact >>
rect 3335 17945 3385 17995
<< pdcontact >>
rect 4505 17945 4555 17995
<< pdcontact >>
rect 4805 17945 4855 17995
<< pdcontact >>
rect 5945 17945 5995 17995
<< pdcontact >>
rect 6245 17945 6295 17995
<< pdcontact >>
rect 7415 17945 7465 17995
<< pdcontact >>
rect 7715 17945 7765 17995
<< pdcontact >>
rect 8015 17945 8065 17995
<< pdcontact >>
rect 8315 17945 8365 17995
<< pdcontact >>
rect 8615 17945 8665 17995
<< pdcontact >>
rect 8915 17945 8965 17995
<< pdcontact >>
rect 9215 17945 9265 17995
<< pdcontact >>
rect 9515 17945 9565 17995
<< psubstratepcontact >>
rect 10535 17945 10585 17995
<< psubstratepcontact >>
rect 10685 17945 10735 17995
<< polycontact >>
rect 995 17855 1045 17905
<< polycontact >>
rect 5075 17855 5125 17905
<< polycontact >>
rect 5675 17855 5725 17905
<< polycontact >>
rect 9755 17855 9805 17905
<< pdcontact >>
rect 1235 17795 1285 17845
<< pdcontact >>
rect 1535 17795 1585 17845
<< pdcontact >>
rect 1835 17795 1885 17845
<< pdcontact >>
rect 2135 17795 2185 17845
<< pdcontact >>
rect 2435 17795 2485 17845
<< pdcontact >>
rect 2735 17795 2785 17845
<< pdcontact >>
rect 3035 17795 3085 17845
<< pdcontact >>
rect 3335 17795 3385 17845
<< pdcontact >>
rect 4505 17795 4555 17845
<< pdcontact >>
rect 4805 17795 4855 17845
<< pdcontact >>
rect 5945 17795 5995 17845
<< pdcontact >>
rect 6245 17795 6295 17845
<< pdcontact >>
rect 7415 17795 7465 17845
<< pdcontact >>
rect 7715 17795 7765 17845
<< pdcontact >>
rect 8015 17795 8065 17845
<< pdcontact >>
rect 8315 17795 8365 17845
<< pdcontact >>
rect 8615 17795 8665 17845
<< pdcontact >>
rect 8915 17795 8965 17845
<< pdcontact >>
rect 9215 17795 9265 17845
<< pdcontact >>
rect 9515 17795 9565 17845
<< psubstratepcontact >>
rect 65 17705 115 17755
<< psubstratepcontact >>
rect 215 17705 265 17755
<< polycontact >>
rect 995 17705 1045 17755
<< polycontact >>
rect 5075 17705 5125 17755
<< polycontact >>
rect 5675 17705 5725 17755
<< polycontact >>
rect 9755 17705 9805 17755
<< psubstratepcontact >>
rect 10535 17705 10585 17755
<< psubstratepcontact >>
rect 10685 17705 10735 17755
<< nsubstratencontact >>
rect 605 17645 655 17695
<< nsubstratencontact >>
rect 755 17645 805 17695
<< nsubstratencontact >>
rect 5315 17645 5365 17695
<< nsubstratencontact >>
rect 5465 17645 5515 17695
<< nsubstratencontact >>
rect 9995 17645 10045 17695
<< nsubstratencontact >>
rect 10145 17645 10195 17695
<< polycontact >>
rect 995 17555 1045 17605
<< polycontact >>
rect 5075 17555 5125 17605
<< polycontact >>
rect 5675 17555 5725 17605
<< polycontact >>
rect 9755 17555 9805 17605
<< psubstratepcontact >>
rect 65 17465 115 17515
<< psubstratepcontact >>
rect 215 17465 265 17515
<< nsubstratencontact >>
rect 605 17495 655 17545
<< nsubstratencontact >>
rect 755 17495 805 17545
<< pdcontact >>
rect 1265 17495 1315 17545
<< pdcontact >>
rect 1415 17495 1465 17545
<< pdcontact >>
rect 1565 17495 1615 17545
<< pdcontact >>
rect 1715 17495 1765 17545
<< pdcontact >>
rect 1865 17495 1915 17545
<< pdcontact >>
rect 2015 17495 2065 17545
<< pdcontact >>
rect 2165 17495 2215 17545
<< pdcontact >>
rect 2315 17495 2365 17545
<< pdcontact >>
rect 2465 17495 2515 17545
<< pdcontact >>
rect 2615 17495 2665 17545
<< pdcontact >>
rect 2765 17495 2815 17545
<< pdcontact >>
rect 2915 17495 2965 17545
<< pdcontact >>
rect 3065 17495 3115 17545
<< pdcontact >>
rect 3215 17495 3265 17545
<< pdcontact >>
rect 3365 17495 3415 17545
<< pdcontact >>
rect 3515 17495 3565 17545
<< pdcontact >>
rect 3665 17495 3715 17545
<< pdcontact >>
rect 3815 17495 3865 17545
<< pdcontact >>
rect 3965 17495 4015 17545
<< pdcontact >>
rect 4115 17495 4165 17545
<< pdcontact >>
rect 4265 17495 4315 17545
<< pdcontact >>
rect 4415 17495 4465 17545
<< pdcontact >>
rect 4565 17495 4615 17545
<< pdcontact >>
rect 4715 17495 4765 17545
<< pdcontact >>
rect 4865 17495 4915 17545
<< nsubstratencontact >>
rect 5315 17495 5365 17545
<< nsubstratencontact >>
rect 5465 17495 5515 17545
<< pdcontact >>
rect 5885 17495 5935 17545
<< pdcontact >>
rect 6035 17495 6085 17545
<< pdcontact >>
rect 6185 17495 6235 17545
<< pdcontact >>
rect 6335 17495 6385 17545
<< pdcontact >>
rect 6485 17495 6535 17545
<< pdcontact >>
rect 6635 17495 6685 17545
<< pdcontact >>
rect 6785 17495 6835 17545
<< pdcontact >>
rect 6935 17495 6985 17545
<< pdcontact >>
rect 7085 17495 7135 17545
<< pdcontact >>
rect 7235 17495 7285 17545
<< pdcontact >>
rect 7385 17495 7435 17545
<< pdcontact >>
rect 7535 17495 7585 17545
<< pdcontact >>
rect 7685 17495 7735 17545
<< pdcontact >>
rect 7835 17495 7885 17545
<< pdcontact >>
rect 7985 17495 8035 17545
<< pdcontact >>
rect 8135 17495 8185 17545
<< pdcontact >>
rect 8285 17495 8335 17545
<< pdcontact >>
rect 8435 17495 8485 17545
<< pdcontact >>
rect 8585 17495 8635 17545
<< pdcontact >>
rect 8735 17495 8785 17545
<< pdcontact >>
rect 8885 17495 8935 17545
<< pdcontact >>
rect 9035 17495 9085 17545
<< pdcontact >>
rect 9185 17495 9235 17545
<< pdcontact >>
rect 9335 17495 9385 17545
<< pdcontact >>
rect 9485 17495 9535 17545
<< nsubstratencontact >>
rect 9995 17495 10045 17545
<< nsubstratencontact >>
rect 10145 17495 10195 17545
<< psubstratepcontact >>
rect 10535 17465 10585 17515
<< psubstratepcontact >>
rect 10685 17465 10735 17515
<< polycontact >>
rect 995 17405 1045 17455
<< polycontact >>
rect 5075 17405 5125 17455
<< polycontact >>
rect 5675 17405 5725 17455
<< polycontact >>
rect 9755 17405 9805 17455
<< nsubstratencontact >>
rect 605 17345 655 17395
<< nsubstratencontact >>
rect 755 17345 805 17395
<< pdcontact >>
rect 1265 17345 1315 17395
<< pdcontact >>
rect 1415 17345 1465 17395
<< pdcontact >>
rect 1565 17345 1615 17395
<< pdcontact >>
rect 1715 17345 1765 17395
<< pdcontact >>
rect 1865 17345 1915 17395
<< pdcontact >>
rect 2015 17345 2065 17395
<< pdcontact >>
rect 2165 17345 2215 17395
<< pdcontact >>
rect 2315 17345 2365 17395
<< pdcontact >>
rect 2465 17345 2515 17395
<< pdcontact >>
rect 2615 17345 2665 17395
<< pdcontact >>
rect 2765 17345 2815 17395
<< pdcontact >>
rect 2915 17345 2965 17395
<< pdcontact >>
rect 3065 17345 3115 17395
<< pdcontact >>
rect 3215 17345 3265 17395
<< pdcontact >>
rect 3365 17345 3415 17395
<< pdcontact >>
rect 3515 17345 3565 17395
<< pdcontact >>
rect 3665 17345 3715 17395
<< pdcontact >>
rect 3815 17345 3865 17395
<< pdcontact >>
rect 3965 17345 4015 17395
<< pdcontact >>
rect 4115 17345 4165 17395
<< pdcontact >>
rect 4265 17345 4315 17395
<< pdcontact >>
rect 4415 17345 4465 17395
<< pdcontact >>
rect 4565 17345 4615 17395
<< pdcontact >>
rect 4715 17345 4765 17395
<< pdcontact >>
rect 4865 17345 4915 17395
<< nsubstratencontact >>
rect 5315 17345 5365 17395
<< nsubstratencontact >>
rect 5465 17345 5515 17395
<< pdcontact >>
rect 5885 17345 5935 17395
<< pdcontact >>
rect 6035 17345 6085 17395
<< pdcontact >>
rect 6185 17345 6235 17395
<< pdcontact >>
rect 6335 17345 6385 17395
<< pdcontact >>
rect 6485 17345 6535 17395
<< pdcontact >>
rect 6635 17345 6685 17395
<< pdcontact >>
rect 6785 17345 6835 17395
<< pdcontact >>
rect 6935 17345 6985 17395
<< pdcontact >>
rect 7085 17345 7135 17395
<< pdcontact >>
rect 7235 17345 7285 17395
<< pdcontact >>
rect 7385 17345 7435 17395
<< pdcontact >>
rect 7535 17345 7585 17395
<< pdcontact >>
rect 7685 17345 7735 17395
<< pdcontact >>
rect 7835 17345 7885 17395
<< pdcontact >>
rect 7985 17345 8035 17395
<< pdcontact >>
rect 8135 17345 8185 17395
<< pdcontact >>
rect 8285 17345 8335 17395
<< pdcontact >>
rect 8435 17345 8485 17395
<< pdcontact >>
rect 8585 17345 8635 17395
<< pdcontact >>
rect 8735 17345 8785 17395
<< pdcontact >>
rect 8885 17345 8935 17395
<< pdcontact >>
rect 9035 17345 9085 17395
<< pdcontact >>
rect 9185 17345 9235 17395
<< pdcontact >>
rect 9335 17345 9385 17395
<< pdcontact >>
rect 9485 17345 9535 17395
<< nsubstratencontact >>
rect 9995 17345 10045 17395
<< nsubstratencontact >>
rect 10145 17345 10195 17395
<< psubstratepcontact >>
rect 65 17225 115 17275
<< psubstratepcontact >>
rect 215 17225 265 17275
<< polycontact >>
rect 995 17255 1045 17305
<< polycontact >>
rect 5075 17255 5125 17305
<< polycontact >>
rect 5675 17255 5725 17305
<< polycontact >>
rect 9755 17255 9805 17305
<< nsubstratencontact >>
rect 605 17195 655 17245
<< nsubstratencontact >>
rect 755 17195 805 17245
<< pdcontact >>
rect 1265 17195 1315 17245
<< pdcontact >>
rect 1415 17195 1465 17245
<< pdcontact >>
rect 1565 17195 1615 17245
<< pdcontact >>
rect 1715 17195 1765 17245
<< pdcontact >>
rect 1865 17195 1915 17245
<< pdcontact >>
rect 2015 17195 2065 17245
<< pdcontact >>
rect 2165 17195 2215 17245
<< pdcontact >>
rect 2315 17195 2365 17245
<< pdcontact >>
rect 2465 17195 2515 17245
<< pdcontact >>
rect 2615 17195 2665 17245
<< pdcontact >>
rect 2765 17195 2815 17245
<< pdcontact >>
rect 2915 17195 2965 17245
<< pdcontact >>
rect 3065 17195 3115 17245
<< pdcontact >>
rect 3215 17195 3265 17245
<< pdcontact >>
rect 3365 17195 3415 17245
<< pdcontact >>
rect 3515 17195 3565 17245
<< pdcontact >>
rect 3665 17195 3715 17245
<< pdcontact >>
rect 3815 17195 3865 17245
<< pdcontact >>
rect 3965 17195 4015 17245
<< pdcontact >>
rect 4115 17195 4165 17245
<< pdcontact >>
rect 4265 17195 4315 17245
<< pdcontact >>
rect 4415 17195 4465 17245
<< pdcontact >>
rect 4565 17195 4615 17245
<< pdcontact >>
rect 4715 17195 4765 17245
<< pdcontact >>
rect 4865 17195 4915 17245
<< nsubstratencontact >>
rect 5315 17195 5365 17245
<< nsubstratencontact >>
rect 5465 17195 5515 17245
<< pdcontact >>
rect 5885 17195 5935 17245
<< pdcontact >>
rect 6035 17195 6085 17245
<< pdcontact >>
rect 6185 17195 6235 17245
<< pdcontact >>
rect 6335 17195 6385 17245
<< pdcontact >>
rect 6485 17195 6535 17245
<< pdcontact >>
rect 6635 17195 6685 17245
<< pdcontact >>
rect 6785 17195 6835 17245
<< pdcontact >>
rect 6935 17195 6985 17245
<< pdcontact >>
rect 7085 17195 7135 17245
<< pdcontact >>
rect 7235 17195 7285 17245
<< pdcontact >>
rect 7385 17195 7435 17245
<< pdcontact >>
rect 7535 17195 7585 17245
<< pdcontact >>
rect 7685 17195 7735 17245
<< pdcontact >>
rect 7835 17195 7885 17245
<< pdcontact >>
rect 7985 17195 8035 17245
<< pdcontact >>
rect 8135 17195 8185 17245
<< pdcontact >>
rect 8285 17195 8335 17245
<< pdcontact >>
rect 8435 17195 8485 17245
<< pdcontact >>
rect 8585 17195 8635 17245
<< pdcontact >>
rect 8735 17195 8785 17245
<< pdcontact >>
rect 8885 17195 8935 17245
<< pdcontact >>
rect 9035 17195 9085 17245
<< pdcontact >>
rect 9185 17195 9235 17245
<< pdcontact >>
rect 9335 17195 9385 17245
<< pdcontact >>
rect 9485 17195 9535 17245
<< nsubstratencontact >>
rect 9995 17195 10045 17245
<< nsubstratencontact >>
rect 10145 17195 10195 17245
<< psubstratepcontact >>
rect 10535 17225 10585 17275
<< psubstratepcontact >>
rect 10685 17225 10735 17275
<< polycontact >>
rect 995 17105 1045 17155
<< polycontact >>
rect 5075 17105 5125 17155
<< polycontact >>
rect 5675 17105 5725 17155
<< polycontact >>
rect 9755 17105 9805 17155
<< nsubstratencontact >>
rect 605 17045 655 17095
<< nsubstratencontact >>
rect 755 17045 805 17095
<< pdcontact >>
rect 1265 17045 1315 17095
<< pdcontact >>
rect 1415 17045 1465 17095
<< pdcontact >>
rect 1565 17045 1615 17095
<< pdcontact >>
rect 1715 17045 1765 17095
<< pdcontact >>
rect 1865 17045 1915 17095
<< pdcontact >>
rect 2015 17045 2065 17095
<< pdcontact >>
rect 2165 17045 2215 17095
<< pdcontact >>
rect 2315 17045 2365 17095
<< pdcontact >>
rect 2465 17045 2515 17095
<< pdcontact >>
rect 2615 17045 2665 17095
<< pdcontact >>
rect 2765 17045 2815 17095
<< pdcontact >>
rect 2915 17045 2965 17095
<< pdcontact >>
rect 3065 17045 3115 17095
<< pdcontact >>
rect 3215 17045 3265 17095
<< pdcontact >>
rect 3365 17045 3415 17095
<< pdcontact >>
rect 3515 17045 3565 17095
<< pdcontact >>
rect 3665 17045 3715 17095
<< pdcontact >>
rect 3815 17045 3865 17095
<< pdcontact >>
rect 3965 17045 4015 17095
<< pdcontact >>
rect 4115 17045 4165 17095
<< pdcontact >>
rect 4265 17045 4315 17095
<< pdcontact >>
rect 4415 17045 4465 17095
<< pdcontact >>
rect 4565 17045 4615 17095
<< pdcontact >>
rect 4715 17045 4765 17095
<< pdcontact >>
rect 4865 17045 4915 17095
<< nsubstratencontact >>
rect 5315 17045 5365 17095
<< nsubstratencontact >>
rect 5465 17045 5515 17095
<< pdcontact >>
rect 5885 17045 5935 17095
<< pdcontact >>
rect 6035 17045 6085 17095
<< pdcontact >>
rect 6185 17045 6235 17095
<< pdcontact >>
rect 6335 17045 6385 17095
<< pdcontact >>
rect 6485 17045 6535 17095
<< pdcontact >>
rect 6635 17045 6685 17095
<< pdcontact >>
rect 6785 17045 6835 17095
<< pdcontact >>
rect 6935 17045 6985 17095
<< pdcontact >>
rect 7085 17045 7135 17095
<< pdcontact >>
rect 7235 17045 7285 17095
<< pdcontact >>
rect 7385 17045 7435 17095
<< pdcontact >>
rect 7535 17045 7585 17095
<< pdcontact >>
rect 7685 17045 7735 17095
<< pdcontact >>
rect 7835 17045 7885 17095
<< pdcontact >>
rect 7985 17045 8035 17095
<< pdcontact >>
rect 8135 17045 8185 17095
<< pdcontact >>
rect 8285 17045 8335 17095
<< pdcontact >>
rect 8435 17045 8485 17095
<< pdcontact >>
rect 8585 17045 8635 17095
<< pdcontact >>
rect 8735 17045 8785 17095
<< pdcontact >>
rect 8885 17045 8935 17095
<< pdcontact >>
rect 9035 17045 9085 17095
<< pdcontact >>
rect 9185 17045 9235 17095
<< pdcontact >>
rect 9335 17045 9385 17095
<< pdcontact >>
rect 9485 17045 9535 17095
<< nsubstratencontact >>
rect 9995 17045 10045 17095
<< nsubstratencontact >>
rect 10145 17045 10195 17095
<< psubstratepcontact >>
rect 65 16985 115 17035
<< psubstratepcontact >>
rect 215 16985 265 17035
<< psubstratepcontact >>
rect 10535 16985 10585 17035
<< psubstratepcontact >>
rect 10685 16985 10735 17035
<< nsubstratencontact >>
rect 605 16895 655 16945
<< nsubstratencontact >>
rect 755 16895 805 16945
<< polycontact >>
rect 995 16925 1045 16975
<< pdcontact >>
rect 1265 16895 1315 16945
<< pdcontact >>
rect 1415 16895 1465 16945
<< pdcontact >>
rect 1565 16895 1615 16945
<< pdcontact >>
rect 1715 16895 1765 16945
<< pdcontact >>
rect 1865 16895 1915 16945
<< pdcontact >>
rect 2015 16895 2065 16945
<< pdcontact >>
rect 2165 16895 2215 16945
<< pdcontact >>
rect 2315 16895 2365 16945
<< pdcontact >>
rect 2465 16895 2515 16945
<< pdcontact >>
rect 2615 16895 2665 16945
<< pdcontact >>
rect 2765 16895 2815 16945
<< pdcontact >>
rect 2915 16895 2965 16945
<< pdcontact >>
rect 3065 16895 3115 16945
<< pdcontact >>
rect 3215 16895 3265 16945
<< pdcontact >>
rect 3365 16895 3415 16945
<< pdcontact >>
rect 3515 16895 3565 16945
<< pdcontact >>
rect 3665 16895 3715 16945
<< pdcontact >>
rect 3815 16895 3865 16945
<< pdcontact >>
rect 3965 16895 4015 16945
<< pdcontact >>
rect 4115 16895 4165 16945
<< pdcontact >>
rect 4265 16895 4315 16945
<< pdcontact >>
rect 4415 16895 4465 16945
<< pdcontact >>
rect 4565 16895 4615 16945
<< pdcontact >>
rect 4715 16895 4765 16945
<< pdcontact >>
rect 4865 16895 4915 16945
<< polycontact >>
rect 5075 16925 5125 16975
<< nsubstratencontact >>
rect 5315 16895 5365 16945
<< nsubstratencontact >>
rect 5465 16895 5515 16945
<< polycontact >>
rect 5675 16925 5725 16975
<< pdcontact >>
rect 5885 16895 5935 16945
<< pdcontact >>
rect 6035 16895 6085 16945
<< pdcontact >>
rect 6185 16895 6235 16945
<< pdcontact >>
rect 6335 16895 6385 16945
<< pdcontact >>
rect 6485 16895 6535 16945
<< pdcontact >>
rect 6635 16895 6685 16945
<< pdcontact >>
rect 6785 16895 6835 16945
<< pdcontact >>
rect 6935 16895 6985 16945
<< pdcontact >>
rect 7085 16895 7135 16945
<< pdcontact >>
rect 7235 16895 7285 16945
<< pdcontact >>
rect 7385 16895 7435 16945
<< pdcontact >>
rect 7535 16895 7585 16945
<< pdcontact >>
rect 7685 16895 7735 16945
<< pdcontact >>
rect 7835 16895 7885 16945
<< pdcontact >>
rect 7985 16895 8035 16945
<< pdcontact >>
rect 8135 16895 8185 16945
<< pdcontact >>
rect 8285 16895 8335 16945
<< pdcontact >>
rect 8435 16895 8485 16945
<< pdcontact >>
rect 8585 16895 8635 16945
<< pdcontact >>
rect 8735 16895 8785 16945
<< pdcontact >>
rect 8885 16895 8935 16945
<< pdcontact >>
rect 9035 16895 9085 16945
<< pdcontact >>
rect 9185 16895 9235 16945
<< pdcontact >>
rect 9335 16895 9385 16945
<< pdcontact >>
rect 9485 16895 9535 16945
<< polycontact >>
rect 9755 16925 9805 16975
<< nsubstratencontact >>
rect 9995 16895 10045 16945
<< nsubstratencontact >>
rect 10145 16895 10195 16945
<< psubstratepcontact >>
rect 65 16745 115 16795
<< psubstratepcontact >>
rect 215 16745 265 16795
<< nsubstratencontact >>
rect 605 16745 655 16795
<< nsubstratencontact >>
rect 755 16745 805 16795
<< polycontact >>
rect 995 16775 1045 16825
<< pdcontact >>
rect 1265 16745 1315 16795
<< pdcontact >>
rect 1415 16745 1465 16795
<< pdcontact >>
rect 1565 16745 1615 16795
<< pdcontact >>
rect 1715 16745 1765 16795
<< pdcontact >>
rect 1865 16745 1915 16795
<< pdcontact >>
rect 2015 16745 2065 16795
<< pdcontact >>
rect 2165 16745 2215 16795
<< pdcontact >>
rect 2315 16745 2365 16795
<< pdcontact >>
rect 2465 16745 2515 16795
<< pdcontact >>
rect 2615 16745 2665 16795
<< pdcontact >>
rect 2765 16745 2815 16795
<< pdcontact >>
rect 2915 16745 2965 16795
<< pdcontact >>
rect 3065 16745 3115 16795
<< pdcontact >>
rect 3215 16745 3265 16795
<< pdcontact >>
rect 3365 16745 3415 16795
<< pdcontact >>
rect 3515 16745 3565 16795
<< pdcontact >>
rect 3665 16745 3715 16795
<< pdcontact >>
rect 3815 16745 3865 16795
<< pdcontact >>
rect 3965 16745 4015 16795
<< pdcontact >>
rect 4115 16745 4165 16795
<< pdcontact >>
rect 4265 16745 4315 16795
<< pdcontact >>
rect 4415 16745 4465 16795
<< pdcontact >>
rect 4565 16745 4615 16795
<< pdcontact >>
rect 4715 16745 4765 16795
<< pdcontact >>
rect 4865 16745 4915 16795
<< polycontact >>
rect 5075 16775 5125 16825
<< nsubstratencontact >>
rect 5315 16745 5365 16795
<< nsubstratencontact >>
rect 5465 16745 5515 16795
<< polycontact >>
rect 5675 16775 5725 16825
<< pdcontact >>
rect 5885 16745 5935 16795
<< pdcontact >>
rect 6035 16745 6085 16795
<< pdcontact >>
rect 6185 16745 6235 16795
<< pdcontact >>
rect 6335 16745 6385 16795
<< pdcontact >>
rect 6485 16745 6535 16795
<< pdcontact >>
rect 6635 16745 6685 16795
<< pdcontact >>
rect 6785 16745 6835 16795
<< pdcontact >>
rect 6935 16745 6985 16795
<< pdcontact >>
rect 7085 16745 7135 16795
<< pdcontact >>
rect 7235 16745 7285 16795
<< pdcontact >>
rect 7385 16745 7435 16795
<< pdcontact >>
rect 7535 16745 7585 16795
<< pdcontact >>
rect 7685 16745 7735 16795
<< pdcontact >>
rect 7835 16745 7885 16795
<< pdcontact >>
rect 7985 16745 8035 16795
<< pdcontact >>
rect 8135 16745 8185 16795
<< pdcontact >>
rect 8285 16745 8335 16795
<< pdcontact >>
rect 8435 16745 8485 16795
<< pdcontact >>
rect 8585 16745 8635 16795
<< pdcontact >>
rect 8735 16745 8785 16795
<< pdcontact >>
rect 8885 16745 8935 16795
<< pdcontact >>
rect 9035 16745 9085 16795
<< pdcontact >>
rect 9185 16745 9235 16795
<< pdcontact >>
rect 9335 16745 9385 16795
<< pdcontact >>
rect 9485 16745 9535 16795
<< polycontact >>
rect 9755 16775 9805 16825
<< nsubstratencontact >>
rect 9995 16745 10045 16795
<< nsubstratencontact >>
rect 10145 16745 10195 16795
<< psubstratepcontact >>
rect 10535 16745 10585 16795
<< psubstratepcontact >>
rect 10685 16745 10735 16795
<< nsubstratencontact >>
rect 605 16595 655 16645
<< nsubstratencontact >>
rect 755 16595 805 16645
<< polycontact >>
rect 995 16625 1045 16675
<< pdcontact >>
rect 1265 16595 1315 16645
<< pdcontact >>
rect 1415 16595 1465 16645
<< pdcontact >>
rect 1565 16595 1615 16645
<< pdcontact >>
rect 1715 16595 1765 16645
<< pdcontact >>
rect 1865 16595 1915 16645
<< pdcontact >>
rect 2015 16595 2065 16645
<< pdcontact >>
rect 2165 16595 2215 16645
<< pdcontact >>
rect 2315 16595 2365 16645
<< pdcontact >>
rect 2465 16595 2515 16645
<< pdcontact >>
rect 2615 16595 2665 16645
<< pdcontact >>
rect 2765 16595 2815 16645
<< pdcontact >>
rect 2915 16595 2965 16645
<< pdcontact >>
rect 3065 16595 3115 16645
<< pdcontact >>
rect 3215 16595 3265 16645
<< pdcontact >>
rect 3365 16595 3415 16645
<< pdcontact >>
rect 3515 16595 3565 16645
<< pdcontact >>
rect 3665 16595 3715 16645
<< pdcontact >>
rect 3815 16595 3865 16645
<< pdcontact >>
rect 3965 16595 4015 16645
<< pdcontact >>
rect 4115 16595 4165 16645
<< pdcontact >>
rect 4265 16595 4315 16645
<< pdcontact >>
rect 4415 16595 4465 16645
<< pdcontact >>
rect 4565 16595 4615 16645
<< pdcontact >>
rect 4715 16595 4765 16645
<< pdcontact >>
rect 4865 16595 4915 16645
<< polycontact >>
rect 5075 16625 5125 16675
<< nsubstratencontact >>
rect 5315 16595 5365 16645
<< nsubstratencontact >>
rect 5465 16595 5515 16645
<< polycontact >>
rect 5675 16625 5725 16675
<< pdcontact >>
rect 5885 16595 5935 16645
<< pdcontact >>
rect 6035 16595 6085 16645
<< pdcontact >>
rect 6185 16595 6235 16645
<< pdcontact >>
rect 6335 16595 6385 16645
<< pdcontact >>
rect 6485 16595 6535 16645
<< pdcontact >>
rect 6635 16595 6685 16645
<< pdcontact >>
rect 6785 16595 6835 16645
<< pdcontact >>
rect 6935 16595 6985 16645
<< pdcontact >>
rect 7085 16595 7135 16645
<< pdcontact >>
rect 7235 16595 7285 16645
<< pdcontact >>
rect 7385 16595 7435 16645
<< pdcontact >>
rect 7535 16595 7585 16645
<< pdcontact >>
rect 7685 16595 7735 16645
<< pdcontact >>
rect 7835 16595 7885 16645
<< pdcontact >>
rect 7985 16595 8035 16645
<< pdcontact >>
rect 8135 16595 8185 16645
<< pdcontact >>
rect 8285 16595 8335 16645
<< pdcontact >>
rect 8435 16595 8485 16645
<< pdcontact >>
rect 8585 16595 8635 16645
<< pdcontact >>
rect 8735 16595 8785 16645
<< pdcontact >>
rect 8885 16595 8935 16645
<< pdcontact >>
rect 9035 16595 9085 16645
<< pdcontact >>
rect 9185 16595 9235 16645
<< pdcontact >>
rect 9335 16595 9385 16645
<< pdcontact >>
rect 9485 16595 9535 16645
<< polycontact >>
rect 9755 16625 9805 16675
<< nsubstratencontact >>
rect 9995 16595 10045 16645
<< nsubstratencontact >>
rect 10145 16595 10195 16645
<< psubstratepcontact >>
rect 65 16475 115 16525
<< psubstratepcontact >>
rect 215 16475 265 16525
<< nsubstratencontact >>
rect 605 16445 655 16495
<< nsubstratencontact >>
rect 755 16445 805 16495
<< polycontact >>
rect 995 16475 1045 16525
<< pdcontact >>
rect 1265 16445 1315 16495
<< pdcontact >>
rect 1415 16445 1465 16495
<< pdcontact >>
rect 1565 16445 1615 16495
<< pdcontact >>
rect 1715 16445 1765 16495
<< pdcontact >>
rect 1865 16445 1915 16495
<< pdcontact >>
rect 2015 16445 2065 16495
<< pdcontact >>
rect 2165 16445 2215 16495
<< pdcontact >>
rect 2315 16445 2365 16495
<< pdcontact >>
rect 2465 16445 2515 16495
<< pdcontact >>
rect 2615 16445 2665 16495
<< pdcontact >>
rect 2765 16445 2815 16495
<< pdcontact >>
rect 2915 16445 2965 16495
<< pdcontact >>
rect 3065 16445 3115 16495
<< pdcontact >>
rect 3215 16445 3265 16495
<< pdcontact >>
rect 3365 16445 3415 16495
<< pdcontact >>
rect 3515 16445 3565 16495
<< pdcontact >>
rect 3665 16445 3715 16495
<< pdcontact >>
rect 3815 16445 3865 16495
<< pdcontact >>
rect 3965 16445 4015 16495
<< pdcontact >>
rect 4115 16445 4165 16495
<< pdcontact >>
rect 4265 16445 4315 16495
<< pdcontact >>
rect 4415 16445 4465 16495
<< pdcontact >>
rect 4565 16445 4615 16495
<< pdcontact >>
rect 4715 16445 4765 16495
<< pdcontact >>
rect 4865 16445 4915 16495
<< polycontact >>
rect 5075 16475 5125 16525
<< nsubstratencontact >>
rect 5315 16445 5365 16495
<< nsubstratencontact >>
rect 5465 16445 5515 16495
<< polycontact >>
rect 5675 16475 5725 16525
<< pdcontact >>
rect 5885 16445 5935 16495
<< pdcontact >>
rect 6035 16445 6085 16495
<< pdcontact >>
rect 6185 16445 6235 16495
<< pdcontact >>
rect 6335 16445 6385 16495
<< pdcontact >>
rect 6485 16445 6535 16495
<< pdcontact >>
rect 6635 16445 6685 16495
<< pdcontact >>
rect 6785 16445 6835 16495
<< pdcontact >>
rect 6935 16445 6985 16495
<< pdcontact >>
rect 7085 16445 7135 16495
<< pdcontact >>
rect 7235 16445 7285 16495
<< pdcontact >>
rect 7385 16445 7435 16495
<< pdcontact >>
rect 7535 16445 7585 16495
<< pdcontact >>
rect 7685 16445 7735 16495
<< pdcontact >>
rect 7835 16445 7885 16495
<< pdcontact >>
rect 7985 16445 8035 16495
<< pdcontact >>
rect 8135 16445 8185 16495
<< pdcontact >>
rect 8285 16445 8335 16495
<< pdcontact >>
rect 8435 16445 8485 16495
<< pdcontact >>
rect 8585 16445 8635 16495
<< pdcontact >>
rect 8735 16445 8785 16495
<< pdcontact >>
rect 8885 16445 8935 16495
<< pdcontact >>
rect 9035 16445 9085 16495
<< pdcontact >>
rect 9185 16445 9235 16495
<< pdcontact >>
rect 9335 16445 9385 16495
<< pdcontact >>
rect 9485 16445 9535 16495
<< polycontact >>
rect 9755 16475 9805 16525
<< nsubstratencontact >>
rect 9995 16445 10045 16495
<< nsubstratencontact >>
rect 10145 16445 10195 16495
<< psubstratepcontact >>
rect 10535 16475 10585 16525
<< psubstratepcontact >>
rect 10685 16475 10735 16525
<< nsubstratencontact >>
rect 605 16295 655 16345
<< nsubstratencontact >>
rect 755 16295 805 16345
<< polycontact >>
rect 995 16325 1045 16375
<< polycontact >>
rect 5075 16325 5125 16375
<< nsubstratencontact >>
rect 5315 16295 5365 16345
<< nsubstratencontact >>
rect 5465 16295 5515 16345
<< polycontact >>
rect 5675 16325 5725 16375
<< polycontact >>
rect 9755 16325 9805 16375
<< nsubstratencontact >>
rect 9995 16295 10045 16345
<< nsubstratencontact >>
rect 10145 16295 10195 16345
<< psubstratepcontact >>
rect 65 16235 115 16285
<< psubstratepcontact >>
rect 215 16235 265 16285
<< psubstratepcontact >>
rect 10535 16235 10585 16285
<< psubstratepcontact >>
rect 10685 16235 10735 16285
<< polycontact >>
rect 995 16175 1045 16225
<< pdcontact >>
rect 1235 16145 1285 16195
<< pdcontact >>
rect 1535 16145 1585 16195
<< pdcontact >>
rect 1835 16145 1885 16195
<< pdcontact >>
rect 2135 16145 2185 16195
<< pdcontact >>
rect 2435 16145 2485 16195
<< pdcontact >>
rect 2735 16145 2785 16195
<< pdcontact >>
rect 3035 16145 3085 16195
<< pdcontact >>
rect 3335 16145 3385 16195
<< pdcontact >>
rect 4505 16145 4555 16195
<< pdcontact >>
rect 4805 16145 4855 16195
<< polycontact >>
rect 5075 16175 5125 16225
<< polycontact >>
rect 5675 16175 5725 16225
<< pdcontact >>
rect 5945 16145 5995 16195
<< pdcontact >>
rect 6245 16145 6295 16195
<< pdcontact >>
rect 7415 16145 7465 16195
<< pdcontact >>
rect 7715 16145 7765 16195
<< pdcontact >>
rect 8015 16145 8065 16195
<< pdcontact >>
rect 8315 16145 8365 16195
<< pdcontact >>
rect 8615 16145 8665 16195
<< pdcontact >>
rect 8915 16145 8965 16195
<< pdcontact >>
rect 9215 16145 9265 16195
<< pdcontact >>
rect 9515 16145 9565 16195
<< polycontact >>
rect 9755 16175 9805 16225
<< psubstratepcontact >>
rect 65 15995 115 16045
<< psubstratepcontact >>
rect 215 15995 265 16045
<< polycontact >>
rect 995 16025 1045 16075
<< pdcontact >>
rect 1235 15995 1285 16045
<< pdcontact >>
rect 1535 15995 1585 16045
<< pdcontact >>
rect 1835 15995 1885 16045
<< pdcontact >>
rect 2135 15995 2185 16045
<< pdcontact >>
rect 2435 15995 2485 16045
<< pdcontact >>
rect 2735 15995 2785 16045
<< pdcontact >>
rect 3035 15995 3085 16045
<< pdcontact >>
rect 3335 15995 3385 16045
<< pdcontact >>
rect 4505 15995 4555 16045
<< pdcontact >>
rect 4805 15995 4855 16045
<< polycontact >>
rect 5075 16025 5125 16075
<< polycontact >>
rect 5675 16025 5725 16075
<< pdcontact >>
rect 5945 15995 5995 16045
<< pdcontact >>
rect 6245 15995 6295 16045
<< pdcontact >>
rect 7415 15995 7465 16045
<< pdcontact >>
rect 7715 15995 7765 16045
<< pdcontact >>
rect 8015 15995 8065 16045
<< pdcontact >>
rect 8315 15995 8365 16045
<< pdcontact >>
rect 8615 15995 8665 16045
<< pdcontact >>
rect 8915 15995 8965 16045
<< pdcontact >>
rect 9215 15995 9265 16045
<< pdcontact >>
rect 9515 15995 9565 16045
<< polycontact >>
rect 9755 16025 9805 16075
<< psubstratepcontact >>
rect 10535 15995 10585 16045
<< psubstratepcontact >>
rect 10685 15995 10735 16045
<< polycontact >>
rect 995 15875 1045 15925
<< pdcontact >>
rect 1235 15845 1285 15895
<< pdcontact >>
rect 1535 15845 1585 15895
<< pdcontact >>
rect 1835 15845 1885 15895
<< pdcontact >>
rect 2135 15845 2185 15895
<< pdcontact >>
rect 2435 15845 2485 15895
<< pdcontact >>
rect 2735 15845 2785 15895
<< pdcontact >>
rect 3035 15845 3085 15895
<< pdcontact >>
rect 3335 15845 3385 15895
<< pdcontact >>
rect 4505 15845 4555 15895
<< pdcontact >>
rect 4805 15845 4855 15895
<< polycontact >>
rect 5075 15875 5125 15925
<< polycontact >>
rect 5675 15875 5725 15925
<< pdcontact >>
rect 5945 15845 5995 15895
<< pdcontact >>
rect 6245 15845 6295 15895
<< pdcontact >>
rect 7415 15845 7465 15895
<< pdcontact >>
rect 7715 15845 7765 15895
<< pdcontact >>
rect 8015 15845 8065 15895
<< pdcontact >>
rect 8315 15845 8365 15895
<< pdcontact >>
rect 8615 15845 8665 15895
<< pdcontact >>
rect 8915 15845 8965 15895
<< pdcontact >>
rect 9215 15845 9265 15895
<< pdcontact >>
rect 9515 15845 9565 15895
<< polycontact >>
rect 9755 15875 9805 15925
<< psubstratepcontact >>
rect 65 15755 115 15805
<< psubstratepcontact >>
rect 215 15755 265 15805
<< nsubstratencontact >>
rect 605 15695 655 15745
<< nsubstratencontact >>
rect 755 15695 805 15745
<< polycontact >>
rect 995 15725 1045 15775
<< polycontact >>
rect 5075 15725 5125 15775
<< nsubstratencontact >>
rect 5315 15695 5365 15745
<< nsubstratencontact >>
rect 5465 15695 5515 15745
<< polycontact >>
rect 5675 15725 5725 15775
<< polycontact >>
rect 9755 15725 9805 15775
<< psubstratepcontact >>
rect 10535 15755 10585 15805
<< psubstratepcontact >>
rect 10685 15755 10735 15805
<< nsubstratencontact >>
rect 9995 15695 10045 15745
<< nsubstratencontact >>
rect 10145 15695 10195 15745
<< psubstratepcontact >>
rect 65 15515 115 15565
<< psubstratepcontact >>
rect 215 15515 265 15565
<< nsubstratencontact >>
rect 605 15545 655 15595
<< nsubstratencontact >>
rect 755 15545 805 15595
<< polycontact >>
rect 995 15575 1045 15625
<< pdcontact >>
rect 1265 15545 1315 15595
<< pdcontact >>
rect 1415 15545 1465 15595
<< pdcontact >>
rect 1565 15545 1615 15595
<< pdcontact >>
rect 1715 15545 1765 15595
<< pdcontact >>
rect 1865 15545 1915 15595
<< pdcontact >>
rect 2015 15545 2065 15595
<< pdcontact >>
rect 2165 15545 2215 15595
<< pdcontact >>
rect 2315 15545 2365 15595
<< pdcontact >>
rect 2465 15545 2515 15595
<< pdcontact >>
rect 2615 15545 2665 15595
<< pdcontact >>
rect 2765 15545 2815 15595
<< pdcontact >>
rect 2915 15545 2965 15595
<< pdcontact >>
rect 3065 15545 3115 15595
<< pdcontact >>
rect 3215 15545 3265 15595
<< pdcontact >>
rect 3365 15545 3415 15595
<< pdcontact >>
rect 3515 15545 3565 15595
<< pdcontact >>
rect 3665 15545 3715 15595
<< pdcontact >>
rect 3815 15545 3865 15595
<< pdcontact >>
rect 3965 15545 4015 15595
<< pdcontact >>
rect 4115 15545 4165 15595
<< pdcontact >>
rect 4265 15545 4315 15595
<< pdcontact >>
rect 4415 15545 4465 15595
<< pdcontact >>
rect 4565 15545 4615 15595
<< pdcontact >>
rect 4715 15545 4765 15595
<< pdcontact >>
rect 4865 15545 4915 15595
<< polycontact >>
rect 5075 15575 5125 15625
<< nsubstratencontact >>
rect 5315 15545 5365 15595
<< nsubstratencontact >>
rect 5465 15545 5515 15595
<< polycontact >>
rect 5675 15575 5725 15625
<< pdcontact >>
rect 5885 15545 5935 15595
<< pdcontact >>
rect 6035 15545 6085 15595
<< pdcontact >>
rect 6185 15545 6235 15595
<< pdcontact >>
rect 6335 15545 6385 15595
<< pdcontact >>
rect 6485 15545 6535 15595
<< pdcontact >>
rect 6635 15545 6685 15595
<< pdcontact >>
rect 6785 15545 6835 15595
<< pdcontact >>
rect 6935 15545 6985 15595
<< pdcontact >>
rect 7085 15545 7135 15595
<< pdcontact >>
rect 7235 15545 7285 15595
<< pdcontact >>
rect 7385 15545 7435 15595
<< pdcontact >>
rect 7535 15545 7585 15595
<< pdcontact >>
rect 7685 15545 7735 15595
<< pdcontact >>
rect 7835 15545 7885 15595
<< pdcontact >>
rect 7985 15545 8035 15595
<< pdcontact >>
rect 8135 15545 8185 15595
<< pdcontact >>
rect 8285 15545 8335 15595
<< pdcontact >>
rect 8435 15545 8485 15595
<< pdcontact >>
rect 8585 15545 8635 15595
<< pdcontact >>
rect 8735 15545 8785 15595
<< pdcontact >>
rect 8885 15545 8935 15595
<< pdcontact >>
rect 9035 15545 9085 15595
<< pdcontact >>
rect 9185 15545 9235 15595
<< pdcontact >>
rect 9335 15545 9385 15595
<< pdcontact >>
rect 9485 15545 9535 15595
<< polycontact >>
rect 9755 15575 9805 15625
<< nsubstratencontact >>
rect 9995 15545 10045 15595
<< nsubstratencontact >>
rect 10145 15545 10195 15595
<< psubstratepcontact >>
rect 10535 15515 10585 15565
<< psubstratepcontact >>
rect 10685 15515 10735 15565
<< nsubstratencontact >>
rect 605 15395 655 15445
<< nsubstratencontact >>
rect 755 15395 805 15445
<< polycontact >>
rect 995 15425 1045 15475
<< pdcontact >>
rect 1265 15395 1315 15445
<< pdcontact >>
rect 1415 15395 1465 15445
<< pdcontact >>
rect 1565 15395 1615 15445
<< pdcontact >>
rect 1715 15395 1765 15445
<< pdcontact >>
rect 1865 15395 1915 15445
<< pdcontact >>
rect 2015 15395 2065 15445
<< pdcontact >>
rect 2165 15395 2215 15445
<< pdcontact >>
rect 2315 15395 2365 15445
<< pdcontact >>
rect 2465 15395 2515 15445
<< pdcontact >>
rect 2615 15395 2665 15445
<< pdcontact >>
rect 2765 15395 2815 15445
<< pdcontact >>
rect 2915 15395 2965 15445
<< pdcontact >>
rect 3065 15395 3115 15445
<< pdcontact >>
rect 3215 15395 3265 15445
<< pdcontact >>
rect 3365 15395 3415 15445
<< pdcontact >>
rect 3515 15395 3565 15445
<< pdcontact >>
rect 3665 15395 3715 15445
<< pdcontact >>
rect 3815 15395 3865 15445
<< pdcontact >>
rect 3965 15395 4015 15445
<< pdcontact >>
rect 4115 15395 4165 15445
<< pdcontact >>
rect 4265 15395 4315 15445
<< pdcontact >>
rect 4415 15395 4465 15445
<< pdcontact >>
rect 4565 15395 4615 15445
<< pdcontact >>
rect 4715 15395 4765 15445
<< pdcontact >>
rect 4865 15395 4915 15445
<< polycontact >>
rect 5075 15425 5125 15475
<< nsubstratencontact >>
rect 5315 15395 5365 15445
<< nsubstratencontact >>
rect 5465 15395 5515 15445
<< polycontact >>
rect 5675 15425 5725 15475
<< pdcontact >>
rect 5885 15395 5935 15445
<< pdcontact >>
rect 6035 15395 6085 15445
<< pdcontact >>
rect 6185 15395 6235 15445
<< pdcontact >>
rect 6335 15395 6385 15445
<< pdcontact >>
rect 6485 15395 6535 15445
<< pdcontact >>
rect 6635 15395 6685 15445
<< pdcontact >>
rect 6785 15395 6835 15445
<< pdcontact >>
rect 6935 15395 6985 15445
<< pdcontact >>
rect 7085 15395 7135 15445
<< pdcontact >>
rect 7235 15395 7285 15445
<< pdcontact >>
rect 7385 15395 7435 15445
<< pdcontact >>
rect 7535 15395 7585 15445
<< pdcontact >>
rect 7685 15395 7735 15445
<< pdcontact >>
rect 7835 15395 7885 15445
<< pdcontact >>
rect 7985 15395 8035 15445
<< pdcontact >>
rect 8135 15395 8185 15445
<< pdcontact >>
rect 8285 15395 8335 15445
<< pdcontact >>
rect 8435 15395 8485 15445
<< pdcontact >>
rect 8585 15395 8635 15445
<< pdcontact >>
rect 8735 15395 8785 15445
<< pdcontact >>
rect 8885 15395 8935 15445
<< pdcontact >>
rect 9035 15395 9085 15445
<< pdcontact >>
rect 9185 15395 9235 15445
<< pdcontact >>
rect 9335 15395 9385 15445
<< pdcontact >>
rect 9485 15395 9535 15445
<< polycontact >>
rect 9755 15425 9805 15475
<< nsubstratencontact >>
rect 9995 15395 10045 15445
<< nsubstratencontact >>
rect 10145 15395 10195 15445
<< psubstratepcontact >>
rect 65 15275 115 15325
<< psubstratepcontact >>
rect 215 15275 265 15325
<< nsubstratencontact >>
rect 605 15245 655 15295
<< nsubstratencontact >>
rect 755 15245 805 15295
<< polycontact >>
rect 995 15275 1045 15325
<< pdcontact >>
rect 1265 15245 1315 15295
<< pdcontact >>
rect 1415 15245 1465 15295
<< pdcontact >>
rect 1565 15245 1615 15295
<< pdcontact >>
rect 1715 15245 1765 15295
<< pdcontact >>
rect 1865 15245 1915 15295
<< pdcontact >>
rect 2015 15245 2065 15295
<< pdcontact >>
rect 2165 15245 2215 15295
<< pdcontact >>
rect 2315 15245 2365 15295
<< pdcontact >>
rect 2465 15245 2515 15295
<< pdcontact >>
rect 2615 15245 2665 15295
<< pdcontact >>
rect 2765 15245 2815 15295
<< pdcontact >>
rect 2915 15245 2965 15295
<< pdcontact >>
rect 3065 15245 3115 15295
<< pdcontact >>
rect 3215 15245 3265 15295
<< pdcontact >>
rect 3365 15245 3415 15295
<< pdcontact >>
rect 3515 15245 3565 15295
<< pdcontact >>
rect 3665 15245 3715 15295
<< pdcontact >>
rect 3815 15245 3865 15295
<< pdcontact >>
rect 3965 15245 4015 15295
<< pdcontact >>
rect 4115 15245 4165 15295
<< pdcontact >>
rect 4265 15245 4315 15295
<< pdcontact >>
rect 4415 15245 4465 15295
<< pdcontact >>
rect 4565 15245 4615 15295
<< pdcontact >>
rect 4715 15245 4765 15295
<< pdcontact >>
rect 4865 15245 4915 15295
<< polycontact >>
rect 5075 15275 5125 15325
<< nsubstratencontact >>
rect 5315 15245 5365 15295
<< nsubstratencontact >>
rect 5465 15245 5515 15295
<< polycontact >>
rect 5675 15275 5725 15325
<< pdcontact >>
rect 5885 15245 5935 15295
<< pdcontact >>
rect 6035 15245 6085 15295
<< pdcontact >>
rect 6185 15245 6235 15295
<< pdcontact >>
rect 6335 15245 6385 15295
<< pdcontact >>
rect 6485 15245 6535 15295
<< pdcontact >>
rect 6635 15245 6685 15295
<< pdcontact >>
rect 6785 15245 6835 15295
<< pdcontact >>
rect 6935 15245 6985 15295
<< pdcontact >>
rect 7085 15245 7135 15295
<< pdcontact >>
rect 7235 15245 7285 15295
<< pdcontact >>
rect 7385 15245 7435 15295
<< pdcontact >>
rect 7535 15245 7585 15295
<< pdcontact >>
rect 7685 15245 7735 15295
<< pdcontact >>
rect 7835 15245 7885 15295
<< pdcontact >>
rect 7985 15245 8035 15295
<< pdcontact >>
rect 8135 15245 8185 15295
<< pdcontact >>
rect 8285 15245 8335 15295
<< pdcontact >>
rect 8435 15245 8485 15295
<< pdcontact >>
rect 8585 15245 8635 15295
<< pdcontact >>
rect 8735 15245 8785 15295
<< pdcontact >>
rect 8885 15245 8935 15295
<< pdcontact >>
rect 9035 15245 9085 15295
<< pdcontact >>
rect 9185 15245 9235 15295
<< pdcontact >>
rect 9335 15245 9385 15295
<< pdcontact >>
rect 9485 15245 9535 15295
<< polycontact >>
rect 9755 15275 9805 15325
<< nsubstratencontact >>
rect 9995 15245 10045 15295
<< nsubstratencontact >>
rect 10145 15245 10195 15295
<< psubstratepcontact >>
rect 10535 15275 10585 15325
<< psubstratepcontact >>
rect 10685 15275 10735 15325
<< nsubstratencontact >>
rect 605 15095 655 15145
<< nsubstratencontact >>
rect 755 15095 805 15145
<< polycontact >>
rect 995 15125 1045 15175
<< pdcontact >>
rect 1265 15095 1315 15145
<< pdcontact >>
rect 1415 15095 1465 15145
<< pdcontact >>
rect 1565 15095 1615 15145
<< pdcontact >>
rect 1715 15095 1765 15145
<< pdcontact >>
rect 1865 15095 1915 15145
<< pdcontact >>
rect 2015 15095 2065 15145
<< pdcontact >>
rect 2165 15095 2215 15145
<< pdcontact >>
rect 2315 15095 2365 15145
<< pdcontact >>
rect 2465 15095 2515 15145
<< pdcontact >>
rect 2615 15095 2665 15145
<< pdcontact >>
rect 2765 15095 2815 15145
<< pdcontact >>
rect 2915 15095 2965 15145
<< pdcontact >>
rect 3065 15095 3115 15145
<< pdcontact >>
rect 3215 15095 3265 15145
<< pdcontact >>
rect 3365 15095 3415 15145
<< pdcontact >>
rect 3515 15095 3565 15145
<< pdcontact >>
rect 3665 15095 3715 15145
<< pdcontact >>
rect 3815 15095 3865 15145
<< pdcontact >>
rect 3965 15095 4015 15145
<< pdcontact >>
rect 4115 15095 4165 15145
<< pdcontact >>
rect 4265 15095 4315 15145
<< pdcontact >>
rect 4415 15095 4465 15145
<< pdcontact >>
rect 4565 15095 4615 15145
<< pdcontact >>
rect 4715 15095 4765 15145
<< pdcontact >>
rect 4865 15095 4915 15145
<< polycontact >>
rect 5075 15125 5125 15175
<< nsubstratencontact >>
rect 5315 15095 5365 15145
<< nsubstratencontact >>
rect 5465 15095 5515 15145
<< polycontact >>
rect 5675 15125 5725 15175
<< pdcontact >>
rect 5885 15095 5935 15145
<< pdcontact >>
rect 6035 15095 6085 15145
<< pdcontact >>
rect 6185 15095 6235 15145
<< pdcontact >>
rect 6335 15095 6385 15145
<< pdcontact >>
rect 6485 15095 6535 15145
<< pdcontact >>
rect 6635 15095 6685 15145
<< pdcontact >>
rect 6785 15095 6835 15145
<< pdcontact >>
rect 6935 15095 6985 15145
<< pdcontact >>
rect 7085 15095 7135 15145
<< pdcontact >>
rect 7235 15095 7285 15145
<< pdcontact >>
rect 7385 15095 7435 15145
<< pdcontact >>
rect 7535 15095 7585 15145
<< pdcontact >>
rect 7685 15095 7735 15145
<< pdcontact >>
rect 7835 15095 7885 15145
<< pdcontact >>
rect 7985 15095 8035 15145
<< pdcontact >>
rect 8135 15095 8185 15145
<< pdcontact >>
rect 8285 15095 8335 15145
<< pdcontact >>
rect 8435 15095 8485 15145
<< pdcontact >>
rect 8585 15095 8635 15145
<< pdcontact >>
rect 8735 15095 8785 15145
<< pdcontact >>
rect 8885 15095 8935 15145
<< pdcontact >>
rect 9035 15095 9085 15145
<< pdcontact >>
rect 9185 15095 9235 15145
<< pdcontact >>
rect 9335 15095 9385 15145
<< pdcontact >>
rect 9485 15095 9535 15145
<< polycontact >>
rect 9755 15125 9805 15175
<< nsubstratencontact >>
rect 9995 15095 10045 15145
<< nsubstratencontact >>
rect 10145 15095 10195 15145
<< psubstratepcontact >>
rect 65 15035 115 15085
<< psubstratepcontact >>
rect 215 15035 265 15085
<< psubstratepcontact >>
rect 10535 15035 10585 15085
<< psubstratepcontact >>
rect 10685 15035 10735 15085
<< nsubstratencontact >>
rect 605 14945 655 14995
<< nsubstratencontact >>
rect 755 14945 805 14995
<< polycontact >>
rect 995 14975 1045 15025
<< pdcontact >>
rect 1265 14945 1315 14995
<< pdcontact >>
rect 1415 14945 1465 14995
<< pdcontact >>
rect 1565 14945 1615 14995
<< pdcontact >>
rect 1715 14945 1765 14995
<< pdcontact >>
rect 1865 14945 1915 14995
<< pdcontact >>
rect 2015 14945 2065 14995
<< pdcontact >>
rect 2165 14945 2215 14995
<< pdcontact >>
rect 2315 14945 2365 14995
<< pdcontact >>
rect 2465 14945 2515 14995
<< pdcontact >>
rect 2615 14945 2665 14995
<< pdcontact >>
rect 2765 14945 2815 14995
<< pdcontact >>
rect 2915 14945 2965 14995
<< pdcontact >>
rect 3065 14945 3115 14995
<< pdcontact >>
rect 3215 14945 3265 14995
<< pdcontact >>
rect 3365 14945 3415 14995
<< pdcontact >>
rect 3515 14945 3565 14995
<< pdcontact >>
rect 3665 14945 3715 14995
<< pdcontact >>
rect 3815 14945 3865 14995
<< pdcontact >>
rect 3965 14945 4015 14995
<< pdcontact >>
rect 4115 14945 4165 14995
<< pdcontact >>
rect 4265 14945 4315 14995
<< pdcontact >>
rect 4415 14945 4465 14995
<< pdcontact >>
rect 4565 14945 4615 14995
<< pdcontact >>
rect 4715 14945 4765 14995
<< pdcontact >>
rect 4865 14945 4915 14995
<< polycontact >>
rect 5075 14975 5125 15025
<< nsubstratencontact >>
rect 5315 14945 5365 14995
<< nsubstratencontact >>
rect 5465 14945 5515 14995
<< polycontact >>
rect 5675 14975 5725 15025
<< pdcontact >>
rect 5885 14945 5935 14995
<< pdcontact >>
rect 6035 14945 6085 14995
<< pdcontact >>
rect 6185 14945 6235 14995
<< pdcontact >>
rect 6335 14945 6385 14995
<< pdcontact >>
rect 6485 14945 6535 14995
<< pdcontact >>
rect 6635 14945 6685 14995
<< pdcontact >>
rect 6785 14945 6835 14995
<< pdcontact >>
rect 6935 14945 6985 14995
<< pdcontact >>
rect 7085 14945 7135 14995
<< pdcontact >>
rect 7235 14945 7285 14995
<< pdcontact >>
rect 7385 14945 7435 14995
<< pdcontact >>
rect 7535 14945 7585 14995
<< pdcontact >>
rect 7685 14945 7735 14995
<< pdcontact >>
rect 7835 14945 7885 14995
<< pdcontact >>
rect 7985 14945 8035 14995
<< pdcontact >>
rect 8135 14945 8185 14995
<< pdcontact >>
rect 8285 14945 8335 14995
<< pdcontact >>
rect 8435 14945 8485 14995
<< pdcontact >>
rect 8585 14945 8635 14995
<< pdcontact >>
rect 8735 14945 8785 14995
<< pdcontact >>
rect 8885 14945 8935 14995
<< pdcontact >>
rect 9035 14945 9085 14995
<< pdcontact >>
rect 9185 14945 9235 14995
<< pdcontact >>
rect 9335 14945 9385 14995
<< pdcontact >>
rect 9485 14945 9535 14995
<< polycontact >>
rect 9755 14975 9805 15025
<< nsubstratencontact >>
rect 9995 14945 10045 14995
<< nsubstratencontact >>
rect 10145 14945 10195 14995
<< psubstratepcontact >>
rect 65 14795 115 14845
<< psubstratepcontact >>
rect 215 14795 265 14845
<< nsubstratencontact >>
rect 605 14795 655 14845
<< nsubstratencontact >>
rect 755 14795 805 14845
<< polycontact >>
rect 995 14825 1045 14875
<< pdcontact >>
rect 1265 14795 1315 14845
<< pdcontact >>
rect 1415 14795 1465 14845
<< pdcontact >>
rect 1565 14795 1615 14845
<< pdcontact >>
rect 1715 14795 1765 14845
<< pdcontact >>
rect 1865 14795 1915 14845
<< pdcontact >>
rect 2015 14795 2065 14845
<< pdcontact >>
rect 2165 14795 2215 14845
<< pdcontact >>
rect 2315 14795 2365 14845
<< pdcontact >>
rect 2465 14795 2515 14845
<< pdcontact >>
rect 2615 14795 2665 14845
<< pdcontact >>
rect 2765 14795 2815 14845
<< pdcontact >>
rect 2915 14795 2965 14845
<< pdcontact >>
rect 3065 14795 3115 14845
<< pdcontact >>
rect 3215 14795 3265 14845
<< pdcontact >>
rect 3365 14795 3415 14845
<< pdcontact >>
rect 3515 14795 3565 14845
<< pdcontact >>
rect 3665 14795 3715 14845
<< pdcontact >>
rect 3815 14795 3865 14845
<< pdcontact >>
rect 3965 14795 4015 14845
<< pdcontact >>
rect 4115 14795 4165 14845
<< pdcontact >>
rect 4265 14795 4315 14845
<< pdcontact >>
rect 4415 14795 4465 14845
<< pdcontact >>
rect 4565 14795 4615 14845
<< pdcontact >>
rect 4715 14795 4765 14845
<< pdcontact >>
rect 4865 14795 4915 14845
<< polycontact >>
rect 5075 14825 5125 14875
<< nsubstratencontact >>
rect 5315 14795 5365 14845
<< nsubstratencontact >>
rect 5465 14795 5515 14845
<< polycontact >>
rect 5675 14825 5725 14875
<< pdcontact >>
rect 5885 14795 5935 14845
<< pdcontact >>
rect 6035 14795 6085 14845
<< pdcontact >>
rect 6185 14795 6235 14845
<< pdcontact >>
rect 6335 14795 6385 14845
<< pdcontact >>
rect 6485 14795 6535 14845
<< pdcontact >>
rect 6635 14795 6685 14845
<< pdcontact >>
rect 6785 14795 6835 14845
<< pdcontact >>
rect 6935 14795 6985 14845
<< pdcontact >>
rect 7085 14795 7135 14845
<< pdcontact >>
rect 7235 14795 7285 14845
<< pdcontact >>
rect 7385 14795 7435 14845
<< pdcontact >>
rect 7535 14795 7585 14845
<< pdcontact >>
rect 7685 14795 7735 14845
<< pdcontact >>
rect 7835 14795 7885 14845
<< pdcontact >>
rect 7985 14795 8035 14845
<< pdcontact >>
rect 8135 14795 8185 14845
<< pdcontact >>
rect 8285 14795 8335 14845
<< pdcontact >>
rect 8435 14795 8485 14845
<< pdcontact >>
rect 8585 14795 8635 14845
<< pdcontact >>
rect 8735 14795 8785 14845
<< pdcontact >>
rect 8885 14795 8935 14845
<< pdcontact >>
rect 9035 14795 9085 14845
<< pdcontact >>
rect 9185 14795 9235 14845
<< pdcontact >>
rect 9335 14795 9385 14845
<< pdcontact >>
rect 9485 14795 9535 14845
<< polycontact >>
rect 9755 14825 9805 14875
<< nsubstratencontact >>
rect 9995 14795 10045 14845
<< nsubstratencontact >>
rect 10145 14795 10195 14845
<< psubstratepcontact >>
rect 10535 14795 10585 14845
<< psubstratepcontact >>
rect 10685 14795 10735 14845
<< nsubstratencontact >>
rect 605 14645 655 14695
<< nsubstratencontact >>
rect 755 14645 805 14695
<< polycontact >>
rect 995 14675 1045 14725
<< pdcontact >>
rect 1265 14645 1315 14695
<< pdcontact >>
rect 1415 14645 1465 14695
<< pdcontact >>
rect 1565 14645 1615 14695
<< pdcontact >>
rect 1715 14645 1765 14695
<< pdcontact >>
rect 1865 14645 1915 14695
<< pdcontact >>
rect 2015 14645 2065 14695
<< pdcontact >>
rect 2165 14645 2215 14695
<< pdcontact >>
rect 2315 14645 2365 14695
<< pdcontact >>
rect 2465 14645 2515 14695
<< pdcontact >>
rect 2615 14645 2665 14695
<< pdcontact >>
rect 2765 14645 2815 14695
<< pdcontact >>
rect 2915 14645 2965 14695
<< pdcontact >>
rect 3065 14645 3115 14695
<< pdcontact >>
rect 3215 14645 3265 14695
<< pdcontact >>
rect 3365 14645 3415 14695
<< pdcontact >>
rect 3515 14645 3565 14695
<< pdcontact >>
rect 3665 14645 3715 14695
<< pdcontact >>
rect 3815 14645 3865 14695
<< pdcontact >>
rect 3965 14645 4015 14695
<< pdcontact >>
rect 4115 14645 4165 14695
<< pdcontact >>
rect 4265 14645 4315 14695
<< pdcontact >>
rect 4415 14645 4465 14695
<< pdcontact >>
rect 4565 14645 4615 14695
<< pdcontact >>
rect 4715 14645 4765 14695
<< pdcontact >>
rect 4865 14645 4915 14695
<< polycontact >>
rect 5075 14675 5125 14725
<< nsubstratencontact >>
rect 5315 14645 5365 14695
<< nsubstratencontact >>
rect 5465 14645 5515 14695
<< polycontact >>
rect 5675 14675 5725 14725
<< pdcontact >>
rect 5885 14645 5935 14695
<< pdcontact >>
rect 6035 14645 6085 14695
<< pdcontact >>
rect 6185 14645 6235 14695
<< pdcontact >>
rect 6335 14645 6385 14695
<< pdcontact >>
rect 6485 14645 6535 14695
<< pdcontact >>
rect 6635 14645 6685 14695
<< pdcontact >>
rect 6785 14645 6835 14695
<< pdcontact >>
rect 6935 14645 6985 14695
<< pdcontact >>
rect 7085 14645 7135 14695
<< pdcontact >>
rect 7235 14645 7285 14695
<< pdcontact >>
rect 7385 14645 7435 14695
<< pdcontact >>
rect 7535 14645 7585 14695
<< pdcontact >>
rect 7685 14645 7735 14695
<< pdcontact >>
rect 7835 14645 7885 14695
<< pdcontact >>
rect 7985 14645 8035 14695
<< pdcontact >>
rect 8135 14645 8185 14695
<< pdcontact >>
rect 8285 14645 8335 14695
<< pdcontact >>
rect 8435 14645 8485 14695
<< pdcontact >>
rect 8585 14645 8635 14695
<< pdcontact >>
rect 8735 14645 8785 14695
<< pdcontact >>
rect 8885 14645 8935 14695
<< pdcontact >>
rect 9035 14645 9085 14695
<< pdcontact >>
rect 9185 14645 9235 14695
<< pdcontact >>
rect 9335 14645 9385 14695
<< pdcontact >>
rect 9485 14645 9535 14695
<< polycontact >>
rect 9755 14675 9805 14725
<< nsubstratencontact >>
rect 9995 14645 10045 14695
<< nsubstratencontact >>
rect 10145 14645 10195 14695
<< psubstratepcontact >>
rect 65 14555 115 14605
<< psubstratepcontact >>
rect 215 14555 265 14605
<< nsubstratencontact >>
rect 605 14495 655 14545
<< nsubstratencontact >>
rect 755 14495 805 14545
<< polycontact >>
rect 995 14525 1045 14575
<< pdcontact >>
rect 1265 14495 1315 14545
<< pdcontact >>
rect 1415 14495 1465 14545
<< pdcontact >>
rect 1565 14495 1615 14545
<< pdcontact >>
rect 1715 14495 1765 14545
<< pdcontact >>
rect 1865 14495 1915 14545
<< pdcontact >>
rect 2015 14495 2065 14545
<< pdcontact >>
rect 2165 14495 2215 14545
<< pdcontact >>
rect 2315 14495 2365 14545
<< pdcontact >>
rect 2465 14495 2515 14545
<< pdcontact >>
rect 2615 14495 2665 14545
<< pdcontact >>
rect 2765 14495 2815 14545
<< pdcontact >>
rect 2915 14495 2965 14545
<< pdcontact >>
rect 3065 14495 3115 14545
<< pdcontact >>
rect 3215 14495 3265 14545
<< pdcontact >>
rect 3365 14495 3415 14545
<< pdcontact >>
rect 3515 14495 3565 14545
<< pdcontact >>
rect 3665 14495 3715 14545
<< pdcontact >>
rect 3815 14495 3865 14545
<< pdcontact >>
rect 3965 14495 4015 14545
<< pdcontact >>
rect 4115 14495 4165 14545
<< pdcontact >>
rect 4265 14495 4315 14545
<< pdcontact >>
rect 4415 14495 4465 14545
<< pdcontact >>
rect 4565 14495 4615 14545
<< pdcontact >>
rect 4715 14495 4765 14545
<< pdcontact >>
rect 4865 14495 4915 14545
<< polycontact >>
rect 5075 14525 5125 14575
<< nsubstratencontact >>
rect 5315 14495 5365 14545
<< nsubstratencontact >>
rect 5465 14495 5515 14545
<< polycontact >>
rect 5675 14525 5725 14575
<< pdcontact >>
rect 5885 14495 5935 14545
<< pdcontact >>
rect 6035 14495 6085 14545
<< pdcontact >>
rect 6185 14495 6235 14545
<< pdcontact >>
rect 6335 14495 6385 14545
<< pdcontact >>
rect 6485 14495 6535 14545
<< pdcontact >>
rect 6635 14495 6685 14545
<< pdcontact >>
rect 6785 14495 6835 14545
<< pdcontact >>
rect 6935 14495 6985 14545
<< pdcontact >>
rect 7085 14495 7135 14545
<< pdcontact >>
rect 7235 14495 7285 14545
<< pdcontact >>
rect 7385 14495 7435 14545
<< pdcontact >>
rect 7535 14495 7585 14545
<< pdcontact >>
rect 7685 14495 7735 14545
<< pdcontact >>
rect 7835 14495 7885 14545
<< pdcontact >>
rect 7985 14495 8035 14545
<< pdcontact >>
rect 8135 14495 8185 14545
<< pdcontact >>
rect 8285 14495 8335 14545
<< pdcontact >>
rect 8435 14495 8485 14545
<< pdcontact >>
rect 8585 14495 8635 14545
<< pdcontact >>
rect 8735 14495 8785 14545
<< pdcontact >>
rect 8885 14495 8935 14545
<< pdcontact >>
rect 9035 14495 9085 14545
<< pdcontact >>
rect 9185 14495 9235 14545
<< pdcontact >>
rect 9335 14495 9385 14545
<< pdcontact >>
rect 9485 14495 9535 14545
<< polycontact >>
rect 9755 14525 9805 14575
<< psubstratepcontact >>
rect 10535 14555 10585 14605
<< psubstratepcontact >>
rect 10685 14555 10735 14605
<< nsubstratencontact >>
rect 9995 14495 10045 14545
<< nsubstratencontact >>
rect 10145 14495 10195 14545
<< psubstratepcontact >>
rect 65 14315 115 14365
<< psubstratepcontact >>
rect 215 14315 265 14365
<< nsubstratencontact >>
rect 605 14345 655 14395
<< nsubstratencontact >>
rect 755 14345 805 14395
<< polycontact >>
rect 995 14375 1045 14425
<< polycontact >>
rect 5075 14375 5125 14425
<< nsubstratencontact >>
rect 5315 14345 5365 14395
<< nsubstratencontact >>
rect 5465 14345 5515 14395
<< polycontact >>
rect 5675 14375 5725 14425
<< polycontact >>
rect 9755 14375 9805 14425
<< nsubstratencontact >>
rect 9995 14345 10045 14395
<< nsubstratencontact >>
rect 10145 14345 10195 14395
<< psubstratepcontact >>
rect 10535 14315 10585 14365
<< psubstratepcontact >>
rect 10685 14315 10735 14365
<< pdcontact >>
rect 1235 14195 1285 14245
<< pdcontact >>
rect 1535 14195 1585 14245
<< pdcontact >>
rect 1835 14195 1885 14245
<< pdcontact >>
rect 2135 14195 2185 14245
<< pdcontact >>
rect 2435 14195 2485 14245
<< pdcontact >>
rect 2735 14195 2785 14245
<< pdcontact >>
rect 3035 14195 3085 14245
<< pdcontact >>
rect 3335 14195 3385 14245
<< pdcontact >>
rect 4505 14195 4555 14245
<< pdcontact >>
rect 4805 14195 4855 14245
<< pdcontact >>
rect 5945 14195 5995 14245
<< pdcontact >>
rect 6245 14195 6295 14245
<< pdcontact >>
rect 7415 14195 7465 14245
<< pdcontact >>
rect 7715 14195 7765 14245
<< pdcontact >>
rect 8015 14195 8065 14245
<< pdcontact >>
rect 8315 14195 8365 14245
<< pdcontact >>
rect 8615 14195 8665 14245
<< pdcontact >>
rect 8915 14195 8965 14245
<< pdcontact >>
rect 9215 14195 9265 14245
<< pdcontact >>
rect 9515 14195 9565 14245
<< psubstratepcontact >>
rect 65 14075 115 14125
<< psubstratepcontact >>
rect 215 14075 265 14125
<< pdcontact >>
rect 1235 14045 1285 14095
<< pdcontact >>
rect 1535 14045 1585 14095
<< pdcontact >>
rect 1835 14045 1885 14095
<< pdcontact >>
rect 2135 14045 2185 14095
<< pdcontact >>
rect 2435 14045 2485 14095
<< pdcontact >>
rect 2735 14045 2785 14095
<< pdcontact >>
rect 3035 14045 3085 14095
<< pdcontact >>
rect 3335 14045 3385 14095
<< pdcontact >>
rect 4505 14045 4555 14095
<< pdcontact >>
rect 4805 14045 4855 14095
<< pdcontact >>
rect 5945 14045 5995 14095
<< pdcontact >>
rect 6245 14045 6295 14095
<< pdcontact >>
rect 7415 14045 7465 14095
<< pdcontact >>
rect 7715 14045 7765 14095
<< pdcontact >>
rect 8015 14045 8065 14095
<< pdcontact >>
rect 8315 14045 8365 14095
<< pdcontact >>
rect 8615 14045 8665 14095
<< pdcontact >>
rect 8915 14045 8965 14095
<< pdcontact >>
rect 9215 14045 9265 14095
<< pdcontact >>
rect 9515 14045 9565 14095
<< psubstratepcontact >>
rect 10535 14075 10585 14125
<< psubstratepcontact >>
rect 10685 14075 10735 14125
<< nsubstratencontact >>
rect 1235 13895 1285 13945
<< nsubstratencontact >>
rect 1535 13895 1585 13945
<< nsubstratencontact >>
rect 1835 13895 1885 13945
<< nsubstratencontact >>
rect 2135 13895 2185 13945
<< nsubstratencontact >>
rect 2435 13895 2485 13945
<< nsubstratencontact >>
rect 2735 13895 2785 13945
<< nsubstratencontact >>
rect 3035 13895 3085 13945
<< nsubstratencontact >>
rect 3335 13895 3385 13945
<< nsubstratencontact >>
rect 4505 13895 4555 13945
<< nsubstratencontact >>
rect 4805 13895 4855 13945
<< nsubstratencontact >>
rect 5945 13895 5995 13945
<< nsubstratencontact >>
rect 6245 13895 6295 13945
<< nsubstratencontact >>
rect 7415 13895 7465 13945
<< nsubstratencontact >>
rect 7715 13895 7765 13945
<< nsubstratencontact >>
rect 8015 13895 8065 13945
<< nsubstratencontact >>
rect 8315 13895 8365 13945
<< nsubstratencontact >>
rect 8615 13895 8665 13945
<< nsubstratencontact >>
rect 8915 13895 8965 13945
<< nsubstratencontact >>
rect 9215 13895 9265 13945
<< nsubstratencontact >>
rect 9515 13895 9565 13945
<< psubstratepcontact >>
rect 65 13835 115 13885
<< psubstratepcontact >>
rect 215 13835 265 13885
<< psubstratepcontact >>
rect 10535 13835 10585 13885
<< psubstratepcontact >>
rect 10685 13835 10735 13885
<< psubstratepcontact >>
rect 65 13595 115 13645
<< psubstratepcontact >>
rect 215 13595 265 13645
<< psubstratepcontact >>
rect 10535 13595 10585 13645
<< psubstratepcontact >>
rect 10685 13595 10735 13645
<< psubstratepcontact >>
rect 275 13355 325 13405
<< psubstratepcontact >>
rect 515 13355 565 13405
<< psubstratepcontact >>
rect 755 13355 805 13405
<< psubstratepcontact >>
rect 1235 13355 1285 13405
<< psubstratepcontact >>
rect 1475 13355 1525 13405
<< psubstratepcontact >>
rect 1715 13355 1765 13405
<< psubstratepcontact >>
rect 1955 13355 2005 13405
<< psubstratepcontact >>
rect 2195 13355 2245 13405
<< psubstratepcontact >>
rect 2435 13355 2485 13405
<< psubstratepcontact >>
rect 2675 13355 2725 13405
<< psubstratepcontact >>
rect 2915 13355 2965 13405
<< psubstratepcontact >>
rect 3155 13355 3205 13405
<< psubstratepcontact >>
rect 3395 13355 3445 13405
<< psubstratepcontact >>
rect 4505 13355 4555 13405
<< psubstratepcontact >>
rect 4745 13355 4795 13405
<< psubstratepcontact >>
rect 5435 13355 5485 13405
<< psubstratepcontact >>
rect 5945 13355 5995 13405
<< psubstratepcontact >>
rect 6185 13355 6235 13405
<< psubstratepcontact >>
rect 7355 13355 7405 13405
<< psubstratepcontact >>
rect 7595 13355 7645 13405
<< psubstratepcontact >>
rect 7835 13355 7885 13405
<< psubstratepcontact >>
rect 8075 13355 8125 13405
<< psubstratepcontact >>
rect 8315 13355 8365 13405
<< psubstratepcontact >>
rect 8555 13355 8605 13405
<< psubstratepcontact >>
rect 8795 13355 8845 13405
<< psubstratepcontact >>
rect 9035 13355 9085 13405
<< psubstratepcontact >>
rect 9275 13355 9325 13405
<< psubstratepcontact >>
rect 9515 13355 9565 13405
<< psubstratepcontact >>
rect 9995 13355 10045 13405
<< psubstratepcontact >>
rect 10235 13355 10285 13405
<< psubstratepcontact >>
rect 10475 13355 10525 13405
<< psubstratepcontact >>
rect 275 13205 325 13255
<< psubstratepcontact >>
rect 515 13205 565 13255
<< psubstratepcontact >>
rect 755 13205 805 13255
<< psubstratepcontact >>
rect 1235 13205 1285 13255
<< psubstratepcontact >>
rect 1475 13205 1525 13255
<< psubstratepcontact >>
rect 1715 13205 1765 13255
<< psubstratepcontact >>
rect 1955 13205 2005 13255
<< psubstratepcontact >>
rect 2195 13205 2245 13255
<< psubstratepcontact >>
rect 2435 13205 2485 13255
<< psubstratepcontact >>
rect 2675 13205 2725 13255
<< psubstratepcontact >>
rect 2915 13205 2965 13255
<< psubstratepcontact >>
rect 3155 13205 3205 13255
<< psubstratepcontact >>
rect 3395 13205 3445 13255
<< psubstratepcontact >>
rect 4505 13205 4555 13255
<< psubstratepcontact >>
rect 4745 13205 4795 13255
<< psubstratepcontact >>
rect 5435 13205 5485 13255
<< psubstratepcontact >>
rect 5945 13205 5995 13255
<< psubstratepcontact >>
rect 6185 13205 6235 13255
<< psubstratepcontact >>
rect 7355 13205 7405 13255
<< psubstratepcontact >>
rect 7595 13205 7645 13255
<< psubstratepcontact >>
rect 7835 13205 7885 13255
<< psubstratepcontact >>
rect 8075 13205 8125 13255
<< psubstratepcontact >>
rect 8315 13205 8365 13255
<< psubstratepcontact >>
rect 8555 13205 8605 13255
<< psubstratepcontact >>
rect 8795 13205 8845 13255
<< psubstratepcontact >>
rect 9035 13205 9085 13255
<< psubstratepcontact >>
rect 9275 13205 9325 13255
<< psubstratepcontact >>
rect 9515 13205 9565 13255
<< psubstratepcontact >>
rect 9995 13205 10045 13255
<< psubstratepcontact >>
rect 10235 13205 10285 13255
<< psubstratepcontact >>
rect 10475 13205 10525 13255
<< nsubstratencontact >>
rect 275 12845 325 12895
<< nsubstratencontact >>
rect 515 12845 565 12895
<< nsubstratencontact >>
rect 755 12845 805 12895
<< nsubstratencontact >>
rect 1235 12845 1285 12895
<< nsubstratencontact >>
rect 1475 12845 1525 12895
<< nsubstratencontact >>
rect 1715 12845 1765 12895
<< nsubstratencontact >>
rect 1955 12845 2005 12895
<< nsubstratencontact >>
rect 2195 12845 2245 12895
<< nsubstratencontact >>
rect 2435 12845 2485 12895
<< nsubstratencontact >>
rect 2675 12845 2725 12895
<< nsubstratencontact >>
rect 2915 12845 2965 12895
<< nsubstratencontact >>
rect 3155 12845 3205 12895
<< nsubstratencontact >>
rect 3395 12845 3445 12895
<< nsubstratencontact >>
rect 4505 12845 4555 12895
<< nsubstratencontact >>
rect 4745 12845 4795 12895
<< nsubstratencontact >>
rect 5435 12845 5485 12895
<< nsubstratencontact >>
rect 5945 12845 5995 12895
<< nsubstratencontact >>
rect 6185 12845 6235 12895
<< nsubstratencontact >>
rect 7355 12845 7405 12895
<< nsubstratencontact >>
rect 7595 12845 7645 12895
<< nsubstratencontact >>
rect 7835 12845 7885 12895
<< nsubstratencontact >>
rect 8075 12845 8125 12895
<< nsubstratencontact >>
rect 8315 12845 8365 12895
<< nsubstratencontact >>
rect 8555 12845 8605 12895
<< nsubstratencontact >>
rect 8795 12845 8845 12895
<< nsubstratencontact >>
rect 9035 12845 9085 12895
<< nsubstratencontact >>
rect 9275 12845 9325 12895
<< nsubstratencontact >>
rect 9515 12845 9565 12895
<< nsubstratencontact >>
rect 9995 12845 10045 12895
<< nsubstratencontact >>
rect 10235 12845 10285 12895
<< nsubstratencontact >>
rect 10475 12845 10525 12895
<< nsubstratencontact >>
rect 275 12695 325 12745
<< nsubstratencontact >>
rect 515 12695 565 12745
<< nsubstratencontact >>
rect 755 12695 805 12745
<< nsubstratencontact >>
rect 1235 12695 1285 12745
<< nsubstratencontact >>
rect 1475 12695 1525 12745
<< nsubstratencontact >>
rect 1715 12695 1765 12745
<< nsubstratencontact >>
rect 1955 12695 2005 12745
<< nsubstratencontact >>
rect 2195 12695 2245 12745
<< nsubstratencontact >>
rect 2435 12695 2485 12745
<< nsubstratencontact >>
rect 2675 12695 2725 12745
<< nsubstratencontact >>
rect 2915 12695 2965 12745
<< nsubstratencontact >>
rect 3155 12695 3205 12745
<< nsubstratencontact >>
rect 3395 12695 3445 12745
<< nsubstratencontact >>
rect 4505 12695 4555 12745
<< nsubstratencontact >>
rect 4745 12695 4795 12745
<< nsubstratencontact >>
rect 5435 12695 5485 12745
<< nsubstratencontact >>
rect 5945 12695 5995 12745
<< nsubstratencontact >>
rect 6185 12695 6235 12745
<< nsubstratencontact >>
rect 7355 12695 7405 12745
<< nsubstratencontact >>
rect 7595 12695 7645 12745
<< nsubstratencontact >>
rect 7835 12695 7885 12745
<< nsubstratencontact >>
rect 8075 12695 8125 12745
<< nsubstratencontact >>
rect 8315 12695 8365 12745
<< nsubstratencontact >>
rect 8555 12695 8605 12745
<< nsubstratencontact >>
rect 8795 12695 8845 12745
<< nsubstratencontact >>
rect 9035 12695 9085 12745
<< nsubstratencontact >>
rect 9275 12695 9325 12745
<< nsubstratencontact >>
rect 9515 12695 9565 12745
<< nsubstratencontact >>
rect 9995 12695 10045 12745
<< nsubstratencontact >>
rect 10235 12695 10285 12745
<< nsubstratencontact >>
rect 10475 12695 10525 12745
<< psubstratepcontact >>
rect 275 12005 325 12055
<< psubstratepcontact >>
rect 515 12005 565 12055
<< psubstratepcontact >>
rect 755 12005 805 12055
<< psubstratepcontact >>
rect 995 12005 1045 12055
<< psubstratepcontact >>
rect 1235 12005 1285 12055
<< psubstratepcontact >>
rect 1475 12005 1525 12055
<< psubstratepcontact >>
rect 1715 12005 1765 12055
<< psubstratepcontact >>
rect 1955 12005 2005 12055
<< psubstratepcontact >>
rect 2195 12005 2245 12055
<< psubstratepcontact >>
rect 2435 12005 2485 12055
<< psubstratepcontact >>
rect 2675 12005 2725 12055
<< psubstratepcontact >>
rect 2915 12005 2965 12055
<< psubstratepcontact >>
rect 3155 12005 3205 12055
<< psubstratepcontact >>
rect 3395 12005 3445 12055
<< psubstratepcontact >>
rect 4505 12005 4555 12055
<< psubstratepcontact >>
rect 4745 12005 4795 12055
<< psubstratepcontact >>
rect 5435 12005 5485 12055
<< psubstratepcontact >>
rect 5945 12005 5995 12055
<< psubstratepcontact >>
rect 6185 12005 6235 12055
<< psubstratepcontact >>
rect 7355 12005 7405 12055
<< psubstratepcontact >>
rect 7595 12005 7645 12055
<< psubstratepcontact >>
rect 7835 12005 7885 12055
<< psubstratepcontact >>
rect 8075 12005 8125 12055
<< psubstratepcontact >>
rect 8315 12005 8365 12055
<< psubstratepcontact >>
rect 8555 12005 8605 12055
<< psubstratepcontact >>
rect 8795 12005 8845 12055
<< psubstratepcontact >>
rect 9035 12005 9085 12055
<< psubstratepcontact >>
rect 9275 12005 9325 12055
<< psubstratepcontact >>
rect 9515 12005 9565 12055
<< psubstratepcontact >>
rect 9755 12005 9805 12055
<< psubstratepcontact >>
rect 9995 12005 10045 12055
<< psubstratepcontact >>
rect 10235 12005 10285 12055
<< psubstratepcontact >>
rect 10475 12005 10525 12055
<< psubstratepcontact >>
rect 275 11855 325 11905
<< psubstratepcontact >>
rect 515 11855 565 11905
<< psubstratepcontact >>
rect 755 11855 805 11905
<< psubstratepcontact >>
rect 995 11855 1045 11905
<< psubstratepcontact >>
rect 1235 11855 1285 11905
<< psubstratepcontact >>
rect 1475 11855 1525 11905
<< psubstratepcontact >>
rect 1715 11855 1765 11905
<< psubstratepcontact >>
rect 1955 11855 2005 11905
<< psubstratepcontact >>
rect 2195 11855 2245 11905
<< psubstratepcontact >>
rect 2435 11855 2485 11905
<< psubstratepcontact >>
rect 2675 11855 2725 11905
<< psubstratepcontact >>
rect 2915 11855 2965 11905
<< psubstratepcontact >>
rect 3155 11855 3205 11905
<< psubstratepcontact >>
rect 3395 11855 3445 11905
<< psubstratepcontact >>
rect 4505 11855 4555 11905
<< psubstratepcontact >>
rect 4745 11855 4795 11905
<< psubstratepcontact >>
rect 5435 11855 5485 11905
<< psubstratepcontact >>
rect 5945 11855 5995 11905
<< psubstratepcontact >>
rect 6185 11855 6235 11905
<< psubstratepcontact >>
rect 7355 11855 7405 11905
<< psubstratepcontact >>
rect 7595 11855 7645 11905
<< psubstratepcontact >>
rect 7835 11855 7885 11905
<< psubstratepcontact >>
rect 8075 11855 8125 11905
<< psubstratepcontact >>
rect 8315 11855 8365 11905
<< psubstratepcontact >>
rect 8555 11855 8605 11905
<< psubstratepcontact >>
rect 8795 11855 8845 11905
<< psubstratepcontact >>
rect 9035 11855 9085 11905
<< psubstratepcontact >>
rect 9275 11855 9325 11905
<< psubstratepcontact >>
rect 9515 11855 9565 11905
<< psubstratepcontact >>
rect 9755 11855 9805 11905
<< psubstratepcontact >>
rect 9995 11855 10045 11905
<< psubstratepcontact >>
rect 10235 11855 10285 11905
<< psubstratepcontact >>
rect 10475 11855 10525 11905
<< nsubstratencontact >>
rect 65 11495 115 11545
<< nsubstratencontact >>
rect 275 11495 325 11545
<< nsubstratencontact >>
rect 515 11495 565 11545
<< nsubstratencontact >>
rect 755 11495 805 11545
<< nsubstratencontact >>
rect 995 11495 1045 11545
<< nsubstratencontact >>
rect 1235 11495 1285 11545
<< nsubstratencontact >>
rect 1475 11495 1525 11545
<< nsubstratencontact >>
rect 1715 11495 1765 11545
<< nsubstratencontact >>
rect 1955 11495 2005 11545
<< nsubstratencontact >>
rect 2195 11495 2245 11545
<< nsubstratencontact >>
rect 2435 11495 2485 11545
<< nsubstratencontact >>
rect 2675 11495 2725 11545
<< nsubstratencontact >>
rect 2915 11495 2965 11545
<< nsubstratencontact >>
rect 3155 11495 3205 11545
<< nsubstratencontact >>
rect 3395 11495 3445 11545
<< nsubstratencontact >>
rect 4505 11495 4555 11545
<< nsubstratencontact >>
rect 4745 11495 4795 11545
<< nsubstratencontact >>
rect 4985 11495 5035 11545
<< nsubstratencontact >>
rect 5225 11495 5275 11545
<< nsubstratencontact >>
rect 5435 11495 5485 11545
<< nsubstratencontact >>
rect 5675 11495 5725 11545
<< nsubstratencontact >>
rect 5945 11495 5995 11545
<< nsubstratencontact >>
rect 6185 11495 6235 11545
<< nsubstratencontact >>
rect 7355 11495 7405 11545
<< nsubstratencontact >>
rect 7595 11495 7645 11545
<< nsubstratencontact >>
rect 7835 11495 7885 11545
<< nsubstratencontact >>
rect 8075 11495 8125 11545
<< nsubstratencontact >>
rect 8315 11495 8365 11545
<< nsubstratencontact >>
rect 8555 11495 8605 11545
<< nsubstratencontact >>
rect 8795 11495 8845 11545
<< nsubstratencontact >>
rect 9035 11495 9085 11545
<< nsubstratencontact >>
rect 9275 11495 9325 11545
<< nsubstratencontact >>
rect 9515 11495 9565 11545
<< nsubstratencontact >>
rect 9755 11495 9805 11545
<< nsubstratencontact >>
rect 9995 11495 10045 11545
<< nsubstratencontact >>
rect 10235 11495 10285 11545
<< nsubstratencontact >>
rect 10475 11495 10525 11545
<< nsubstratencontact >>
rect 10715 11495 10765 11545
<< nsubstratencontact >>
rect 65 11345 115 11395
<< nsubstratencontact >>
rect 275 11345 325 11395
<< nsubstratencontact >>
rect 515 11345 565 11395
<< nsubstratencontact >>
rect 755 11345 805 11395
<< nsubstratencontact >>
rect 995 11345 1045 11395
<< nsubstratencontact >>
rect 1235 11345 1285 11395
<< nsubstratencontact >>
rect 1475 11345 1525 11395
<< nsubstratencontact >>
rect 1715 11345 1765 11395
<< nsubstratencontact >>
rect 1955 11345 2005 11395
<< nsubstratencontact >>
rect 2195 11345 2245 11395
<< nsubstratencontact >>
rect 2435 11345 2485 11395
<< nsubstratencontact >>
rect 2675 11345 2725 11395
<< nsubstratencontact >>
rect 2915 11345 2965 11395
<< nsubstratencontact >>
rect 3155 11345 3205 11395
<< nsubstratencontact >>
rect 3395 11345 3445 11395
<< nsubstratencontact >>
rect 4505 11345 4555 11395
<< nsubstratencontact >>
rect 4745 11345 4795 11395
<< nsubstratencontact >>
rect 4985 11345 5035 11395
<< nsubstratencontact >>
rect 5225 11345 5275 11395
<< nsubstratencontact >>
rect 5435 11345 5485 11395
<< nsubstratencontact >>
rect 5675 11345 5725 11395
<< nsubstratencontact >>
rect 5945 11345 5995 11395
<< nsubstratencontact >>
rect 6185 11345 6235 11395
<< nsubstratencontact >>
rect 7355 11345 7405 11395
<< nsubstratencontact >>
rect 7595 11345 7645 11395
<< nsubstratencontact >>
rect 7835 11345 7885 11395
<< nsubstratencontact >>
rect 8075 11345 8125 11395
<< nsubstratencontact >>
rect 8315 11345 8365 11395
<< nsubstratencontact >>
rect 8555 11345 8605 11395
<< nsubstratencontact >>
rect 8795 11345 8845 11395
<< nsubstratencontact >>
rect 9035 11345 9085 11395
<< nsubstratencontact >>
rect 9275 11345 9325 11395
<< nsubstratencontact >>
rect 9515 11345 9565 11395
<< nsubstratencontact >>
rect 9755 11345 9805 11395
<< nsubstratencontact >>
rect 9995 11345 10045 11395
<< nsubstratencontact >>
rect 10235 11345 10285 11395
<< nsubstratencontact >>
rect 10475 11345 10525 11395
<< nsubstratencontact >>
rect 10715 11345 10765 11395
<< nsubstratencontact >>
rect 65 11105 115 11155
<< nsubstratencontact >>
rect 215 11105 265 11155
<< nsubstratencontact >>
rect 10535 11105 10585 11155
<< nsubstratencontact >>
rect 10685 11105 10735 11155
<< nsubstratencontact >>
rect 65 10865 115 10915
<< nsubstratencontact >>
rect 215 10865 265 10915
<< nsubstratencontact >>
rect 10535 10865 10585 10915
<< nsubstratencontact >>
rect 10685 10865 10735 10915
<< psubstratepcontact >>
rect 1235 10805 1285 10855
<< psubstratepcontact >>
rect 1535 10805 1585 10855
<< psubstratepcontact >>
rect 1835 10805 1885 10855
<< psubstratepcontact >>
rect 2135 10805 2185 10855
<< psubstratepcontact >>
rect 2435 10805 2485 10855
<< psubstratepcontact >>
rect 2735 10805 2785 10855
<< psubstratepcontact >>
rect 3035 10805 3085 10855
<< psubstratepcontact >>
rect 3335 10805 3385 10855
<< psubstratepcontact >>
rect 4625 10805 4675 10855
<< psubstratepcontact >>
rect 6125 10805 6175 10855
<< psubstratepcontact >>
rect 7415 10805 7465 10855
<< psubstratepcontact >>
rect 7715 10805 7765 10855
<< psubstratepcontact >>
rect 8015 10805 8065 10855
<< psubstratepcontact >>
rect 8315 10805 8365 10855
<< psubstratepcontact >>
rect 8615 10805 8665 10855
<< psubstratepcontact >>
rect 8915 10805 8965 10855
<< psubstratepcontact >>
rect 9215 10805 9265 10855
<< psubstratepcontact >>
rect 9515 10805 9565 10855
<< nsubstratencontact >>
rect 65 10625 115 10675
<< nsubstratencontact >>
rect 215 10625 265 10675
<< ndcontact >>
rect 1235 10655 1285 10705
<< ndcontact >>
rect 1535 10655 1585 10705
<< ndcontact >>
rect 1835 10655 1885 10705
<< ndcontact >>
rect 2135 10655 2185 10705
<< ndcontact >>
rect 2435 10655 2485 10705
<< ndcontact >>
rect 2735 10655 2785 10705
<< ndcontact >>
rect 3035 10655 3085 10705
<< ndcontact >>
rect 3335 10655 3385 10705
<< ndcontact >>
rect 4625 10655 4675 10705
<< ndcontact >>
rect 6125 10655 6175 10705
<< ndcontact >>
rect 7415 10655 7465 10705
<< ndcontact >>
rect 7715 10655 7765 10705
<< ndcontact >>
rect 8015 10655 8065 10705
<< ndcontact >>
rect 8315 10655 8365 10705
<< ndcontact >>
rect 8615 10655 8665 10705
<< ndcontact >>
rect 8915 10655 8965 10705
<< ndcontact >>
rect 9215 10655 9265 10705
<< ndcontact >>
rect 9515 10655 9565 10705
<< nsubstratencontact >>
rect 10535 10625 10585 10675
<< nsubstratencontact >>
rect 10685 10625 10735 10675
<< ndcontact >>
rect 1235 10505 1285 10555
<< ndcontact >>
rect 1535 10505 1585 10555
<< ndcontact >>
rect 1835 10505 1885 10555
<< ndcontact >>
rect 2135 10505 2185 10555
<< ndcontact >>
rect 2435 10505 2485 10555
<< ndcontact >>
rect 2735 10505 2785 10555
<< ndcontact >>
rect 3035 10505 3085 10555
<< ndcontact >>
rect 3335 10505 3385 10555
<< ndcontact >>
rect 4625 10505 4675 10555
<< ndcontact >>
rect 6125 10505 6175 10555
<< ndcontact >>
rect 7415 10505 7465 10555
<< ndcontact >>
rect 7715 10505 7765 10555
<< ndcontact >>
rect 8015 10505 8065 10555
<< ndcontact >>
rect 8315 10505 8365 10555
<< ndcontact >>
rect 8615 10505 8665 10555
<< ndcontact >>
rect 8915 10505 8965 10555
<< ndcontact >>
rect 9215 10505 9265 10555
<< ndcontact >>
rect 9515 10505 9565 10555
<< nsubstratencontact >>
rect 65 10385 115 10435
<< nsubstratencontact >>
rect 215 10385 265 10435
<< psubstratepcontact >>
rect 605 10355 655 10405
<< psubstratepcontact >>
rect 755 10355 805 10405
<< psubstratepcontact >>
rect 5315 10355 5365 10405
<< psubstratepcontact >>
rect 5465 10355 5515 10405
<< psubstratepcontact >>
rect 9995 10355 10045 10405
<< psubstratepcontact >>
rect 10145 10355 10195 10405
<< nsubstratencontact >>
rect 10535 10385 10585 10435
<< nsubstratencontact >>
rect 10685 10385 10735 10435
<< polycontact >>
rect 995 10265 1045 10315
<< polycontact >>
rect 4865 10265 4915 10315
<< polycontact >>
rect 5885 10265 5935 10315
<< polycontact >>
rect 9755 10265 9805 10315
<< psubstratepcontact >>
rect 605 10205 655 10255
<< psubstratepcontact >>
rect 755 10205 805 10255
<< ndcontact >>
rect 1265 10205 1315 10255
<< ndcontact >>
rect 1415 10205 1465 10255
<< ndcontact >>
rect 1565 10205 1615 10255
<< ndcontact >>
rect 1715 10205 1765 10255
<< ndcontact >>
rect 1865 10205 1915 10255
<< ndcontact >>
rect 2015 10205 2065 10255
<< ndcontact >>
rect 2165 10205 2215 10255
<< ndcontact >>
rect 2315 10205 2365 10255
<< ndcontact >>
rect 2465 10205 2515 10255
<< ndcontact >>
rect 2615 10205 2665 10255
<< ndcontact >>
rect 2765 10205 2815 10255
<< ndcontact >>
rect 2915 10205 2965 10255
<< ndcontact >>
rect 3065 10205 3115 10255
<< ndcontact >>
rect 3215 10205 3265 10255
<< ndcontact >>
rect 3365 10205 3415 10255
<< ndcontact >>
rect 3515 10205 3565 10255
<< ndcontact >>
rect 3665 10205 3715 10255
<< ndcontact >>
rect 3815 10205 3865 10255
<< ndcontact >>
rect 3965 10205 4015 10255
<< ndcontact >>
rect 4115 10205 4165 10255
<< ndcontact >>
rect 4265 10205 4315 10255
<< ndcontact >>
rect 4415 10205 4465 10255
<< ndcontact >>
rect 4565 10205 4615 10255
<< psubstratepcontact >>
rect 5315 10205 5365 10255
<< psubstratepcontact >>
rect 5465 10205 5515 10255
<< ndcontact >>
rect 6185 10205 6235 10255
<< ndcontact >>
rect 6335 10205 6385 10255
<< ndcontact >>
rect 6485 10205 6535 10255
<< ndcontact >>
rect 6635 10205 6685 10255
<< ndcontact >>
rect 6785 10205 6835 10255
<< ndcontact >>
rect 6935 10205 6985 10255
<< ndcontact >>
rect 7085 10205 7135 10255
<< ndcontact >>
rect 7235 10205 7285 10255
<< ndcontact >>
rect 7385 10205 7435 10255
<< ndcontact >>
rect 7535 10205 7585 10255
<< ndcontact >>
rect 7685 10205 7735 10255
<< ndcontact >>
rect 7835 10205 7885 10255
<< ndcontact >>
rect 7985 10205 8035 10255
<< ndcontact >>
rect 8135 10205 8185 10255
<< ndcontact >>
rect 8285 10205 8335 10255
<< ndcontact >>
rect 8435 10205 8485 10255
<< ndcontact >>
rect 8585 10205 8635 10255
<< ndcontact >>
rect 8735 10205 8785 10255
<< ndcontact >>
rect 8885 10205 8935 10255
<< ndcontact >>
rect 9035 10205 9085 10255
<< ndcontact >>
rect 9185 10205 9235 10255
<< ndcontact >>
rect 9335 10205 9385 10255
<< ndcontact >>
rect 9485 10205 9535 10255
<< psubstratepcontact >>
rect 9995 10205 10045 10255
<< psubstratepcontact >>
rect 10145 10205 10195 10255
<< nsubstratencontact >>
rect 65 10145 115 10195
<< nsubstratencontact >>
rect 215 10145 265 10195
<< polycontact >>
rect 995 10115 1045 10165
<< polycontact >>
rect 4865 10115 4915 10165
<< polycontact >>
rect 5885 10115 5935 10165
<< polycontact >>
rect 9755 10115 9805 10165
<< nsubstratencontact >>
rect 10535 10145 10585 10195
<< nsubstratencontact >>
rect 10685 10145 10735 10195
<< psubstratepcontact >>
rect 605 10055 655 10105
<< psubstratepcontact >>
rect 755 10055 805 10105
<< ndcontact >>
rect 1265 10055 1315 10105
<< ndcontact >>
rect 1415 10055 1465 10105
<< ndcontact >>
rect 1565 10055 1615 10105
<< ndcontact >>
rect 1715 10055 1765 10105
<< ndcontact >>
rect 1865 10055 1915 10105
<< ndcontact >>
rect 2015 10055 2065 10105
<< ndcontact >>
rect 2165 10055 2215 10105
<< ndcontact >>
rect 2315 10055 2365 10105
<< ndcontact >>
rect 2465 10055 2515 10105
<< ndcontact >>
rect 2615 10055 2665 10105
<< ndcontact >>
rect 2765 10055 2815 10105
<< ndcontact >>
rect 2915 10055 2965 10105
<< ndcontact >>
rect 3065 10055 3115 10105
<< ndcontact >>
rect 3215 10055 3265 10105
<< ndcontact >>
rect 3365 10055 3415 10105
<< ndcontact >>
rect 3515 10055 3565 10105
<< ndcontact >>
rect 3665 10055 3715 10105
<< ndcontact >>
rect 3815 10055 3865 10105
<< ndcontact >>
rect 3965 10055 4015 10105
<< ndcontact >>
rect 4115 10055 4165 10105
<< ndcontact >>
rect 4265 10055 4315 10105
<< ndcontact >>
rect 4415 10055 4465 10105
<< ndcontact >>
rect 4565 10055 4615 10105
<< psubstratepcontact >>
rect 5315 10055 5365 10105
<< psubstratepcontact >>
rect 5465 10055 5515 10105
<< ndcontact >>
rect 6185 10055 6235 10105
<< ndcontact >>
rect 6335 10055 6385 10105
<< ndcontact >>
rect 6485 10055 6535 10105
<< ndcontact >>
rect 6635 10055 6685 10105
<< ndcontact >>
rect 6785 10055 6835 10105
<< ndcontact >>
rect 6935 10055 6985 10105
<< ndcontact >>
rect 7085 10055 7135 10105
<< ndcontact >>
rect 7235 10055 7285 10105
<< ndcontact >>
rect 7385 10055 7435 10105
<< ndcontact >>
rect 7535 10055 7585 10105
<< ndcontact >>
rect 7685 10055 7735 10105
<< ndcontact >>
rect 7835 10055 7885 10105
<< ndcontact >>
rect 7985 10055 8035 10105
<< ndcontact >>
rect 8135 10055 8185 10105
<< ndcontact >>
rect 8285 10055 8335 10105
<< ndcontact >>
rect 8435 10055 8485 10105
<< ndcontact >>
rect 8585 10055 8635 10105
<< ndcontact >>
rect 8735 10055 8785 10105
<< ndcontact >>
rect 8885 10055 8935 10105
<< ndcontact >>
rect 9035 10055 9085 10105
<< ndcontact >>
rect 9185 10055 9235 10105
<< ndcontact >>
rect 9335 10055 9385 10105
<< ndcontact >>
rect 9485 10055 9535 10105
<< psubstratepcontact >>
rect 9995 10055 10045 10105
<< psubstratepcontact >>
rect 10145 10055 10195 10105
<< polycontact >>
rect 995 9965 1045 10015
<< polycontact >>
rect 4865 9965 4915 10015
<< polycontact >>
rect 5885 9965 5935 10015
<< polycontact >>
rect 9755 9965 9805 10015
<< nsubstratencontact >>
rect 65 9905 115 9955
<< nsubstratencontact >>
rect 215 9905 265 9955
<< psubstratepcontact >>
rect 605 9905 655 9955
<< psubstratepcontact >>
rect 755 9905 805 9955
<< ndcontact >>
rect 1265 9905 1315 9955
<< ndcontact >>
rect 1415 9905 1465 9955
<< ndcontact >>
rect 1565 9905 1615 9955
<< ndcontact >>
rect 1715 9905 1765 9955
<< ndcontact >>
rect 1865 9905 1915 9955
<< ndcontact >>
rect 2015 9905 2065 9955
<< ndcontact >>
rect 2165 9905 2215 9955
<< ndcontact >>
rect 2315 9905 2365 9955
<< ndcontact >>
rect 2465 9905 2515 9955
<< ndcontact >>
rect 2615 9905 2665 9955
<< ndcontact >>
rect 2765 9905 2815 9955
<< ndcontact >>
rect 2915 9905 2965 9955
<< ndcontact >>
rect 3065 9905 3115 9955
<< ndcontact >>
rect 3215 9905 3265 9955
<< ndcontact >>
rect 3365 9905 3415 9955
<< ndcontact >>
rect 3515 9905 3565 9955
<< ndcontact >>
rect 3665 9905 3715 9955
<< ndcontact >>
rect 3815 9905 3865 9955
<< ndcontact >>
rect 3965 9905 4015 9955
<< ndcontact >>
rect 4115 9905 4165 9955
<< ndcontact >>
rect 4265 9905 4315 9955
<< ndcontact >>
rect 4415 9905 4465 9955
<< ndcontact >>
rect 4565 9905 4615 9955
<< psubstratepcontact >>
rect 5315 9905 5365 9955
<< psubstratepcontact >>
rect 5465 9905 5515 9955
<< ndcontact >>
rect 6185 9905 6235 9955
<< ndcontact >>
rect 6335 9905 6385 9955
<< ndcontact >>
rect 6485 9905 6535 9955
<< ndcontact >>
rect 6635 9905 6685 9955
<< ndcontact >>
rect 6785 9905 6835 9955
<< ndcontact >>
rect 6935 9905 6985 9955
<< ndcontact >>
rect 7085 9905 7135 9955
<< ndcontact >>
rect 7235 9905 7285 9955
<< ndcontact >>
rect 7385 9905 7435 9955
<< ndcontact >>
rect 7535 9905 7585 9955
<< ndcontact >>
rect 7685 9905 7735 9955
<< ndcontact >>
rect 7835 9905 7885 9955
<< ndcontact >>
rect 7985 9905 8035 9955
<< ndcontact >>
rect 8135 9905 8185 9955
<< ndcontact >>
rect 8285 9905 8335 9955
<< ndcontact >>
rect 8435 9905 8485 9955
<< ndcontact >>
rect 8585 9905 8635 9955
<< ndcontact >>
rect 8735 9905 8785 9955
<< ndcontact >>
rect 8885 9905 8935 9955
<< ndcontact >>
rect 9035 9905 9085 9955
<< ndcontact >>
rect 9185 9905 9235 9955
<< ndcontact >>
rect 9335 9905 9385 9955
<< ndcontact >>
rect 9485 9905 9535 9955
<< psubstratepcontact >>
rect 9995 9905 10045 9955
<< psubstratepcontact >>
rect 10145 9905 10195 9955
<< nsubstratencontact >>
rect 10535 9905 10585 9955
<< nsubstratencontact >>
rect 10685 9905 10735 9955
<< polycontact >>
rect 995 9815 1045 9865
<< polycontact >>
rect 4865 9815 4915 9865
<< polycontact >>
rect 5885 9815 5935 9865
<< polycontact >>
rect 9755 9815 9805 9865
<< psubstratepcontact >>
rect 605 9755 655 9805
<< psubstratepcontact >>
rect 755 9755 805 9805
<< ndcontact >>
rect 1265 9755 1315 9805
<< ndcontact >>
rect 1415 9755 1465 9805
<< ndcontact >>
rect 1565 9755 1615 9805
<< ndcontact >>
rect 1715 9755 1765 9805
<< ndcontact >>
rect 1865 9755 1915 9805
<< ndcontact >>
rect 2015 9755 2065 9805
<< ndcontact >>
rect 2165 9755 2215 9805
<< ndcontact >>
rect 2315 9755 2365 9805
<< ndcontact >>
rect 2465 9755 2515 9805
<< ndcontact >>
rect 2615 9755 2665 9805
<< ndcontact >>
rect 2765 9755 2815 9805
<< ndcontact >>
rect 2915 9755 2965 9805
<< ndcontact >>
rect 3065 9755 3115 9805
<< ndcontact >>
rect 3215 9755 3265 9805
<< ndcontact >>
rect 3365 9755 3415 9805
<< ndcontact >>
rect 3515 9755 3565 9805
<< ndcontact >>
rect 3665 9755 3715 9805
<< ndcontact >>
rect 3815 9755 3865 9805
<< ndcontact >>
rect 3965 9755 4015 9805
<< ndcontact >>
rect 4115 9755 4165 9805
<< ndcontact >>
rect 4265 9755 4315 9805
<< ndcontact >>
rect 4415 9755 4465 9805
<< ndcontact >>
rect 4565 9755 4615 9805
<< psubstratepcontact >>
rect 5315 9755 5365 9805
<< psubstratepcontact >>
rect 5465 9755 5515 9805
<< ndcontact >>
rect 6185 9755 6235 9805
<< ndcontact >>
rect 6335 9755 6385 9805
<< ndcontact >>
rect 6485 9755 6535 9805
<< ndcontact >>
rect 6635 9755 6685 9805
<< ndcontact >>
rect 6785 9755 6835 9805
<< ndcontact >>
rect 6935 9755 6985 9805
<< ndcontact >>
rect 7085 9755 7135 9805
<< ndcontact >>
rect 7235 9755 7285 9805
<< ndcontact >>
rect 7385 9755 7435 9805
<< ndcontact >>
rect 7535 9755 7585 9805
<< ndcontact >>
rect 7685 9755 7735 9805
<< ndcontact >>
rect 7835 9755 7885 9805
<< ndcontact >>
rect 7985 9755 8035 9805
<< ndcontact >>
rect 8135 9755 8185 9805
<< ndcontact >>
rect 8285 9755 8335 9805
<< ndcontact >>
rect 8435 9755 8485 9805
<< ndcontact >>
rect 8585 9755 8635 9805
<< ndcontact >>
rect 8735 9755 8785 9805
<< ndcontact >>
rect 8885 9755 8935 9805
<< ndcontact >>
rect 9035 9755 9085 9805
<< ndcontact >>
rect 9185 9755 9235 9805
<< ndcontact >>
rect 9335 9755 9385 9805
<< ndcontact >>
rect 9485 9755 9535 9805
<< psubstratepcontact >>
rect 9995 9755 10045 9805
<< psubstratepcontact >>
rect 10145 9755 10195 9805
<< nsubstratencontact >>
rect 65 9665 115 9715
<< nsubstratencontact >>
rect 215 9665 265 9715
<< polycontact >>
rect 995 9665 1045 9715
<< polycontact >>
rect 4865 9665 4915 9715
<< polycontact >>
rect 5885 9665 5935 9715
<< polycontact >>
rect 9755 9665 9805 9715
<< nsubstratencontact >>
rect 10535 9665 10585 9715
<< nsubstratencontact >>
rect 10685 9665 10735 9715
<< psubstratepcontact >>
rect 605 9605 655 9655
<< psubstratepcontact >>
rect 755 9605 805 9655
<< ndcontact >>
rect 1265 9605 1315 9655
<< ndcontact >>
rect 1415 9605 1465 9655
<< ndcontact >>
rect 1565 9605 1615 9655
<< ndcontact >>
rect 1715 9605 1765 9655
<< ndcontact >>
rect 1865 9605 1915 9655
<< ndcontact >>
rect 2015 9605 2065 9655
<< ndcontact >>
rect 2165 9605 2215 9655
<< ndcontact >>
rect 2315 9605 2365 9655
<< ndcontact >>
rect 2465 9605 2515 9655
<< ndcontact >>
rect 2615 9605 2665 9655
<< ndcontact >>
rect 2765 9605 2815 9655
<< ndcontact >>
rect 2915 9605 2965 9655
<< ndcontact >>
rect 3065 9605 3115 9655
<< ndcontact >>
rect 3215 9605 3265 9655
<< ndcontact >>
rect 3365 9605 3415 9655
<< ndcontact >>
rect 3515 9605 3565 9655
<< ndcontact >>
rect 3665 9605 3715 9655
<< ndcontact >>
rect 3815 9605 3865 9655
<< ndcontact >>
rect 3965 9605 4015 9655
<< ndcontact >>
rect 4115 9605 4165 9655
<< ndcontact >>
rect 4265 9605 4315 9655
<< ndcontact >>
rect 4415 9605 4465 9655
<< ndcontact >>
rect 4565 9605 4615 9655
<< psubstratepcontact >>
rect 5315 9605 5365 9655
<< psubstratepcontact >>
rect 5465 9605 5515 9655
<< ndcontact >>
rect 6185 9605 6235 9655
<< ndcontact >>
rect 6335 9605 6385 9655
<< ndcontact >>
rect 6485 9605 6535 9655
<< ndcontact >>
rect 6635 9605 6685 9655
<< ndcontact >>
rect 6785 9605 6835 9655
<< ndcontact >>
rect 6935 9605 6985 9655
<< ndcontact >>
rect 7085 9605 7135 9655
<< ndcontact >>
rect 7235 9605 7285 9655
<< ndcontact >>
rect 7385 9605 7435 9655
<< ndcontact >>
rect 7535 9605 7585 9655
<< ndcontact >>
rect 7685 9605 7735 9655
<< ndcontact >>
rect 7835 9605 7885 9655
<< ndcontact >>
rect 7985 9605 8035 9655
<< ndcontact >>
rect 8135 9605 8185 9655
<< ndcontact >>
rect 8285 9605 8335 9655
<< ndcontact >>
rect 8435 9605 8485 9655
<< ndcontact >>
rect 8585 9605 8635 9655
<< ndcontact >>
rect 8735 9605 8785 9655
<< ndcontact >>
rect 8885 9605 8935 9655
<< ndcontact >>
rect 9035 9605 9085 9655
<< ndcontact >>
rect 9185 9605 9235 9655
<< ndcontact >>
rect 9335 9605 9385 9655
<< ndcontact >>
rect 9485 9605 9535 9655
<< psubstratepcontact >>
rect 9995 9605 10045 9655
<< psubstratepcontact >>
rect 10145 9605 10195 9655
<< polycontact >>
rect 995 9515 1045 9565
<< polycontact >>
rect 4865 9515 4915 9565
<< polycontact >>
rect 5885 9515 5935 9565
<< polycontact >>
rect 9755 9515 9805 9565
<< nsubstratencontact >>
rect 65 9425 115 9475
<< nsubstratencontact >>
rect 215 9425 265 9475
<< psubstratepcontact >>
rect 605 9455 655 9505
<< psubstratepcontact >>
rect 755 9455 805 9505
<< ndcontact >>
rect 1265 9455 1315 9505
<< ndcontact >>
rect 1415 9455 1465 9505
<< ndcontact >>
rect 1565 9455 1615 9505
<< ndcontact >>
rect 1715 9455 1765 9505
<< ndcontact >>
rect 1865 9455 1915 9505
<< ndcontact >>
rect 2015 9455 2065 9505
<< ndcontact >>
rect 2165 9455 2215 9505
<< ndcontact >>
rect 2315 9455 2365 9505
<< ndcontact >>
rect 2465 9455 2515 9505
<< ndcontact >>
rect 2615 9455 2665 9505
<< ndcontact >>
rect 2765 9455 2815 9505
<< ndcontact >>
rect 2915 9455 2965 9505
<< ndcontact >>
rect 3065 9455 3115 9505
<< ndcontact >>
rect 3215 9455 3265 9505
<< ndcontact >>
rect 3365 9455 3415 9505
<< ndcontact >>
rect 3515 9455 3565 9505
<< ndcontact >>
rect 3665 9455 3715 9505
<< ndcontact >>
rect 3815 9455 3865 9505
<< ndcontact >>
rect 3965 9455 4015 9505
<< ndcontact >>
rect 4115 9455 4165 9505
<< ndcontact >>
rect 4265 9455 4315 9505
<< ndcontact >>
rect 4415 9455 4465 9505
<< ndcontact >>
rect 4565 9455 4615 9505
<< psubstratepcontact >>
rect 5315 9455 5365 9505
<< psubstratepcontact >>
rect 5465 9455 5515 9505
<< ndcontact >>
rect 6185 9455 6235 9505
<< ndcontact >>
rect 6335 9455 6385 9505
<< ndcontact >>
rect 6485 9455 6535 9505
<< ndcontact >>
rect 6635 9455 6685 9505
<< ndcontact >>
rect 6785 9455 6835 9505
<< ndcontact >>
rect 6935 9455 6985 9505
<< ndcontact >>
rect 7085 9455 7135 9505
<< ndcontact >>
rect 7235 9455 7285 9505
<< ndcontact >>
rect 7385 9455 7435 9505
<< ndcontact >>
rect 7535 9455 7585 9505
<< ndcontact >>
rect 7685 9455 7735 9505
<< ndcontact >>
rect 7835 9455 7885 9505
<< ndcontact >>
rect 7985 9455 8035 9505
<< ndcontact >>
rect 8135 9455 8185 9505
<< ndcontact >>
rect 8285 9455 8335 9505
<< ndcontact >>
rect 8435 9455 8485 9505
<< ndcontact >>
rect 8585 9455 8635 9505
<< ndcontact >>
rect 8735 9455 8785 9505
<< ndcontact >>
rect 8885 9455 8935 9505
<< ndcontact >>
rect 9035 9455 9085 9505
<< ndcontact >>
rect 9185 9455 9235 9505
<< ndcontact >>
rect 9335 9455 9385 9505
<< ndcontact >>
rect 9485 9455 9535 9505
<< psubstratepcontact >>
rect 9995 9455 10045 9505
<< psubstratepcontact >>
rect 10145 9455 10195 9505
<< nsubstratencontact >>
rect 10535 9425 10585 9475
<< nsubstratencontact >>
rect 10685 9425 10735 9475
<< polycontact >>
rect 995 9365 1045 9415
<< polycontact >>
rect 4865 9365 4915 9415
<< polycontact >>
rect 5885 9365 5935 9415
<< polycontact >>
rect 9755 9365 9805 9415
<< psubstratepcontact >>
rect 605 9305 655 9355
<< psubstratepcontact >>
rect 755 9305 805 9355
<< ndcontact >>
rect 1265 9305 1315 9355
<< ndcontact >>
rect 1415 9305 1465 9355
<< ndcontact >>
rect 1565 9305 1615 9355
<< ndcontact >>
rect 1715 9305 1765 9355
<< ndcontact >>
rect 1865 9305 1915 9355
<< ndcontact >>
rect 2015 9305 2065 9355
<< ndcontact >>
rect 2165 9305 2215 9355
<< ndcontact >>
rect 2315 9305 2365 9355
<< ndcontact >>
rect 2465 9305 2515 9355
<< ndcontact >>
rect 2615 9305 2665 9355
<< ndcontact >>
rect 2765 9305 2815 9355
<< ndcontact >>
rect 2915 9305 2965 9355
<< ndcontact >>
rect 3065 9305 3115 9355
<< ndcontact >>
rect 3215 9305 3265 9355
<< ndcontact >>
rect 3365 9305 3415 9355
<< ndcontact >>
rect 3515 9305 3565 9355
<< ndcontact >>
rect 3665 9305 3715 9355
<< ndcontact >>
rect 3815 9305 3865 9355
<< ndcontact >>
rect 3965 9305 4015 9355
<< ndcontact >>
rect 4115 9305 4165 9355
<< ndcontact >>
rect 4265 9305 4315 9355
<< ndcontact >>
rect 4415 9305 4465 9355
<< ndcontact >>
rect 4565 9305 4615 9355
<< psubstratepcontact >>
rect 5315 9305 5365 9355
<< psubstratepcontact >>
rect 5465 9305 5515 9355
<< ndcontact >>
rect 6185 9305 6235 9355
<< ndcontact >>
rect 6335 9305 6385 9355
<< ndcontact >>
rect 6485 9305 6535 9355
<< ndcontact >>
rect 6635 9305 6685 9355
<< ndcontact >>
rect 6785 9305 6835 9355
<< ndcontact >>
rect 6935 9305 6985 9355
<< ndcontact >>
rect 7085 9305 7135 9355
<< ndcontact >>
rect 7235 9305 7285 9355
<< ndcontact >>
rect 7385 9305 7435 9355
<< ndcontact >>
rect 7535 9305 7585 9355
<< ndcontact >>
rect 7685 9305 7735 9355
<< ndcontact >>
rect 7835 9305 7885 9355
<< ndcontact >>
rect 7985 9305 8035 9355
<< ndcontact >>
rect 8135 9305 8185 9355
<< ndcontact >>
rect 8285 9305 8335 9355
<< ndcontact >>
rect 8435 9305 8485 9355
<< ndcontact >>
rect 8585 9305 8635 9355
<< ndcontact >>
rect 8735 9305 8785 9355
<< ndcontact >>
rect 8885 9305 8935 9355
<< ndcontact >>
rect 9035 9305 9085 9355
<< ndcontact >>
rect 9185 9305 9235 9355
<< ndcontact >>
rect 9335 9305 9385 9355
<< ndcontact >>
rect 9485 9305 9535 9355
<< psubstratepcontact >>
rect 9995 9305 10045 9355
<< psubstratepcontact >>
rect 10145 9305 10195 9355
<< nsubstratencontact >>
rect 65 9185 115 9235
<< nsubstratencontact >>
rect 215 9185 265 9235
<< polycontact >>
rect 995 9215 1045 9265
<< polycontact >>
rect 4865 9215 4915 9265
<< polycontact >>
rect 5885 9215 5935 9265
<< polycontact >>
rect 9755 9215 9805 9265
<< psubstratepcontact >>
rect 605 9155 655 9205
<< psubstratepcontact >>
rect 755 9155 805 9205
<< ndcontact >>
rect 1265 9155 1315 9205
<< ndcontact >>
rect 1415 9155 1465 9205
<< ndcontact >>
rect 1565 9155 1615 9205
<< ndcontact >>
rect 1715 9155 1765 9205
<< ndcontact >>
rect 1865 9155 1915 9205
<< ndcontact >>
rect 2015 9155 2065 9205
<< ndcontact >>
rect 2165 9155 2215 9205
<< ndcontact >>
rect 2315 9155 2365 9205
<< ndcontact >>
rect 2465 9155 2515 9205
<< ndcontact >>
rect 2615 9155 2665 9205
<< ndcontact >>
rect 2765 9155 2815 9205
<< ndcontact >>
rect 2915 9155 2965 9205
<< ndcontact >>
rect 3065 9155 3115 9205
<< ndcontact >>
rect 3215 9155 3265 9205
<< ndcontact >>
rect 3365 9155 3415 9205
<< ndcontact >>
rect 3515 9155 3565 9205
<< ndcontact >>
rect 3665 9155 3715 9205
<< ndcontact >>
rect 3815 9155 3865 9205
<< ndcontact >>
rect 3965 9155 4015 9205
<< ndcontact >>
rect 4115 9155 4165 9205
<< ndcontact >>
rect 4265 9155 4315 9205
<< ndcontact >>
rect 4415 9155 4465 9205
<< ndcontact >>
rect 4565 9155 4615 9205
<< psubstratepcontact >>
rect 5315 9155 5365 9205
<< psubstratepcontact >>
rect 5465 9155 5515 9205
<< ndcontact >>
rect 6185 9155 6235 9205
<< ndcontact >>
rect 6335 9155 6385 9205
<< ndcontact >>
rect 6485 9155 6535 9205
<< ndcontact >>
rect 6635 9155 6685 9205
<< ndcontact >>
rect 6785 9155 6835 9205
<< ndcontact >>
rect 6935 9155 6985 9205
<< ndcontact >>
rect 7085 9155 7135 9205
<< ndcontact >>
rect 7235 9155 7285 9205
<< ndcontact >>
rect 7385 9155 7435 9205
<< ndcontact >>
rect 7535 9155 7585 9205
<< ndcontact >>
rect 7685 9155 7735 9205
<< ndcontact >>
rect 7835 9155 7885 9205
<< ndcontact >>
rect 7985 9155 8035 9205
<< ndcontact >>
rect 8135 9155 8185 9205
<< ndcontact >>
rect 8285 9155 8335 9205
<< ndcontact >>
rect 8435 9155 8485 9205
<< ndcontact >>
rect 8585 9155 8635 9205
<< ndcontact >>
rect 8735 9155 8785 9205
<< ndcontact >>
rect 8885 9155 8935 9205
<< ndcontact >>
rect 9035 9155 9085 9205
<< ndcontact >>
rect 9185 9155 9235 9205
<< ndcontact >>
rect 9335 9155 9385 9205
<< ndcontact >>
rect 9485 9155 9535 9205
<< psubstratepcontact >>
rect 9995 9155 10045 9205
<< psubstratepcontact >>
rect 10145 9155 10195 9205
<< nsubstratencontact >>
rect 10535 9185 10585 9235
<< nsubstratencontact >>
rect 10685 9185 10735 9235
<< polycontact >>
rect 995 9065 1045 9115
<< polycontact >>
rect 4865 9065 4915 9115
<< polycontact >>
rect 5885 9065 5935 9115
<< polycontact >>
rect 9755 9065 9805 9115
<< psubstratepcontact >>
rect 605 9005 655 9055
<< psubstratepcontact >>
rect 755 9005 805 9055
<< psubstratepcontact >>
rect 5315 9005 5365 9055
<< psubstratepcontact >>
rect 5465 9005 5515 9055
<< psubstratepcontact >>
rect 9995 9005 10045 9055
<< psubstratepcontact >>
rect 10145 9005 10195 9055
<< nsubstratencontact >>
rect 65 8945 115 8995
<< nsubstratencontact >>
rect 215 8945 265 8995
<< polycontact >>
rect 995 8915 1045 8965
<< polycontact >>
rect 4865 8915 4915 8965
<< polycontact >>
rect 5885 8915 5935 8965
<< polycontact >>
rect 9755 8915 9805 8965
<< nsubstratencontact >>
rect 10535 8945 10585 8995
<< nsubstratencontact >>
rect 10685 8945 10735 8995
<< ndcontact >>
rect 1235 8855 1285 8905
<< ndcontact >>
rect 1535 8855 1585 8905
<< ndcontact >>
rect 1835 8855 1885 8905
<< ndcontact >>
rect 2135 8855 2185 8905
<< ndcontact >>
rect 2435 8855 2485 8905
<< ndcontact >>
rect 2735 8855 2785 8905
<< ndcontact >>
rect 3035 8855 3085 8905
<< ndcontact >>
rect 3335 8855 3385 8905
<< ndcontact >>
rect 4625 8855 4675 8905
<< ndcontact >>
rect 6125 8855 6175 8905
<< ndcontact >>
rect 7415 8855 7465 8905
<< ndcontact >>
rect 7715 8855 7765 8905
<< ndcontact >>
rect 8015 8855 8065 8905
<< ndcontact >>
rect 8315 8855 8365 8905
<< ndcontact >>
rect 8615 8855 8665 8905
<< ndcontact >>
rect 8915 8855 8965 8905
<< ndcontact >>
rect 9215 8855 9265 8905
<< ndcontact >>
rect 9515 8855 9565 8905
<< polycontact >>
rect 995 8765 1045 8815
<< polycontact >>
rect 4865 8765 4915 8815
<< polycontact >>
rect 5885 8765 5935 8815
<< polycontact >>
rect 9755 8765 9805 8815
<< nsubstratencontact >>
rect 65 8705 115 8755
<< nsubstratencontact >>
rect 215 8705 265 8755
<< ndcontact >>
rect 1235 8705 1285 8755
<< ndcontact >>
rect 1535 8705 1585 8755
<< ndcontact >>
rect 1835 8705 1885 8755
<< ndcontact >>
rect 2135 8705 2185 8755
<< ndcontact >>
rect 2435 8705 2485 8755
<< ndcontact >>
rect 2735 8705 2785 8755
<< ndcontact >>
rect 3035 8705 3085 8755
<< ndcontact >>
rect 3335 8705 3385 8755
<< ndcontact >>
rect 4625 8705 4675 8755
<< ndcontact >>
rect 6125 8705 6175 8755
<< ndcontact >>
rect 7415 8705 7465 8755
<< ndcontact >>
rect 7715 8705 7765 8755
<< ndcontact >>
rect 8015 8705 8065 8755
<< ndcontact >>
rect 8315 8705 8365 8755
<< ndcontact >>
rect 8615 8705 8665 8755
<< ndcontact >>
rect 8915 8705 8965 8755
<< ndcontact >>
rect 9215 8705 9265 8755
<< ndcontact >>
rect 9515 8705 9565 8755
<< nsubstratencontact >>
rect 10535 8705 10585 8755
<< nsubstratencontact >>
rect 10685 8705 10735 8755
<< polycontact >>
rect 995 8615 1045 8665
<< polycontact >>
rect 4865 8615 4915 8665
<< polycontact >>
rect 5885 8615 5935 8665
<< polycontact >>
rect 9755 8615 9805 8665
<< ndcontact >>
rect 1235 8555 1285 8605
<< ndcontact >>
rect 1535 8555 1585 8605
<< ndcontact >>
rect 1835 8555 1885 8605
<< ndcontact >>
rect 2135 8555 2185 8605
<< ndcontact >>
rect 2435 8555 2485 8605
<< ndcontact >>
rect 2735 8555 2785 8605
<< ndcontact >>
rect 3035 8555 3085 8605
<< ndcontact >>
rect 3335 8555 3385 8605
<< ndcontact >>
rect 4625 8555 4675 8605
<< ndcontact >>
rect 6125 8555 6175 8605
<< ndcontact >>
rect 7415 8555 7465 8605
<< ndcontact >>
rect 7715 8555 7765 8605
<< ndcontact >>
rect 8015 8555 8065 8605
<< ndcontact >>
rect 8315 8555 8365 8605
<< ndcontact >>
rect 8615 8555 8665 8605
<< ndcontact >>
rect 8915 8555 8965 8605
<< ndcontact >>
rect 9215 8555 9265 8605
<< ndcontact >>
rect 9515 8555 9565 8605
<< nsubstratencontact >>
rect 65 8465 115 8515
<< nsubstratencontact >>
rect 215 8465 265 8515
<< polycontact >>
rect 995 8465 1045 8515
<< polycontact >>
rect 4865 8465 4915 8515
<< polycontact >>
rect 5885 8465 5935 8515
<< polycontact >>
rect 9755 8465 9805 8515
<< nsubstratencontact >>
rect 10535 8465 10585 8515
<< nsubstratencontact >>
rect 10685 8465 10735 8515
<< psubstratepcontact >>
rect 605 8405 655 8455
<< psubstratepcontact >>
rect 755 8405 805 8455
<< psubstratepcontact >>
rect 5315 8405 5365 8455
<< psubstratepcontact >>
rect 5465 8405 5515 8455
<< psubstratepcontact >>
rect 9995 8405 10045 8455
<< psubstratepcontact >>
rect 10145 8405 10195 8455
<< polycontact >>
rect 995 8315 1045 8365
<< polycontact >>
rect 4865 8315 4915 8365
<< polycontact >>
rect 5885 8315 5935 8365
<< polycontact >>
rect 9755 8315 9805 8365
<< nsubstratencontact >>
rect 65 8225 115 8275
<< nsubstratencontact >>
rect 215 8225 265 8275
<< psubstratepcontact >>
rect 605 8255 655 8305
<< psubstratepcontact >>
rect 755 8255 805 8305
<< ndcontact >>
rect 1265 8255 1315 8305
<< ndcontact >>
rect 1415 8255 1465 8305
<< ndcontact >>
rect 1565 8255 1615 8305
<< ndcontact >>
rect 1715 8255 1765 8305
<< ndcontact >>
rect 1865 8255 1915 8305
<< ndcontact >>
rect 2015 8255 2065 8305
<< ndcontact >>
rect 2165 8255 2215 8305
<< ndcontact >>
rect 2315 8255 2365 8305
<< ndcontact >>
rect 2465 8255 2515 8305
<< ndcontact >>
rect 2615 8255 2665 8305
<< ndcontact >>
rect 2765 8255 2815 8305
<< ndcontact >>
rect 2915 8255 2965 8305
<< ndcontact >>
rect 3065 8255 3115 8305
<< ndcontact >>
rect 3215 8255 3265 8305
<< ndcontact >>
rect 3365 8255 3415 8305
<< ndcontact >>
rect 3515 8255 3565 8305
<< ndcontact >>
rect 3665 8255 3715 8305
<< ndcontact >>
rect 3815 8255 3865 8305
<< ndcontact >>
rect 3965 8255 4015 8305
<< ndcontact >>
rect 4115 8255 4165 8305
<< ndcontact >>
rect 4265 8255 4315 8305
<< ndcontact >>
rect 4415 8255 4465 8305
<< ndcontact >>
rect 4565 8255 4615 8305
<< psubstratepcontact >>
rect 5315 8255 5365 8305
<< psubstratepcontact >>
rect 5465 8255 5515 8305
<< ndcontact >>
rect 6185 8255 6235 8305
<< ndcontact >>
rect 6335 8255 6385 8305
<< ndcontact >>
rect 6485 8255 6535 8305
<< ndcontact >>
rect 6635 8255 6685 8305
<< ndcontact >>
rect 6785 8255 6835 8305
<< ndcontact >>
rect 6935 8255 6985 8305
<< ndcontact >>
rect 7085 8255 7135 8305
<< ndcontact >>
rect 7235 8255 7285 8305
<< ndcontact >>
rect 7385 8255 7435 8305
<< ndcontact >>
rect 7535 8255 7585 8305
<< ndcontact >>
rect 7685 8255 7735 8305
<< ndcontact >>
rect 7835 8255 7885 8305
<< ndcontact >>
rect 7985 8255 8035 8305
<< ndcontact >>
rect 8135 8255 8185 8305
<< ndcontact >>
rect 8285 8255 8335 8305
<< ndcontact >>
rect 8435 8255 8485 8305
<< ndcontact >>
rect 8585 8255 8635 8305
<< ndcontact >>
rect 8735 8255 8785 8305
<< ndcontact >>
rect 8885 8255 8935 8305
<< ndcontact >>
rect 9035 8255 9085 8305
<< ndcontact >>
rect 9185 8255 9235 8305
<< ndcontact >>
rect 9335 8255 9385 8305
<< ndcontact >>
rect 9485 8255 9535 8305
<< psubstratepcontact >>
rect 9995 8255 10045 8305
<< psubstratepcontact >>
rect 10145 8255 10195 8305
<< nsubstratencontact >>
rect 10535 8225 10585 8275
<< nsubstratencontact >>
rect 10685 8225 10735 8275
<< polycontact >>
rect 995 8165 1045 8215
<< polycontact >>
rect 4865 8165 4915 8215
<< polycontact >>
rect 5885 8165 5935 8215
<< polycontact >>
rect 9755 8165 9805 8215
<< psubstratepcontact >>
rect 605 8105 655 8155
<< psubstratepcontact >>
rect 755 8105 805 8155
<< ndcontact >>
rect 1265 8105 1315 8155
<< ndcontact >>
rect 1415 8105 1465 8155
<< ndcontact >>
rect 1565 8105 1615 8155
<< ndcontact >>
rect 1715 8105 1765 8155
<< ndcontact >>
rect 1865 8105 1915 8155
<< ndcontact >>
rect 2015 8105 2065 8155
<< ndcontact >>
rect 2165 8105 2215 8155
<< ndcontact >>
rect 2315 8105 2365 8155
<< ndcontact >>
rect 2465 8105 2515 8155
<< ndcontact >>
rect 2615 8105 2665 8155
<< ndcontact >>
rect 2765 8105 2815 8155
<< ndcontact >>
rect 2915 8105 2965 8155
<< ndcontact >>
rect 3065 8105 3115 8155
<< ndcontact >>
rect 3215 8105 3265 8155
<< ndcontact >>
rect 3365 8105 3415 8155
<< ndcontact >>
rect 3515 8105 3565 8155
<< ndcontact >>
rect 3665 8105 3715 8155
<< ndcontact >>
rect 3815 8105 3865 8155
<< ndcontact >>
rect 3965 8105 4015 8155
<< ndcontact >>
rect 4115 8105 4165 8155
<< ndcontact >>
rect 4265 8105 4315 8155
<< ndcontact >>
rect 4415 8105 4465 8155
<< ndcontact >>
rect 4565 8105 4615 8155
<< psubstratepcontact >>
rect 5315 8105 5365 8155
<< psubstratepcontact >>
rect 5465 8105 5515 8155
<< ndcontact >>
rect 6185 8105 6235 8155
<< ndcontact >>
rect 6335 8105 6385 8155
<< ndcontact >>
rect 6485 8105 6535 8155
<< ndcontact >>
rect 6635 8105 6685 8155
<< ndcontact >>
rect 6785 8105 6835 8155
<< ndcontact >>
rect 6935 8105 6985 8155
<< ndcontact >>
rect 7085 8105 7135 8155
<< ndcontact >>
rect 7235 8105 7285 8155
<< ndcontact >>
rect 7385 8105 7435 8155
<< ndcontact >>
rect 7535 8105 7585 8155
<< ndcontact >>
rect 7685 8105 7735 8155
<< ndcontact >>
rect 7835 8105 7885 8155
<< ndcontact >>
rect 7985 8105 8035 8155
<< ndcontact >>
rect 8135 8105 8185 8155
<< ndcontact >>
rect 8285 8105 8335 8155
<< ndcontact >>
rect 8435 8105 8485 8155
<< ndcontact >>
rect 8585 8105 8635 8155
<< ndcontact >>
rect 8735 8105 8785 8155
<< ndcontact >>
rect 8885 8105 8935 8155
<< ndcontact >>
rect 9035 8105 9085 8155
<< ndcontact >>
rect 9185 8105 9235 8155
<< ndcontact >>
rect 9335 8105 9385 8155
<< ndcontact >>
rect 9485 8105 9535 8155
<< psubstratepcontact >>
rect 9995 8105 10045 8155
<< psubstratepcontact >>
rect 10145 8105 10195 8155
<< nsubstratencontact >>
rect 65 7985 115 8035
<< nsubstratencontact >>
rect 215 7985 265 8035
<< polycontact >>
rect 995 8015 1045 8065
<< polycontact >>
rect 4865 8015 4915 8065
<< polycontact >>
rect 5885 8015 5935 8065
<< polycontact >>
rect 9755 8015 9805 8065
<< psubstratepcontact >>
rect 605 7955 655 8005
<< psubstratepcontact >>
rect 755 7955 805 8005
<< ndcontact >>
rect 1265 7955 1315 8005
<< ndcontact >>
rect 1415 7955 1465 8005
<< ndcontact >>
rect 1565 7955 1615 8005
<< ndcontact >>
rect 1715 7955 1765 8005
<< ndcontact >>
rect 1865 7955 1915 8005
<< ndcontact >>
rect 2015 7955 2065 8005
<< ndcontact >>
rect 2165 7955 2215 8005
<< ndcontact >>
rect 2315 7955 2365 8005
<< ndcontact >>
rect 2465 7955 2515 8005
<< ndcontact >>
rect 2615 7955 2665 8005
<< ndcontact >>
rect 2765 7955 2815 8005
<< ndcontact >>
rect 2915 7955 2965 8005
<< ndcontact >>
rect 3065 7955 3115 8005
<< ndcontact >>
rect 3215 7955 3265 8005
<< ndcontact >>
rect 3365 7955 3415 8005
<< ndcontact >>
rect 3515 7955 3565 8005
<< ndcontact >>
rect 3665 7955 3715 8005
<< ndcontact >>
rect 3815 7955 3865 8005
<< ndcontact >>
rect 3965 7955 4015 8005
<< ndcontact >>
rect 4115 7955 4165 8005
<< ndcontact >>
rect 4265 7955 4315 8005
<< ndcontact >>
rect 4415 7955 4465 8005
<< ndcontact >>
rect 4565 7955 4615 8005
<< psubstratepcontact >>
rect 5315 7955 5365 8005
<< psubstratepcontact >>
rect 5465 7955 5515 8005
<< ndcontact >>
rect 6185 7955 6235 8005
<< ndcontact >>
rect 6335 7955 6385 8005
<< ndcontact >>
rect 6485 7955 6535 8005
<< ndcontact >>
rect 6635 7955 6685 8005
<< ndcontact >>
rect 6785 7955 6835 8005
<< ndcontact >>
rect 6935 7955 6985 8005
<< ndcontact >>
rect 7085 7955 7135 8005
<< ndcontact >>
rect 7235 7955 7285 8005
<< ndcontact >>
rect 7385 7955 7435 8005
<< ndcontact >>
rect 7535 7955 7585 8005
<< ndcontact >>
rect 7685 7955 7735 8005
<< ndcontact >>
rect 7835 7955 7885 8005
<< ndcontact >>
rect 7985 7955 8035 8005
<< ndcontact >>
rect 8135 7955 8185 8005
<< ndcontact >>
rect 8285 7955 8335 8005
<< ndcontact >>
rect 8435 7955 8485 8005
<< ndcontact >>
rect 8585 7955 8635 8005
<< ndcontact >>
rect 8735 7955 8785 8005
<< ndcontact >>
rect 8885 7955 8935 8005
<< ndcontact >>
rect 9035 7955 9085 8005
<< ndcontact >>
rect 9185 7955 9235 8005
<< ndcontact >>
rect 9335 7955 9385 8005
<< ndcontact >>
rect 9485 7955 9535 8005
<< psubstratepcontact >>
rect 9995 7955 10045 8005
<< psubstratepcontact >>
rect 10145 7955 10195 8005
<< nsubstratencontact >>
rect 10535 7985 10585 8035
<< nsubstratencontact >>
rect 10685 7985 10735 8035
<< polycontact >>
rect 995 7865 1045 7915
<< polycontact >>
rect 4865 7865 4915 7915
<< polycontact >>
rect 5885 7865 5935 7915
<< polycontact >>
rect 9755 7865 9805 7915
<< psubstratepcontact >>
rect 605 7805 655 7855
<< psubstratepcontact >>
rect 755 7805 805 7855
<< ndcontact >>
rect 1265 7805 1315 7855
<< ndcontact >>
rect 1415 7805 1465 7855
<< ndcontact >>
rect 1565 7805 1615 7855
<< ndcontact >>
rect 1715 7805 1765 7855
<< ndcontact >>
rect 1865 7805 1915 7855
<< ndcontact >>
rect 2015 7805 2065 7855
<< ndcontact >>
rect 2165 7805 2215 7855
<< ndcontact >>
rect 2315 7805 2365 7855
<< ndcontact >>
rect 2465 7805 2515 7855
<< ndcontact >>
rect 2615 7805 2665 7855
<< ndcontact >>
rect 2765 7805 2815 7855
<< ndcontact >>
rect 2915 7805 2965 7855
<< ndcontact >>
rect 3065 7805 3115 7855
<< ndcontact >>
rect 3215 7805 3265 7855
<< ndcontact >>
rect 3365 7805 3415 7855
<< ndcontact >>
rect 3515 7805 3565 7855
<< ndcontact >>
rect 3665 7805 3715 7855
<< ndcontact >>
rect 3815 7805 3865 7855
<< ndcontact >>
rect 3965 7805 4015 7855
<< ndcontact >>
rect 4115 7805 4165 7855
<< ndcontact >>
rect 4265 7805 4315 7855
<< ndcontact >>
rect 4415 7805 4465 7855
<< ndcontact >>
rect 4565 7805 4615 7855
<< psubstratepcontact >>
rect 5315 7805 5365 7855
<< psubstratepcontact >>
rect 5465 7805 5515 7855
<< ndcontact >>
rect 6185 7805 6235 7855
<< ndcontact >>
rect 6335 7805 6385 7855
<< ndcontact >>
rect 6485 7805 6535 7855
<< ndcontact >>
rect 6635 7805 6685 7855
<< ndcontact >>
rect 6785 7805 6835 7855
<< ndcontact >>
rect 6935 7805 6985 7855
<< ndcontact >>
rect 7085 7805 7135 7855
<< ndcontact >>
rect 7235 7805 7285 7855
<< ndcontact >>
rect 7385 7805 7435 7855
<< ndcontact >>
rect 7535 7805 7585 7855
<< ndcontact >>
rect 7685 7805 7735 7855
<< ndcontact >>
rect 7835 7805 7885 7855
<< ndcontact >>
rect 7985 7805 8035 7855
<< ndcontact >>
rect 8135 7805 8185 7855
<< ndcontact >>
rect 8285 7805 8335 7855
<< ndcontact >>
rect 8435 7805 8485 7855
<< ndcontact >>
rect 8585 7805 8635 7855
<< ndcontact >>
rect 8735 7805 8785 7855
<< ndcontact >>
rect 8885 7805 8935 7855
<< ndcontact >>
rect 9035 7805 9085 7855
<< ndcontact >>
rect 9185 7805 9235 7855
<< ndcontact >>
rect 9335 7805 9385 7855
<< ndcontact >>
rect 9485 7805 9535 7855
<< psubstratepcontact >>
rect 9995 7805 10045 7855
<< psubstratepcontact >>
rect 10145 7805 10195 7855
<< nsubstratencontact >>
rect 65 7745 115 7795
<< nsubstratencontact >>
rect 215 7745 265 7795
<< nsubstratencontact >>
rect 10535 7745 10585 7795
<< nsubstratencontact >>
rect 10685 7745 10735 7795
<< psubstratepcontact >>
rect 605 7655 655 7705
<< psubstratepcontact >>
rect 755 7655 805 7705
<< polycontact >>
rect 995 7685 1045 7735
<< ndcontact >>
rect 1265 7655 1315 7705
<< ndcontact >>
rect 1415 7655 1465 7705
<< ndcontact >>
rect 1565 7655 1615 7705
<< ndcontact >>
rect 1715 7655 1765 7705
<< ndcontact >>
rect 1865 7655 1915 7705
<< ndcontact >>
rect 2015 7655 2065 7705
<< ndcontact >>
rect 2165 7655 2215 7705
<< ndcontact >>
rect 2315 7655 2365 7705
<< ndcontact >>
rect 2465 7655 2515 7705
<< ndcontact >>
rect 2615 7655 2665 7705
<< ndcontact >>
rect 2765 7655 2815 7705
<< ndcontact >>
rect 2915 7655 2965 7705
<< ndcontact >>
rect 3065 7655 3115 7705
<< ndcontact >>
rect 3215 7655 3265 7705
<< ndcontact >>
rect 3365 7655 3415 7705
<< ndcontact >>
rect 3515 7655 3565 7705
<< ndcontact >>
rect 3665 7655 3715 7705
<< ndcontact >>
rect 3815 7655 3865 7705
<< ndcontact >>
rect 3965 7655 4015 7705
<< ndcontact >>
rect 4115 7655 4165 7705
<< ndcontact >>
rect 4265 7655 4315 7705
<< ndcontact >>
rect 4415 7655 4465 7705
<< ndcontact >>
rect 4565 7655 4615 7705
<< polycontact >>
rect 4865 7685 4915 7735
<< psubstratepcontact >>
rect 5315 7655 5365 7705
<< psubstratepcontact >>
rect 5465 7655 5515 7705
<< polycontact >>
rect 5885 7685 5935 7735
<< ndcontact >>
rect 6185 7655 6235 7705
<< ndcontact >>
rect 6335 7655 6385 7705
<< ndcontact >>
rect 6485 7655 6535 7705
<< ndcontact >>
rect 6635 7655 6685 7705
<< ndcontact >>
rect 6785 7655 6835 7705
<< ndcontact >>
rect 6935 7655 6985 7705
<< ndcontact >>
rect 7085 7655 7135 7705
<< ndcontact >>
rect 7235 7655 7285 7705
<< ndcontact >>
rect 7385 7655 7435 7705
<< ndcontact >>
rect 7535 7655 7585 7705
<< ndcontact >>
rect 7685 7655 7735 7705
<< ndcontact >>
rect 7835 7655 7885 7705
<< ndcontact >>
rect 7985 7655 8035 7705
<< ndcontact >>
rect 8135 7655 8185 7705
<< ndcontact >>
rect 8285 7655 8335 7705
<< ndcontact >>
rect 8435 7655 8485 7705
<< ndcontact >>
rect 8585 7655 8635 7705
<< ndcontact >>
rect 8735 7655 8785 7705
<< ndcontact >>
rect 8885 7655 8935 7705
<< ndcontact >>
rect 9035 7655 9085 7705
<< ndcontact >>
rect 9185 7655 9235 7705
<< ndcontact >>
rect 9335 7655 9385 7705
<< ndcontact >>
rect 9485 7655 9535 7705
<< polycontact >>
rect 9755 7685 9805 7735
<< psubstratepcontact >>
rect 9995 7655 10045 7705
<< psubstratepcontact >>
rect 10145 7655 10195 7705
<< nsubstratencontact >>
rect 65 7505 115 7555
<< nsubstratencontact >>
rect 215 7505 265 7555
<< psubstratepcontact >>
rect 605 7505 655 7555
<< psubstratepcontact >>
rect 755 7505 805 7555
<< polycontact >>
rect 995 7535 1045 7585
<< ndcontact >>
rect 1265 7505 1315 7555
<< ndcontact >>
rect 1415 7505 1465 7555
<< ndcontact >>
rect 1565 7505 1615 7555
<< ndcontact >>
rect 1715 7505 1765 7555
<< ndcontact >>
rect 1865 7505 1915 7555
<< ndcontact >>
rect 2015 7505 2065 7555
<< ndcontact >>
rect 2165 7505 2215 7555
<< ndcontact >>
rect 2315 7505 2365 7555
<< ndcontact >>
rect 2465 7505 2515 7555
<< ndcontact >>
rect 2615 7505 2665 7555
<< ndcontact >>
rect 2765 7505 2815 7555
<< ndcontact >>
rect 2915 7505 2965 7555
<< ndcontact >>
rect 3065 7505 3115 7555
<< ndcontact >>
rect 3215 7505 3265 7555
<< ndcontact >>
rect 3365 7505 3415 7555
<< ndcontact >>
rect 3515 7505 3565 7555
<< ndcontact >>
rect 3665 7505 3715 7555
<< ndcontact >>
rect 3815 7505 3865 7555
<< ndcontact >>
rect 3965 7505 4015 7555
<< ndcontact >>
rect 4115 7505 4165 7555
<< ndcontact >>
rect 4265 7505 4315 7555
<< ndcontact >>
rect 4415 7505 4465 7555
<< ndcontact >>
rect 4565 7505 4615 7555
<< polycontact >>
rect 4865 7535 4915 7585
<< psubstratepcontact >>
rect 5315 7505 5365 7555
<< psubstratepcontact >>
rect 5465 7505 5515 7555
<< polycontact >>
rect 5885 7535 5935 7585
<< ndcontact >>
rect 6185 7505 6235 7555
<< ndcontact >>
rect 6335 7505 6385 7555
<< ndcontact >>
rect 6485 7505 6535 7555
<< ndcontact >>
rect 6635 7505 6685 7555
<< ndcontact >>
rect 6785 7505 6835 7555
<< ndcontact >>
rect 6935 7505 6985 7555
<< ndcontact >>
rect 7085 7505 7135 7555
<< ndcontact >>
rect 7235 7505 7285 7555
<< ndcontact >>
rect 7385 7505 7435 7555
<< ndcontact >>
rect 7535 7505 7585 7555
<< ndcontact >>
rect 7685 7505 7735 7555
<< ndcontact >>
rect 7835 7505 7885 7555
<< ndcontact >>
rect 7985 7505 8035 7555
<< ndcontact >>
rect 8135 7505 8185 7555
<< ndcontact >>
rect 8285 7505 8335 7555
<< ndcontact >>
rect 8435 7505 8485 7555
<< ndcontact >>
rect 8585 7505 8635 7555
<< ndcontact >>
rect 8735 7505 8785 7555
<< ndcontact >>
rect 8885 7505 8935 7555
<< ndcontact >>
rect 9035 7505 9085 7555
<< ndcontact >>
rect 9185 7505 9235 7555
<< ndcontact >>
rect 9335 7505 9385 7555
<< ndcontact >>
rect 9485 7505 9535 7555
<< polycontact >>
rect 9755 7535 9805 7585
<< psubstratepcontact >>
rect 9995 7505 10045 7555
<< psubstratepcontact >>
rect 10145 7505 10195 7555
<< nsubstratencontact >>
rect 10535 7505 10585 7555
<< nsubstratencontact >>
rect 10685 7505 10735 7555
<< psubstratepcontact >>
rect 605 7355 655 7405
<< psubstratepcontact >>
rect 755 7355 805 7405
<< polycontact >>
rect 995 7385 1045 7435
<< ndcontact >>
rect 1265 7355 1315 7405
<< ndcontact >>
rect 1415 7355 1465 7405
<< ndcontact >>
rect 1565 7355 1615 7405
<< ndcontact >>
rect 1715 7355 1765 7405
<< ndcontact >>
rect 1865 7355 1915 7405
<< ndcontact >>
rect 2015 7355 2065 7405
<< ndcontact >>
rect 2165 7355 2215 7405
<< ndcontact >>
rect 2315 7355 2365 7405
<< ndcontact >>
rect 2465 7355 2515 7405
<< ndcontact >>
rect 2615 7355 2665 7405
<< ndcontact >>
rect 2765 7355 2815 7405
<< ndcontact >>
rect 2915 7355 2965 7405
<< ndcontact >>
rect 3065 7355 3115 7405
<< ndcontact >>
rect 3215 7355 3265 7405
<< ndcontact >>
rect 3365 7355 3415 7405
<< ndcontact >>
rect 3515 7355 3565 7405
<< ndcontact >>
rect 3665 7355 3715 7405
<< ndcontact >>
rect 3815 7355 3865 7405
<< ndcontact >>
rect 3965 7355 4015 7405
<< ndcontact >>
rect 4115 7355 4165 7405
<< ndcontact >>
rect 4265 7355 4315 7405
<< ndcontact >>
rect 4415 7355 4465 7405
<< ndcontact >>
rect 4565 7355 4615 7405
<< polycontact >>
rect 4865 7385 4915 7435
<< psubstratepcontact >>
rect 5315 7355 5365 7405
<< psubstratepcontact >>
rect 5465 7355 5515 7405
<< polycontact >>
rect 5885 7385 5935 7435
<< ndcontact >>
rect 6185 7355 6235 7405
<< ndcontact >>
rect 6335 7355 6385 7405
<< ndcontact >>
rect 6485 7355 6535 7405
<< ndcontact >>
rect 6635 7355 6685 7405
<< ndcontact >>
rect 6785 7355 6835 7405
<< ndcontact >>
rect 6935 7355 6985 7405
<< ndcontact >>
rect 7085 7355 7135 7405
<< ndcontact >>
rect 7235 7355 7285 7405
<< ndcontact >>
rect 7385 7355 7435 7405
<< ndcontact >>
rect 7535 7355 7585 7405
<< ndcontact >>
rect 7685 7355 7735 7405
<< ndcontact >>
rect 7835 7355 7885 7405
<< ndcontact >>
rect 7985 7355 8035 7405
<< ndcontact >>
rect 8135 7355 8185 7405
<< ndcontact >>
rect 8285 7355 8335 7405
<< ndcontact >>
rect 8435 7355 8485 7405
<< ndcontact >>
rect 8585 7355 8635 7405
<< ndcontact >>
rect 8735 7355 8785 7405
<< ndcontact >>
rect 8885 7355 8935 7405
<< ndcontact >>
rect 9035 7355 9085 7405
<< ndcontact >>
rect 9185 7355 9235 7405
<< ndcontact >>
rect 9335 7355 9385 7405
<< ndcontact >>
rect 9485 7355 9535 7405
<< polycontact >>
rect 9755 7385 9805 7435
<< psubstratepcontact >>
rect 9995 7355 10045 7405
<< psubstratepcontact >>
rect 10145 7355 10195 7405
<< nsubstratencontact >>
rect 65 7235 115 7285
<< nsubstratencontact >>
rect 215 7235 265 7285
<< psubstratepcontact >>
rect 605 7205 655 7255
<< psubstratepcontact >>
rect 755 7205 805 7255
<< polycontact >>
rect 995 7235 1045 7285
<< ndcontact >>
rect 1265 7205 1315 7255
<< ndcontact >>
rect 1415 7205 1465 7255
<< ndcontact >>
rect 1565 7205 1615 7255
<< ndcontact >>
rect 1715 7205 1765 7255
<< ndcontact >>
rect 1865 7205 1915 7255
<< ndcontact >>
rect 2015 7205 2065 7255
<< ndcontact >>
rect 2165 7205 2215 7255
<< ndcontact >>
rect 2315 7205 2365 7255
<< ndcontact >>
rect 2465 7205 2515 7255
<< ndcontact >>
rect 2615 7205 2665 7255
<< ndcontact >>
rect 2765 7205 2815 7255
<< ndcontact >>
rect 2915 7205 2965 7255
<< ndcontact >>
rect 3065 7205 3115 7255
<< ndcontact >>
rect 3215 7205 3265 7255
<< ndcontact >>
rect 3365 7205 3415 7255
<< ndcontact >>
rect 3515 7205 3565 7255
<< ndcontact >>
rect 3665 7205 3715 7255
<< ndcontact >>
rect 3815 7205 3865 7255
<< ndcontact >>
rect 3965 7205 4015 7255
<< ndcontact >>
rect 4115 7205 4165 7255
<< ndcontact >>
rect 4265 7205 4315 7255
<< ndcontact >>
rect 4415 7205 4465 7255
<< ndcontact >>
rect 4565 7205 4615 7255
<< polycontact >>
rect 4865 7235 4915 7285
<< psubstratepcontact >>
rect 5315 7205 5365 7255
<< psubstratepcontact >>
rect 5465 7205 5515 7255
<< polycontact >>
rect 5885 7235 5935 7285
<< ndcontact >>
rect 6185 7205 6235 7255
<< ndcontact >>
rect 6335 7205 6385 7255
<< ndcontact >>
rect 6485 7205 6535 7255
<< ndcontact >>
rect 6635 7205 6685 7255
<< ndcontact >>
rect 6785 7205 6835 7255
<< ndcontact >>
rect 6935 7205 6985 7255
<< ndcontact >>
rect 7085 7205 7135 7255
<< ndcontact >>
rect 7235 7205 7285 7255
<< ndcontact >>
rect 7385 7205 7435 7255
<< ndcontact >>
rect 7535 7205 7585 7255
<< ndcontact >>
rect 7685 7205 7735 7255
<< ndcontact >>
rect 7835 7205 7885 7255
<< ndcontact >>
rect 7985 7205 8035 7255
<< ndcontact >>
rect 8135 7205 8185 7255
<< ndcontact >>
rect 8285 7205 8335 7255
<< ndcontact >>
rect 8435 7205 8485 7255
<< ndcontact >>
rect 8585 7205 8635 7255
<< ndcontact >>
rect 8735 7205 8785 7255
<< ndcontact >>
rect 8885 7205 8935 7255
<< ndcontact >>
rect 9035 7205 9085 7255
<< ndcontact >>
rect 9185 7205 9235 7255
<< ndcontact >>
rect 9335 7205 9385 7255
<< ndcontact >>
rect 9485 7205 9535 7255
<< polycontact >>
rect 9755 7235 9805 7285
<< psubstratepcontact >>
rect 9995 7205 10045 7255
<< psubstratepcontact >>
rect 10145 7205 10195 7255
<< nsubstratencontact >>
rect 10535 7235 10585 7285
<< nsubstratencontact >>
rect 10685 7235 10735 7285
<< psubstratepcontact >>
rect 605 7055 655 7105
<< psubstratepcontact >>
rect 755 7055 805 7105
<< polycontact >>
rect 995 7085 1045 7135
<< polycontact >>
rect 4865 7085 4915 7135
<< psubstratepcontact >>
rect 5315 7055 5365 7105
<< psubstratepcontact >>
rect 5465 7055 5515 7105
<< polycontact >>
rect 5885 7085 5935 7135
<< polycontact >>
rect 9755 7085 9805 7135
<< psubstratepcontact >>
rect 9995 7055 10045 7105
<< psubstratepcontact >>
rect 10145 7055 10195 7105
<< nsubstratencontact >>
rect 65 6995 115 7045
<< nsubstratencontact >>
rect 215 6995 265 7045
<< nsubstratencontact >>
rect 10535 6995 10585 7045
<< nsubstratencontact >>
rect 10685 6995 10735 7045
<< polycontact >>
rect 995 6935 1045 6985
<< ndcontact >>
rect 1235 6905 1285 6955
<< ndcontact >>
rect 1535 6905 1585 6955
<< ndcontact >>
rect 1835 6905 1885 6955
<< ndcontact >>
rect 2135 6905 2185 6955
<< ndcontact >>
rect 2435 6905 2485 6955
<< ndcontact >>
rect 2735 6905 2785 6955
<< ndcontact >>
rect 3035 6905 3085 6955
<< ndcontact >>
rect 3335 6905 3385 6955
<< ndcontact >>
rect 4625 6905 4675 6955
<< polycontact >>
rect 4865 6935 4915 6985
<< polycontact >>
rect 5885 6935 5935 6985
<< ndcontact >>
rect 6125 6905 6175 6955
<< ndcontact >>
rect 7415 6905 7465 6955
<< ndcontact >>
rect 7715 6905 7765 6955
<< ndcontact >>
rect 8015 6905 8065 6955
<< ndcontact >>
rect 8315 6905 8365 6955
<< ndcontact >>
rect 8615 6905 8665 6955
<< ndcontact >>
rect 8915 6905 8965 6955
<< ndcontact >>
rect 9215 6905 9265 6955
<< ndcontact >>
rect 9515 6905 9565 6955
<< polycontact >>
rect 9755 6935 9805 6985
<< nsubstratencontact >>
rect 65 6755 115 6805
<< nsubstratencontact >>
rect 215 6755 265 6805
<< polycontact >>
rect 995 6785 1045 6835
<< ndcontact >>
rect 1235 6755 1285 6805
<< ndcontact >>
rect 1535 6755 1585 6805
<< ndcontact >>
rect 1835 6755 1885 6805
<< ndcontact >>
rect 2135 6755 2185 6805
<< ndcontact >>
rect 2435 6755 2485 6805
<< ndcontact >>
rect 2735 6755 2785 6805
<< ndcontact >>
rect 3035 6755 3085 6805
<< ndcontact >>
rect 3335 6755 3385 6805
<< ndcontact >>
rect 4625 6755 4675 6805
<< polycontact >>
rect 4865 6785 4915 6835
<< polycontact >>
rect 5885 6785 5935 6835
<< ndcontact >>
rect 6125 6755 6175 6805
<< ndcontact >>
rect 7415 6755 7465 6805
<< ndcontact >>
rect 7715 6755 7765 6805
<< ndcontact >>
rect 8015 6755 8065 6805
<< ndcontact >>
rect 8315 6755 8365 6805
<< ndcontact >>
rect 8615 6755 8665 6805
<< ndcontact >>
rect 8915 6755 8965 6805
<< ndcontact >>
rect 9215 6755 9265 6805
<< ndcontact >>
rect 9515 6755 9565 6805
<< polycontact >>
rect 9755 6785 9805 6835
<< nsubstratencontact >>
rect 10535 6755 10585 6805
<< nsubstratencontact >>
rect 10685 6755 10735 6805
<< polycontact >>
rect 995 6635 1045 6685
<< ndcontact >>
rect 1235 6605 1285 6655
<< ndcontact >>
rect 1535 6605 1585 6655
<< ndcontact >>
rect 1835 6605 1885 6655
<< ndcontact >>
rect 2135 6605 2185 6655
<< ndcontact >>
rect 2435 6605 2485 6655
<< ndcontact >>
rect 2735 6605 2785 6655
<< ndcontact >>
rect 3035 6605 3085 6655
<< ndcontact >>
rect 3335 6605 3385 6655
<< ndcontact >>
rect 4625 6605 4675 6655
<< polycontact >>
rect 4865 6635 4915 6685
<< polycontact >>
rect 5885 6635 5935 6685
<< ndcontact >>
rect 6125 6605 6175 6655
<< ndcontact >>
rect 7415 6605 7465 6655
<< ndcontact >>
rect 7715 6605 7765 6655
<< ndcontact >>
rect 8015 6605 8065 6655
<< ndcontact >>
rect 8315 6605 8365 6655
<< ndcontact >>
rect 8615 6605 8665 6655
<< ndcontact >>
rect 8915 6605 8965 6655
<< ndcontact >>
rect 9215 6605 9265 6655
<< ndcontact >>
rect 9515 6605 9565 6655
<< polycontact >>
rect 9755 6635 9805 6685
<< nsubstratencontact >>
rect 65 6515 115 6565
<< nsubstratencontact >>
rect 215 6515 265 6565
<< psubstratepcontact >>
rect 605 6455 655 6505
<< psubstratepcontact >>
rect 755 6455 805 6505
<< polycontact >>
rect 995 6485 1045 6535
<< polycontact >>
rect 4865 6485 4915 6535
<< psubstratepcontact >>
rect 5315 6455 5365 6505
<< psubstratepcontact >>
rect 5465 6455 5515 6505
<< polycontact >>
rect 5885 6485 5935 6535
<< polycontact >>
rect 9755 6485 9805 6535
<< nsubstratencontact >>
rect 10535 6515 10585 6565
<< nsubstratencontact >>
rect 10685 6515 10735 6565
<< psubstratepcontact >>
rect 9995 6455 10045 6505
<< psubstratepcontact >>
rect 10145 6455 10195 6505
<< nsubstratencontact >>
rect 65 6275 115 6325
<< nsubstratencontact >>
rect 215 6275 265 6325
<< psubstratepcontact >>
rect 605 6305 655 6355
<< psubstratepcontact >>
rect 755 6305 805 6355
<< polycontact >>
rect 995 6335 1045 6385
<< ndcontact >>
rect 1265 6305 1315 6355
<< ndcontact >>
rect 1415 6305 1465 6355
<< ndcontact >>
rect 1565 6305 1615 6355
<< ndcontact >>
rect 1715 6305 1765 6355
<< ndcontact >>
rect 1865 6305 1915 6355
<< ndcontact >>
rect 2015 6305 2065 6355
<< ndcontact >>
rect 2165 6305 2215 6355
<< ndcontact >>
rect 2315 6305 2365 6355
<< ndcontact >>
rect 2465 6305 2515 6355
<< ndcontact >>
rect 2615 6305 2665 6355
<< ndcontact >>
rect 2765 6305 2815 6355
<< ndcontact >>
rect 2915 6305 2965 6355
<< ndcontact >>
rect 3065 6305 3115 6355
<< ndcontact >>
rect 3215 6305 3265 6355
<< ndcontact >>
rect 3365 6305 3415 6355
<< ndcontact >>
rect 3515 6305 3565 6355
<< ndcontact >>
rect 3665 6305 3715 6355
<< ndcontact >>
rect 3815 6305 3865 6355
<< ndcontact >>
rect 3965 6305 4015 6355
<< ndcontact >>
rect 4115 6305 4165 6355
<< ndcontact >>
rect 4265 6305 4315 6355
<< ndcontact >>
rect 4415 6305 4465 6355
<< ndcontact >>
rect 4565 6305 4615 6355
<< polycontact >>
rect 4865 6335 4915 6385
<< psubstratepcontact >>
rect 5315 6305 5365 6355
<< psubstratepcontact >>
rect 5465 6305 5515 6355
<< polycontact >>
rect 5885 6335 5935 6385
<< ndcontact >>
rect 6185 6305 6235 6355
<< ndcontact >>
rect 6335 6305 6385 6355
<< ndcontact >>
rect 6485 6305 6535 6355
<< ndcontact >>
rect 6635 6305 6685 6355
<< ndcontact >>
rect 6785 6305 6835 6355
<< ndcontact >>
rect 6935 6305 6985 6355
<< ndcontact >>
rect 7085 6305 7135 6355
<< ndcontact >>
rect 7235 6305 7285 6355
<< ndcontact >>
rect 7385 6305 7435 6355
<< ndcontact >>
rect 7535 6305 7585 6355
<< ndcontact >>
rect 7685 6305 7735 6355
<< ndcontact >>
rect 7835 6305 7885 6355
<< ndcontact >>
rect 7985 6305 8035 6355
<< ndcontact >>
rect 8135 6305 8185 6355
<< ndcontact >>
rect 8285 6305 8335 6355
<< ndcontact >>
rect 8435 6305 8485 6355
<< ndcontact >>
rect 8585 6305 8635 6355
<< ndcontact >>
rect 8735 6305 8785 6355
<< ndcontact >>
rect 8885 6305 8935 6355
<< ndcontact >>
rect 9035 6305 9085 6355
<< ndcontact >>
rect 9185 6305 9235 6355
<< ndcontact >>
rect 9335 6305 9385 6355
<< ndcontact >>
rect 9485 6305 9535 6355
<< polycontact >>
rect 9755 6335 9805 6385
<< psubstratepcontact >>
rect 9995 6305 10045 6355
<< psubstratepcontact >>
rect 10145 6305 10195 6355
<< nsubstratencontact >>
rect 10535 6275 10585 6325
<< nsubstratencontact >>
rect 10685 6275 10735 6325
<< psubstratepcontact >>
rect 605 6155 655 6205
<< psubstratepcontact >>
rect 755 6155 805 6205
<< polycontact >>
rect 995 6185 1045 6235
<< ndcontact >>
rect 1265 6155 1315 6205
<< ndcontact >>
rect 1415 6155 1465 6205
<< ndcontact >>
rect 1565 6155 1615 6205
<< ndcontact >>
rect 1715 6155 1765 6205
<< ndcontact >>
rect 1865 6155 1915 6205
<< ndcontact >>
rect 2015 6155 2065 6205
<< ndcontact >>
rect 2165 6155 2215 6205
<< ndcontact >>
rect 2315 6155 2365 6205
<< ndcontact >>
rect 2465 6155 2515 6205
<< ndcontact >>
rect 2615 6155 2665 6205
<< ndcontact >>
rect 2765 6155 2815 6205
<< ndcontact >>
rect 2915 6155 2965 6205
<< ndcontact >>
rect 3065 6155 3115 6205
<< ndcontact >>
rect 3215 6155 3265 6205
<< ndcontact >>
rect 3365 6155 3415 6205
<< ndcontact >>
rect 3515 6155 3565 6205
<< ndcontact >>
rect 3665 6155 3715 6205
<< ndcontact >>
rect 3815 6155 3865 6205
<< ndcontact >>
rect 3965 6155 4015 6205
<< ndcontact >>
rect 4115 6155 4165 6205
<< ndcontact >>
rect 4265 6155 4315 6205
<< ndcontact >>
rect 4415 6155 4465 6205
<< ndcontact >>
rect 4565 6155 4615 6205
<< polycontact >>
rect 4865 6185 4915 6235
<< psubstratepcontact >>
rect 5315 6155 5365 6205
<< psubstratepcontact >>
rect 5465 6155 5515 6205
<< polycontact >>
rect 5885 6185 5935 6235
<< ndcontact >>
rect 6185 6155 6235 6205
<< ndcontact >>
rect 6335 6155 6385 6205
<< ndcontact >>
rect 6485 6155 6535 6205
<< ndcontact >>
rect 6635 6155 6685 6205
<< ndcontact >>
rect 6785 6155 6835 6205
<< ndcontact >>
rect 6935 6155 6985 6205
<< ndcontact >>
rect 7085 6155 7135 6205
<< ndcontact >>
rect 7235 6155 7285 6205
<< ndcontact >>
rect 7385 6155 7435 6205
<< ndcontact >>
rect 7535 6155 7585 6205
<< ndcontact >>
rect 7685 6155 7735 6205
<< ndcontact >>
rect 7835 6155 7885 6205
<< ndcontact >>
rect 7985 6155 8035 6205
<< ndcontact >>
rect 8135 6155 8185 6205
<< ndcontact >>
rect 8285 6155 8335 6205
<< ndcontact >>
rect 8435 6155 8485 6205
<< ndcontact >>
rect 8585 6155 8635 6205
<< ndcontact >>
rect 8735 6155 8785 6205
<< ndcontact >>
rect 8885 6155 8935 6205
<< ndcontact >>
rect 9035 6155 9085 6205
<< ndcontact >>
rect 9185 6155 9235 6205
<< ndcontact >>
rect 9335 6155 9385 6205
<< ndcontact >>
rect 9485 6155 9535 6205
<< polycontact >>
rect 9755 6185 9805 6235
<< psubstratepcontact >>
rect 9995 6155 10045 6205
<< psubstratepcontact >>
rect 10145 6155 10195 6205
<< nsubstratencontact >>
rect 65 6035 115 6085
<< nsubstratencontact >>
rect 215 6035 265 6085
<< psubstratepcontact >>
rect 605 6005 655 6055
<< psubstratepcontact >>
rect 755 6005 805 6055
<< polycontact >>
rect 995 6035 1045 6085
<< ndcontact >>
rect 1265 6005 1315 6055
<< ndcontact >>
rect 1415 6005 1465 6055
<< ndcontact >>
rect 1565 6005 1615 6055
<< ndcontact >>
rect 1715 6005 1765 6055
<< ndcontact >>
rect 1865 6005 1915 6055
<< ndcontact >>
rect 2015 6005 2065 6055
<< ndcontact >>
rect 2165 6005 2215 6055
<< ndcontact >>
rect 2315 6005 2365 6055
<< ndcontact >>
rect 2465 6005 2515 6055
<< ndcontact >>
rect 2615 6005 2665 6055
<< ndcontact >>
rect 2765 6005 2815 6055
<< ndcontact >>
rect 2915 6005 2965 6055
<< ndcontact >>
rect 3065 6005 3115 6055
<< ndcontact >>
rect 3215 6005 3265 6055
<< ndcontact >>
rect 3365 6005 3415 6055
<< ndcontact >>
rect 3515 6005 3565 6055
<< ndcontact >>
rect 3665 6005 3715 6055
<< ndcontact >>
rect 3815 6005 3865 6055
<< ndcontact >>
rect 3965 6005 4015 6055
<< ndcontact >>
rect 4115 6005 4165 6055
<< ndcontact >>
rect 4265 6005 4315 6055
<< ndcontact >>
rect 4415 6005 4465 6055
<< ndcontact >>
rect 4565 6005 4615 6055
<< polycontact >>
rect 4865 6035 4915 6085
<< psubstratepcontact >>
rect 5315 6005 5365 6055
<< psubstratepcontact >>
rect 5465 6005 5515 6055
<< polycontact >>
rect 5885 6035 5935 6085
<< ndcontact >>
rect 6185 6005 6235 6055
<< ndcontact >>
rect 6335 6005 6385 6055
<< ndcontact >>
rect 6485 6005 6535 6055
<< ndcontact >>
rect 6635 6005 6685 6055
<< ndcontact >>
rect 6785 6005 6835 6055
<< ndcontact >>
rect 6935 6005 6985 6055
<< ndcontact >>
rect 7085 6005 7135 6055
<< ndcontact >>
rect 7235 6005 7285 6055
<< ndcontact >>
rect 7385 6005 7435 6055
<< ndcontact >>
rect 7535 6005 7585 6055
<< ndcontact >>
rect 7685 6005 7735 6055
<< ndcontact >>
rect 7835 6005 7885 6055
<< ndcontact >>
rect 7985 6005 8035 6055
<< ndcontact >>
rect 8135 6005 8185 6055
<< ndcontact >>
rect 8285 6005 8335 6055
<< ndcontact >>
rect 8435 6005 8485 6055
<< ndcontact >>
rect 8585 6005 8635 6055
<< ndcontact >>
rect 8735 6005 8785 6055
<< ndcontact >>
rect 8885 6005 8935 6055
<< ndcontact >>
rect 9035 6005 9085 6055
<< ndcontact >>
rect 9185 6005 9235 6055
<< ndcontact >>
rect 9335 6005 9385 6055
<< ndcontact >>
rect 9485 6005 9535 6055
<< polycontact >>
rect 9755 6035 9805 6085
<< psubstratepcontact >>
rect 9995 6005 10045 6055
<< psubstratepcontact >>
rect 10145 6005 10195 6055
<< nsubstratencontact >>
rect 10535 6035 10585 6085
<< nsubstratencontact >>
rect 10685 6035 10735 6085
<< psubstratepcontact >>
rect 605 5855 655 5905
<< psubstratepcontact >>
rect 755 5855 805 5905
<< polycontact >>
rect 995 5885 1045 5935
<< ndcontact >>
rect 1265 5855 1315 5905
<< ndcontact >>
rect 1415 5855 1465 5905
<< ndcontact >>
rect 1565 5855 1615 5905
<< ndcontact >>
rect 1715 5855 1765 5905
<< ndcontact >>
rect 1865 5855 1915 5905
<< ndcontact >>
rect 2015 5855 2065 5905
<< ndcontact >>
rect 2165 5855 2215 5905
<< ndcontact >>
rect 2315 5855 2365 5905
<< ndcontact >>
rect 2465 5855 2515 5905
<< ndcontact >>
rect 2615 5855 2665 5905
<< ndcontact >>
rect 2765 5855 2815 5905
<< ndcontact >>
rect 2915 5855 2965 5905
<< ndcontact >>
rect 3065 5855 3115 5905
<< ndcontact >>
rect 3215 5855 3265 5905
<< ndcontact >>
rect 3365 5855 3415 5905
<< ndcontact >>
rect 3515 5855 3565 5905
<< ndcontact >>
rect 3665 5855 3715 5905
<< ndcontact >>
rect 3815 5855 3865 5905
<< ndcontact >>
rect 3965 5855 4015 5905
<< ndcontact >>
rect 4115 5855 4165 5905
<< ndcontact >>
rect 4265 5855 4315 5905
<< ndcontact >>
rect 4415 5855 4465 5905
<< ndcontact >>
rect 4565 5855 4615 5905
<< polycontact >>
rect 4865 5885 4915 5935
<< psubstratepcontact >>
rect 5315 5855 5365 5905
<< psubstratepcontact >>
rect 5465 5855 5515 5905
<< polycontact >>
rect 5885 5885 5935 5935
<< ndcontact >>
rect 6185 5855 6235 5905
<< ndcontact >>
rect 6335 5855 6385 5905
<< ndcontact >>
rect 6485 5855 6535 5905
<< ndcontact >>
rect 6635 5855 6685 5905
<< ndcontact >>
rect 6785 5855 6835 5905
<< ndcontact >>
rect 6935 5855 6985 5905
<< ndcontact >>
rect 7085 5855 7135 5905
<< ndcontact >>
rect 7235 5855 7285 5905
<< ndcontact >>
rect 7385 5855 7435 5905
<< ndcontact >>
rect 7535 5855 7585 5905
<< ndcontact >>
rect 7685 5855 7735 5905
<< ndcontact >>
rect 7835 5855 7885 5905
<< ndcontact >>
rect 7985 5855 8035 5905
<< ndcontact >>
rect 8135 5855 8185 5905
<< ndcontact >>
rect 8285 5855 8335 5905
<< ndcontact >>
rect 8435 5855 8485 5905
<< ndcontact >>
rect 8585 5855 8635 5905
<< ndcontact >>
rect 8735 5855 8785 5905
<< ndcontact >>
rect 8885 5855 8935 5905
<< ndcontact >>
rect 9035 5855 9085 5905
<< ndcontact >>
rect 9185 5855 9235 5905
<< ndcontact >>
rect 9335 5855 9385 5905
<< ndcontact >>
rect 9485 5855 9535 5905
<< polycontact >>
rect 9755 5885 9805 5935
<< psubstratepcontact >>
rect 9995 5855 10045 5905
<< psubstratepcontact >>
rect 10145 5855 10195 5905
<< nsubstratencontact >>
rect 65 5795 115 5845
<< nsubstratencontact >>
rect 215 5795 265 5845
<< nsubstratencontact >>
rect 10535 5795 10585 5845
<< nsubstratencontact >>
rect 10685 5795 10735 5845
<< psubstratepcontact >>
rect 605 5705 655 5755
<< psubstratepcontact >>
rect 755 5705 805 5755
<< polycontact >>
rect 995 5735 1045 5785
<< ndcontact >>
rect 1265 5705 1315 5755
<< ndcontact >>
rect 1415 5705 1465 5755
<< ndcontact >>
rect 1565 5705 1615 5755
<< ndcontact >>
rect 1715 5705 1765 5755
<< ndcontact >>
rect 1865 5705 1915 5755
<< ndcontact >>
rect 2015 5705 2065 5755
<< ndcontact >>
rect 2165 5705 2215 5755
<< ndcontact >>
rect 2315 5705 2365 5755
<< ndcontact >>
rect 2465 5705 2515 5755
<< ndcontact >>
rect 2615 5705 2665 5755
<< ndcontact >>
rect 2765 5705 2815 5755
<< ndcontact >>
rect 2915 5705 2965 5755
<< ndcontact >>
rect 3065 5705 3115 5755
<< ndcontact >>
rect 3215 5705 3265 5755
<< ndcontact >>
rect 3365 5705 3415 5755
<< ndcontact >>
rect 3515 5705 3565 5755
<< ndcontact >>
rect 3665 5705 3715 5755
<< ndcontact >>
rect 3815 5705 3865 5755
<< ndcontact >>
rect 3965 5705 4015 5755
<< ndcontact >>
rect 4115 5705 4165 5755
<< ndcontact >>
rect 4265 5705 4315 5755
<< ndcontact >>
rect 4415 5705 4465 5755
<< ndcontact >>
rect 4565 5705 4615 5755
<< polycontact >>
rect 4865 5735 4915 5785
<< psubstratepcontact >>
rect 5315 5705 5365 5755
<< psubstratepcontact >>
rect 5465 5705 5515 5755
<< polycontact >>
rect 5885 5735 5935 5785
<< ndcontact >>
rect 6185 5705 6235 5755
<< ndcontact >>
rect 6335 5705 6385 5755
<< ndcontact >>
rect 6485 5705 6535 5755
<< ndcontact >>
rect 6635 5705 6685 5755
<< ndcontact >>
rect 6785 5705 6835 5755
<< ndcontact >>
rect 6935 5705 6985 5755
<< ndcontact >>
rect 7085 5705 7135 5755
<< ndcontact >>
rect 7235 5705 7285 5755
<< ndcontact >>
rect 7385 5705 7435 5755
<< ndcontact >>
rect 7535 5705 7585 5755
<< ndcontact >>
rect 7685 5705 7735 5755
<< ndcontact >>
rect 7835 5705 7885 5755
<< ndcontact >>
rect 7985 5705 8035 5755
<< ndcontact >>
rect 8135 5705 8185 5755
<< ndcontact >>
rect 8285 5705 8335 5755
<< ndcontact >>
rect 8435 5705 8485 5755
<< ndcontact >>
rect 8585 5705 8635 5755
<< ndcontact >>
rect 8735 5705 8785 5755
<< ndcontact >>
rect 8885 5705 8935 5755
<< ndcontact >>
rect 9035 5705 9085 5755
<< ndcontact >>
rect 9185 5705 9235 5755
<< ndcontact >>
rect 9335 5705 9385 5755
<< ndcontact >>
rect 9485 5705 9535 5755
<< polycontact >>
rect 9755 5735 9805 5785
<< psubstratepcontact >>
rect 9995 5705 10045 5755
<< psubstratepcontact >>
rect 10145 5705 10195 5755
<< nsubstratencontact >>
rect 65 5555 115 5605
<< nsubstratencontact >>
rect 215 5555 265 5605
<< psubstratepcontact >>
rect 605 5555 655 5605
<< psubstratepcontact >>
rect 755 5555 805 5605
<< polycontact >>
rect 995 5585 1045 5635
<< ndcontact >>
rect 1265 5555 1315 5605
<< ndcontact >>
rect 1415 5555 1465 5605
<< ndcontact >>
rect 1565 5555 1615 5605
<< ndcontact >>
rect 1715 5555 1765 5605
<< ndcontact >>
rect 1865 5555 1915 5605
<< ndcontact >>
rect 2015 5555 2065 5605
<< ndcontact >>
rect 2165 5555 2215 5605
<< ndcontact >>
rect 2315 5555 2365 5605
<< ndcontact >>
rect 2465 5555 2515 5605
<< ndcontact >>
rect 2615 5555 2665 5605
<< ndcontact >>
rect 2765 5555 2815 5605
<< ndcontact >>
rect 2915 5555 2965 5605
<< ndcontact >>
rect 3065 5555 3115 5605
<< ndcontact >>
rect 3215 5555 3265 5605
<< ndcontact >>
rect 3365 5555 3415 5605
<< ndcontact >>
rect 3515 5555 3565 5605
<< ndcontact >>
rect 3665 5555 3715 5605
<< ndcontact >>
rect 3815 5555 3865 5605
<< ndcontact >>
rect 3965 5555 4015 5605
<< ndcontact >>
rect 4115 5555 4165 5605
<< ndcontact >>
rect 4265 5555 4315 5605
<< ndcontact >>
rect 4415 5555 4465 5605
<< ndcontact >>
rect 4565 5555 4615 5605
<< polycontact >>
rect 4865 5585 4915 5635
<< psubstratepcontact >>
rect 5315 5555 5365 5605
<< psubstratepcontact >>
rect 5465 5555 5515 5605
<< polycontact >>
rect 5885 5585 5935 5635
<< ndcontact >>
rect 6185 5555 6235 5605
<< ndcontact >>
rect 6335 5555 6385 5605
<< ndcontact >>
rect 6485 5555 6535 5605
<< ndcontact >>
rect 6635 5555 6685 5605
<< ndcontact >>
rect 6785 5555 6835 5605
<< ndcontact >>
rect 6935 5555 6985 5605
<< ndcontact >>
rect 7085 5555 7135 5605
<< ndcontact >>
rect 7235 5555 7285 5605
<< ndcontact >>
rect 7385 5555 7435 5605
<< ndcontact >>
rect 7535 5555 7585 5605
<< ndcontact >>
rect 7685 5555 7735 5605
<< ndcontact >>
rect 7835 5555 7885 5605
<< ndcontact >>
rect 7985 5555 8035 5605
<< ndcontact >>
rect 8135 5555 8185 5605
<< ndcontact >>
rect 8285 5555 8335 5605
<< ndcontact >>
rect 8435 5555 8485 5605
<< ndcontact >>
rect 8585 5555 8635 5605
<< ndcontact >>
rect 8735 5555 8785 5605
<< ndcontact >>
rect 8885 5555 8935 5605
<< ndcontact >>
rect 9035 5555 9085 5605
<< ndcontact >>
rect 9185 5555 9235 5605
<< ndcontact >>
rect 9335 5555 9385 5605
<< ndcontact >>
rect 9485 5555 9535 5605
<< polycontact >>
rect 9755 5585 9805 5635
<< psubstratepcontact >>
rect 9995 5555 10045 5605
<< psubstratepcontact >>
rect 10145 5555 10195 5605
<< nsubstratencontact >>
rect 10535 5555 10585 5605
<< nsubstratencontact >>
rect 10685 5555 10735 5605
<< psubstratepcontact >>
rect 605 5405 655 5455
<< psubstratepcontact >>
rect 755 5405 805 5455
<< polycontact >>
rect 995 5435 1045 5485
<< ndcontact >>
rect 1265 5405 1315 5455
<< ndcontact >>
rect 1415 5405 1465 5455
<< ndcontact >>
rect 1565 5405 1615 5455
<< ndcontact >>
rect 1715 5405 1765 5455
<< ndcontact >>
rect 1865 5405 1915 5455
<< ndcontact >>
rect 2015 5405 2065 5455
<< ndcontact >>
rect 2165 5405 2215 5455
<< ndcontact >>
rect 2315 5405 2365 5455
<< ndcontact >>
rect 2465 5405 2515 5455
<< ndcontact >>
rect 2615 5405 2665 5455
<< ndcontact >>
rect 2765 5405 2815 5455
<< ndcontact >>
rect 2915 5405 2965 5455
<< ndcontact >>
rect 3065 5405 3115 5455
<< ndcontact >>
rect 3215 5405 3265 5455
<< ndcontact >>
rect 3365 5405 3415 5455
<< ndcontact >>
rect 3515 5405 3565 5455
<< ndcontact >>
rect 3665 5405 3715 5455
<< ndcontact >>
rect 3815 5405 3865 5455
<< ndcontact >>
rect 3965 5405 4015 5455
<< ndcontact >>
rect 4115 5405 4165 5455
<< ndcontact >>
rect 4265 5405 4315 5455
<< ndcontact >>
rect 4415 5405 4465 5455
<< ndcontact >>
rect 4565 5405 4615 5455
<< polycontact >>
rect 4865 5435 4915 5485
<< psubstratepcontact >>
rect 5315 5405 5365 5455
<< psubstratepcontact >>
rect 5465 5405 5515 5455
<< polycontact >>
rect 5885 5435 5935 5485
<< ndcontact >>
rect 6185 5405 6235 5455
<< ndcontact >>
rect 6335 5405 6385 5455
<< ndcontact >>
rect 6485 5405 6535 5455
<< ndcontact >>
rect 6635 5405 6685 5455
<< ndcontact >>
rect 6785 5405 6835 5455
<< ndcontact >>
rect 6935 5405 6985 5455
<< ndcontact >>
rect 7085 5405 7135 5455
<< ndcontact >>
rect 7235 5405 7285 5455
<< ndcontact >>
rect 7385 5405 7435 5455
<< ndcontact >>
rect 7535 5405 7585 5455
<< ndcontact >>
rect 7685 5405 7735 5455
<< ndcontact >>
rect 7835 5405 7885 5455
<< ndcontact >>
rect 7985 5405 8035 5455
<< ndcontact >>
rect 8135 5405 8185 5455
<< ndcontact >>
rect 8285 5405 8335 5455
<< ndcontact >>
rect 8435 5405 8485 5455
<< ndcontact >>
rect 8585 5405 8635 5455
<< ndcontact >>
rect 8735 5405 8785 5455
<< ndcontact >>
rect 8885 5405 8935 5455
<< ndcontact >>
rect 9035 5405 9085 5455
<< ndcontact >>
rect 9185 5405 9235 5455
<< ndcontact >>
rect 9335 5405 9385 5455
<< ndcontact >>
rect 9485 5405 9535 5455
<< polycontact >>
rect 9755 5435 9805 5485
<< psubstratepcontact >>
rect 9995 5405 10045 5455
<< psubstratepcontact >>
rect 10145 5405 10195 5455
<< nsubstratencontact >>
rect 65 5315 115 5365
<< nsubstratencontact >>
rect 215 5315 265 5365
<< psubstratepcontact >>
rect 605 5255 655 5305
<< psubstratepcontact >>
rect 755 5255 805 5305
<< polycontact >>
rect 995 5285 1045 5335
<< ndcontact >>
rect 1265 5255 1315 5305
<< ndcontact >>
rect 1415 5255 1465 5305
<< ndcontact >>
rect 1565 5255 1615 5305
<< ndcontact >>
rect 1715 5255 1765 5305
<< ndcontact >>
rect 1865 5255 1915 5305
<< ndcontact >>
rect 2015 5255 2065 5305
<< ndcontact >>
rect 2165 5255 2215 5305
<< ndcontact >>
rect 2315 5255 2365 5305
<< ndcontact >>
rect 2465 5255 2515 5305
<< ndcontact >>
rect 2615 5255 2665 5305
<< ndcontact >>
rect 2765 5255 2815 5305
<< ndcontact >>
rect 2915 5255 2965 5305
<< ndcontact >>
rect 3065 5255 3115 5305
<< ndcontact >>
rect 3215 5255 3265 5305
<< ndcontact >>
rect 3365 5255 3415 5305
<< ndcontact >>
rect 3515 5255 3565 5305
<< ndcontact >>
rect 3665 5255 3715 5305
<< ndcontact >>
rect 3815 5255 3865 5305
<< ndcontact >>
rect 3965 5255 4015 5305
<< ndcontact >>
rect 4115 5255 4165 5305
<< ndcontact >>
rect 4265 5255 4315 5305
<< ndcontact >>
rect 4415 5255 4465 5305
<< ndcontact >>
rect 4565 5255 4615 5305
<< polycontact >>
rect 4865 5285 4915 5335
<< psubstratepcontact >>
rect 5315 5255 5365 5305
<< psubstratepcontact >>
rect 5465 5255 5515 5305
<< polycontact >>
rect 5885 5285 5935 5335
<< ndcontact >>
rect 6185 5255 6235 5305
<< ndcontact >>
rect 6335 5255 6385 5305
<< ndcontact >>
rect 6485 5255 6535 5305
<< ndcontact >>
rect 6635 5255 6685 5305
<< ndcontact >>
rect 6785 5255 6835 5305
<< ndcontact >>
rect 6935 5255 6985 5305
<< ndcontact >>
rect 7085 5255 7135 5305
<< ndcontact >>
rect 7235 5255 7285 5305
<< ndcontact >>
rect 7385 5255 7435 5305
<< ndcontact >>
rect 7535 5255 7585 5305
<< ndcontact >>
rect 7685 5255 7735 5305
<< ndcontact >>
rect 7835 5255 7885 5305
<< ndcontact >>
rect 7985 5255 8035 5305
<< ndcontact >>
rect 8135 5255 8185 5305
<< ndcontact >>
rect 8285 5255 8335 5305
<< ndcontact >>
rect 8435 5255 8485 5305
<< ndcontact >>
rect 8585 5255 8635 5305
<< ndcontact >>
rect 8735 5255 8785 5305
<< ndcontact >>
rect 8885 5255 8935 5305
<< ndcontact >>
rect 9035 5255 9085 5305
<< ndcontact >>
rect 9185 5255 9235 5305
<< ndcontact >>
rect 9335 5255 9385 5305
<< ndcontact >>
rect 9485 5255 9535 5305
<< polycontact >>
rect 9755 5285 9805 5335
<< nsubstratencontact >>
rect 10535 5315 10585 5365
<< nsubstratencontact >>
rect 10685 5315 10735 5365
<< psubstratepcontact >>
rect 9995 5255 10045 5305
<< psubstratepcontact >>
rect 10145 5255 10195 5305
<< nsubstratencontact >>
rect 65 5075 115 5125
<< nsubstratencontact >>
rect 215 5075 265 5125
<< psubstratepcontact >>
rect 605 5105 655 5155
<< psubstratepcontact >>
rect 755 5105 805 5155
<< polycontact >>
rect 995 5135 1045 5185
<< polycontact >>
rect 4865 5135 4915 5185
<< psubstratepcontact >>
rect 5315 5105 5365 5155
<< psubstratepcontact >>
rect 5465 5105 5515 5155
<< polycontact >>
rect 5885 5135 5935 5185
<< polycontact >>
rect 9755 5135 9805 5185
<< psubstratepcontact >>
rect 9995 5105 10045 5155
<< psubstratepcontact >>
rect 10145 5105 10195 5155
<< nsubstratencontact >>
rect 10535 5075 10585 5125
<< nsubstratencontact >>
rect 10685 5075 10735 5125
<< ndcontact >>
rect 1235 4955 1285 5005
<< ndcontact >>
rect 1535 4955 1585 5005
<< ndcontact >>
rect 1835 4955 1885 5005
<< ndcontact >>
rect 2135 4955 2185 5005
<< ndcontact >>
rect 2435 4955 2485 5005
<< ndcontact >>
rect 2735 4955 2785 5005
<< ndcontact >>
rect 3035 4955 3085 5005
<< ndcontact >>
rect 3335 4955 3385 5005
<< ndcontact >>
rect 4625 4955 4675 5005
<< ndcontact >>
rect 6125 4955 6175 5005
<< ndcontact >>
rect 7415 4955 7465 5005
<< ndcontact >>
rect 7715 4955 7765 5005
<< ndcontact >>
rect 8015 4955 8065 5005
<< ndcontact >>
rect 8315 4955 8365 5005
<< ndcontact >>
rect 8615 4955 8665 5005
<< ndcontact >>
rect 8915 4955 8965 5005
<< ndcontact >>
rect 9215 4955 9265 5005
<< ndcontact >>
rect 9515 4955 9565 5005
<< nsubstratencontact >>
rect 65 4835 115 4885
<< nsubstratencontact >>
rect 215 4835 265 4885
<< ndcontact >>
rect 1235 4805 1285 4855
<< ndcontact >>
rect 1535 4805 1585 4855
<< ndcontact >>
rect 1835 4805 1885 4855
<< ndcontact >>
rect 2135 4805 2185 4855
<< ndcontact >>
rect 2435 4805 2485 4855
<< ndcontact >>
rect 2735 4805 2785 4855
<< ndcontact >>
rect 3035 4805 3085 4855
<< ndcontact >>
rect 3335 4805 3385 4855
<< ndcontact >>
rect 4625 4805 4675 4855
<< ndcontact >>
rect 6125 4805 6175 4855
<< ndcontact >>
rect 7415 4805 7465 4855
<< ndcontact >>
rect 7715 4805 7765 4855
<< ndcontact >>
rect 8015 4805 8065 4855
<< ndcontact >>
rect 8315 4805 8365 4855
<< ndcontact >>
rect 8615 4805 8665 4855
<< ndcontact >>
rect 8915 4805 8965 4855
<< ndcontact >>
rect 9215 4805 9265 4855
<< ndcontact >>
rect 9515 4805 9565 4855
<< nsubstratencontact >>
rect 10535 4835 10585 4885
<< nsubstratencontact >>
rect 10685 4835 10735 4885
<< psubstratepcontact >>
rect 1235 4655 1285 4705
<< psubstratepcontact >>
rect 1535 4655 1585 4705
<< psubstratepcontact >>
rect 1835 4655 1885 4705
<< psubstratepcontact >>
rect 2135 4655 2185 4705
<< psubstratepcontact >>
rect 2435 4655 2485 4705
<< psubstratepcontact >>
rect 2735 4655 2785 4705
<< psubstratepcontact >>
rect 3035 4655 3085 4705
<< psubstratepcontact >>
rect 3335 4655 3385 4705
<< psubstratepcontact >>
rect 4625 4655 4675 4705
<< psubstratepcontact >>
rect 6125 4655 6175 4705
<< psubstratepcontact >>
rect 7415 4655 7465 4705
<< psubstratepcontact >>
rect 7715 4655 7765 4705
<< psubstratepcontact >>
rect 8015 4655 8065 4705
<< psubstratepcontact >>
rect 8315 4655 8365 4705
<< psubstratepcontact >>
rect 8615 4655 8665 4705
<< psubstratepcontact >>
rect 8915 4655 8965 4705
<< psubstratepcontact >>
rect 9215 4655 9265 4705
<< psubstratepcontact >>
rect 9515 4655 9565 4705
<< nsubstratencontact >>
rect 65 4595 115 4645
<< nsubstratencontact >>
rect 215 4595 265 4645
<< nsubstratencontact >>
rect 10535 4595 10585 4645
<< nsubstratencontact >>
rect 10685 4595 10735 4645
<< nsubstratencontact >>
rect 65 4355 115 4405
<< nsubstratencontact >>
rect 215 4355 265 4405
<< nsubstratencontact >>
rect 10535 4355 10585 4405
<< nsubstratencontact >>
rect 10685 4355 10735 4405
<< nsubstratencontact >>
rect 275 4115 325 4165
<< nsubstratencontact >>
rect 515 4115 565 4165
<< nsubstratencontact >>
rect 755 4115 805 4165
<< nsubstratencontact >>
rect 995 4115 1045 4165
<< nsubstratencontact >>
rect 1235 4115 1285 4165
<< nsubstratencontact >>
rect 1475 4115 1525 4165
<< nsubstratencontact >>
rect 1715 4115 1765 4165
<< nsubstratencontact >>
rect 1955 4115 2005 4165
<< nsubstratencontact >>
rect 2195 4115 2245 4165
<< nsubstratencontact >>
rect 2435 4115 2485 4165
<< nsubstratencontact >>
rect 2675 4115 2725 4165
<< nsubstratencontact >>
rect 2915 4115 2965 4165
<< nsubstratencontact >>
rect 3155 4115 3205 4165
<< nsubstratencontact >>
rect 3395 4115 3445 4165
<< nsubstratencontact >>
rect 4595 4115 4645 4165
<< nsubstratencontact >>
rect 4835 4115 4885 4165
<< nsubstratencontact >>
rect 5075 4115 5125 4165
<< nsubstratencontact >>
rect 5315 4115 5365 4165
<< nsubstratencontact >>
rect 5555 4115 5605 4165
<< nsubstratencontact >>
rect 5795 4115 5845 4165
<< nsubstratencontact >>
rect 6155 4115 6205 4165
<< nsubstratencontact >>
rect 7355 4115 7405 4165
<< nsubstratencontact >>
rect 7595 4115 7645 4165
<< nsubstratencontact >>
rect 7835 4115 7885 4165
<< nsubstratencontact >>
rect 8075 4115 8125 4165
<< nsubstratencontact >>
rect 8315 4115 8365 4165
<< nsubstratencontact >>
rect 8555 4115 8605 4165
<< nsubstratencontact >>
rect 8795 4115 8845 4165
<< nsubstratencontact >>
rect 9035 4115 9085 4165
<< nsubstratencontact >>
rect 9275 4115 9325 4165
<< nsubstratencontact >>
rect 9515 4115 9565 4165
<< nsubstratencontact >>
rect 9755 4115 9805 4165
<< nsubstratencontact >>
rect 9995 4115 10045 4165
<< nsubstratencontact >>
rect 10235 4115 10285 4165
<< nsubstratencontact >>
rect 10475 4115 10525 4165
<< nsubstratencontact >>
rect 275 3965 325 4015
<< nsubstratencontact >>
rect 515 3965 565 4015
<< nsubstratencontact >>
rect 755 3965 805 4015
<< nsubstratencontact >>
rect 995 3965 1045 4015
<< nsubstratencontact >>
rect 1235 3965 1285 4015
<< nsubstratencontact >>
rect 1475 3965 1525 4015
<< nsubstratencontact >>
rect 1715 3965 1765 4015
<< nsubstratencontact >>
rect 1955 3965 2005 4015
<< nsubstratencontact >>
rect 2195 3965 2245 4015
<< nsubstratencontact >>
rect 2435 3965 2485 4015
<< nsubstratencontact >>
rect 2675 3965 2725 4015
<< nsubstratencontact >>
rect 2915 3965 2965 4015
<< nsubstratencontact >>
rect 3155 3965 3205 4015
<< nsubstratencontact >>
rect 3395 3965 3445 4015
<< nsubstratencontact >>
rect 4595 3965 4645 4015
<< nsubstratencontact >>
rect 4835 3965 4885 4015
<< nsubstratencontact >>
rect 5075 3965 5125 4015
<< nsubstratencontact >>
rect 5315 3965 5365 4015
<< nsubstratencontact >>
rect 5555 3965 5605 4015
<< nsubstratencontact >>
rect 5795 3965 5845 4015
<< nsubstratencontact >>
rect 6155 3965 6205 4015
<< nsubstratencontact >>
rect 7355 3965 7405 4015
<< nsubstratencontact >>
rect 7595 3965 7645 4015
<< nsubstratencontact >>
rect 7835 3965 7885 4015
<< nsubstratencontact >>
rect 8075 3965 8125 4015
<< nsubstratencontact >>
rect 8315 3965 8365 4015
<< nsubstratencontact >>
rect 8555 3965 8605 4015
<< nsubstratencontact >>
rect 8795 3965 8845 4015
<< nsubstratencontact >>
rect 9035 3965 9085 4015
<< nsubstratencontact >>
rect 9275 3965 9325 4015
<< nsubstratencontact >>
rect 9515 3965 9565 4015
<< nsubstratencontact >>
rect 9755 3965 9805 4015
<< nsubstratencontact >>
rect 9995 3965 10045 4015
<< nsubstratencontact >>
rect 10235 3965 10285 4015
<< nsubstratencontact >>
rect 10475 3965 10525 4015
<< psubstratepcontact >>
rect 275 3605 325 3655
<< psubstratepcontact >>
rect 515 3605 565 3655
<< psubstratepcontact >>
rect 755 3605 805 3655
<< psubstratepcontact >>
rect 995 3605 1045 3655
<< psubstratepcontact >>
rect 1235 3605 1285 3655
<< psubstratepcontact >>
rect 1475 3605 1525 3655
<< psubstratepcontact >>
rect 1715 3605 1765 3655
<< psubstratepcontact >>
rect 1955 3605 2005 3655
<< psubstratepcontact >>
rect 2195 3605 2245 3655
<< psubstratepcontact >>
rect 2435 3605 2485 3655
<< psubstratepcontact >>
rect 2675 3605 2725 3655
<< psubstratepcontact >>
rect 2915 3605 2965 3655
<< psubstratepcontact >>
rect 3155 3605 3205 3655
<< psubstratepcontact >>
rect 3395 3605 3445 3655
<< psubstratepcontact >>
rect 4595 3605 4645 3655
<< psubstratepcontact >>
rect 4835 3605 4885 3655
<< psubstratepcontact >>
rect 5075 3605 5125 3655
<< psubstratepcontact >>
rect 5315 3605 5365 3655
<< psubstratepcontact >>
rect 5555 3605 5605 3655
<< psubstratepcontact >>
rect 5795 3605 5845 3655
<< psubstratepcontact >>
rect 6155 3605 6205 3655
<< psubstratepcontact >>
rect 7355 3605 7405 3655
<< psubstratepcontact >>
rect 7595 3605 7645 3655
<< psubstratepcontact >>
rect 7835 3605 7885 3655
<< psubstratepcontact >>
rect 8075 3605 8125 3655
<< psubstratepcontact >>
rect 8315 3605 8365 3655
<< psubstratepcontact >>
rect 8555 3605 8605 3655
<< psubstratepcontact >>
rect 8795 3605 8845 3655
<< psubstratepcontact >>
rect 9035 3605 9085 3655
<< psubstratepcontact >>
rect 9275 3605 9325 3655
<< psubstratepcontact >>
rect 9515 3605 9565 3655
<< psubstratepcontact >>
rect 9755 3605 9805 3655
<< psubstratepcontact >>
rect 9995 3605 10045 3655
<< psubstratepcontact >>
rect 10235 3605 10285 3655
<< psubstratepcontact >>
rect 10475 3605 10525 3655
<< psubstratepcontact >>
rect 65 3515 115 3565
<< psubstratepcontact >>
rect 10685 3515 10735 3565
<< psubstratepcontact >>
rect 275 3455 325 3505
<< psubstratepcontact >>
rect 515 3455 565 3505
<< psubstratepcontact >>
rect 755 3455 805 3505
<< psubstratepcontact >>
rect 995 3455 1045 3505
<< psubstratepcontact >>
rect 1235 3455 1285 3505
<< psubstratepcontact >>
rect 1475 3455 1525 3505
<< psubstratepcontact >>
rect 1715 3455 1765 3505
<< psubstratepcontact >>
rect 1955 3455 2005 3505
<< psubstratepcontact >>
rect 2195 3455 2245 3505
<< psubstratepcontact >>
rect 2435 3455 2485 3505
<< psubstratepcontact >>
rect 2675 3455 2725 3505
<< psubstratepcontact >>
rect 2915 3455 2965 3505
<< psubstratepcontact >>
rect 3155 3455 3205 3505
<< psubstratepcontact >>
rect 3395 3455 3445 3505
<< psubstratepcontact >>
rect 4595 3455 4645 3505
<< psubstratepcontact >>
rect 4835 3455 4885 3505
<< psubstratepcontact >>
rect 5075 3455 5125 3505
<< psubstratepcontact >>
rect 5315 3455 5365 3505
<< psubstratepcontact >>
rect 5555 3455 5605 3505
<< psubstratepcontact >>
rect 5795 3455 5845 3505
<< psubstratepcontact >>
rect 6155 3455 6205 3505
<< psubstratepcontact >>
rect 7355 3455 7405 3505
<< psubstratepcontact >>
rect 7595 3455 7645 3505
<< psubstratepcontact >>
rect 7835 3455 7885 3505
<< psubstratepcontact >>
rect 8075 3455 8125 3505
<< psubstratepcontact >>
rect 8315 3455 8365 3505
<< psubstratepcontact >>
rect 8555 3455 8605 3505
<< psubstratepcontact >>
rect 8795 3455 8845 3505
<< psubstratepcontact >>
rect 9035 3455 9085 3505
<< psubstratepcontact >>
rect 9275 3455 9325 3505
<< psubstratepcontact >>
rect 9515 3455 9565 3505
<< psubstratepcontact >>
rect 9755 3455 9805 3505
<< psubstratepcontact >>
rect 9995 3455 10045 3505
<< psubstratepcontact >>
rect 10235 3455 10285 3505
<< psubstratepcontact >>
rect 10475 3455 10525 3505
<< psubstratepcontact >>
rect 65 3365 115 3415
<< psubstratepcontact >>
rect 10685 3365 10735 3415
<< psubstratepcontact >>
rect 65 3215 115 3265
<< psubstratepcontact >>
rect 215 3215 265 3265
<< psubstratepcontact >>
rect 10535 3215 10585 3265
<< psubstratepcontact >>
rect 10685 3215 10735 3265
<< psubstratepcontact >>
rect 65 3065 115 3115
<< psubstratepcontact >>
rect 215 3065 265 3115
<< psubstratepcontact >>
rect 10535 3065 10585 3115
<< psubstratepcontact >>
rect 10685 3065 10735 3115
<< psubstratepcontact >>
rect 65 2915 115 2965
<< psubstratepcontact >>
rect 215 2915 265 2965
<< psubstratepcontact >>
rect 10535 2915 10585 2965
<< psubstratepcontact >>
rect 10685 2915 10735 2965
<< psubstratepcontact >>
rect 65 2765 115 2815
<< psubstratepcontact >>
rect 215 2765 265 2815
<< psubstratepcontact >>
rect 10535 2765 10585 2815
<< psubstratepcontact >>
rect 10685 2765 10735 2815
<< psubstratepcontact >>
rect 65 2615 115 2665
<< psubstratepcontact >>
rect 215 2615 265 2665
<< ndcontact >>
rect 1025 2645 1075 2695
<< ndcontact >>
rect 1175 2645 1225 2695
<< ndcontact >>
rect 1325 2645 1375 2695
<< ndcontact >>
rect 1475 2645 1525 2695
<< ndcontact >>
rect 1625 2645 1675 2695
<< ndcontact >>
rect 1775 2645 1825 2695
<< ndcontact >>
rect 1925 2645 1975 2695
<< ndcontact >>
rect 2075 2645 2125 2695
<< ndcontact >>
rect 8675 2645 8725 2695
<< ndcontact >>
rect 8825 2645 8875 2695
<< ndcontact >>
rect 8975 2645 9025 2695
<< ndcontact >>
rect 9125 2645 9175 2695
<< ndcontact >>
rect 9275 2645 9325 2695
<< ndcontact >>
rect 9425 2645 9475 2695
<< ndcontact >>
rect 9575 2645 9625 2695
<< ndcontact >>
rect 9725 2645 9775 2695
<< psubstratepcontact >>
rect 10535 2615 10585 2665
<< psubstratepcontact >>
rect 10685 2615 10735 2665
<< psubstratepcontact >>
rect 65 2465 115 2515
<< psubstratepcontact >>
rect 215 2465 265 2515
<< psubstratepcontact >>
rect 10535 2465 10585 2515
<< psubstratepcontact >>
rect 10685 2465 10735 2515
<< ndcontact >>
rect 905 2405 955 2455
<< ndcontact >>
rect 1055 2405 1105 2455
<< ndcontact >>
rect 1205 2405 1255 2455
<< ndcontact >>
rect 1355 2405 1405 2455
<< ndcontact >>
rect 1505 2405 1555 2455
<< ndcontact >>
rect 1655 2405 1705 2455
<< ndcontact >>
rect 9095 2405 9145 2455
<< ndcontact >>
rect 9245 2405 9295 2455
<< ndcontact >>
rect 9395 2405 9445 2455
<< ndcontact >>
rect 9545 2405 9595 2455
<< ndcontact >>
rect 9695 2405 9745 2455
<< ndcontact >>
rect 9845 2405 9895 2455
<< psubstratepcontact >>
rect 65 2315 115 2365
<< psubstratepcontact >>
rect 215 2315 265 2365
<< polycontact >>
rect 725 2315 775 2365
<< nsubstratencontact >>
rect 2585 2345 2635 2395
<< nsubstratencontact >>
rect 2735 2345 2785 2395
<< nsubstratencontact >>
rect 2885 2345 2935 2395
<< nsubstratencontact >>
rect 3035 2345 3085 2395
<< nsubstratencontact >>
rect 3185 2345 3235 2395
<< nsubstratencontact >>
rect 3335 2345 3385 2395
<< nsubstratencontact >>
rect 3485 2345 3535 2395
<< nsubstratencontact >>
rect 3635 2345 3685 2395
<< nsubstratencontact >>
rect 3785 2345 3835 2395
<< nsubstratencontact >>
rect 3935 2345 3985 2395
<< nsubstratencontact >>
rect 4085 2345 4135 2395
<< nsubstratencontact >>
rect 4235 2345 4285 2395
<< nsubstratencontact >>
rect 4385 2345 4435 2395
<< nsubstratencontact >>
rect 4535 2345 4585 2395
<< nsubstratencontact >>
rect 4685 2345 4735 2395
<< nsubstratencontact >>
rect 4835 2345 4885 2395
<< nsubstratencontact >>
rect 4985 2345 5035 2395
<< nsubstratencontact >>
rect 5135 2345 5185 2395
<< nsubstratencontact >>
rect 5285 2345 5335 2395
<< nsubstratencontact >>
rect 5435 2345 5485 2395
<< nsubstratencontact >>
rect 5585 2345 5635 2395
<< nsubstratencontact >>
rect 5735 2345 5785 2395
<< nsubstratencontact >>
rect 5885 2345 5935 2395
<< nsubstratencontact >>
rect 6035 2345 6085 2395
<< nsubstratencontact >>
rect 6185 2345 6235 2395
<< nsubstratencontact >>
rect 6335 2345 6385 2395
<< nsubstratencontact >>
rect 6485 2345 6535 2395
<< nsubstratencontact >>
rect 6635 2345 6685 2395
<< nsubstratencontact >>
rect 6785 2345 6835 2395
<< nsubstratencontact >>
rect 6935 2345 6985 2395
<< nsubstratencontact >>
rect 7085 2345 7135 2395
<< nsubstratencontact >>
rect 7235 2345 7285 2395
<< nsubstratencontact >>
rect 7385 2345 7435 2395
<< nsubstratencontact >>
rect 7535 2345 7585 2395
<< nsubstratencontact >>
rect 7685 2345 7735 2395
<< nsubstratencontact >>
rect 7835 2345 7885 2395
<< nsubstratencontact >>
rect 7985 2345 8035 2395
<< nsubstratencontact >>
rect 8135 2345 8185 2395
<< polycontact >>
rect 10025 2315 10075 2365
<< psubstratepcontact >>
rect 10535 2315 10585 2365
<< psubstratepcontact >>
rect 10685 2315 10735 2365
<< psubstratepcontact >>
rect 65 2165 115 2215
<< psubstratepcontact >>
rect 215 2165 265 2215
<< polycontact >>
rect 725 2165 775 2215
<< ndcontact >>
rect 1475 2165 1525 2215
<< ndcontact >>
rect 1625 2165 1675 2215
<< ndcontact >>
rect 1775 2165 1825 2215
<< ndcontact >>
rect 1925 2165 1975 2215
<< ndcontact >>
rect 2075 2165 2125 2215
<< nsubstratencontact >>
rect 2585 2195 2635 2245
<< nsubstratencontact >>
rect 2735 2195 2785 2245
<< nsubstratencontact >>
rect 2885 2195 2935 2245
<< nsubstratencontact >>
rect 3035 2195 3085 2245
<< nsubstratencontact >>
rect 3185 2195 3235 2245
<< nsubstratencontact >>
rect 3335 2195 3385 2245
<< nsubstratencontact >>
rect 3485 2195 3535 2245
<< nsubstratencontact >>
rect 3635 2195 3685 2245
<< nsubstratencontact >>
rect 3785 2195 3835 2245
<< nsubstratencontact >>
rect 3935 2195 3985 2245
<< nsubstratencontact >>
rect 4085 2195 4135 2245
<< nsubstratencontact >>
rect 4235 2195 4285 2245
<< nsubstratencontact >>
rect 4385 2195 4435 2245
<< nsubstratencontact >>
rect 4535 2195 4585 2245
<< nsubstratencontact >>
rect 4685 2195 4735 2245
<< nsubstratencontact >>
rect 4835 2195 4885 2245
<< nsubstratencontact >>
rect 4985 2195 5035 2245
<< nsubstratencontact >>
rect 5135 2195 5185 2245
<< nsubstratencontact >>
rect 5285 2195 5335 2245
<< nsubstratencontact >>
rect 5435 2195 5485 2245
<< nsubstratencontact >>
rect 5585 2195 5635 2245
<< nsubstratencontact >>
rect 5735 2195 5785 2245
<< nsubstratencontact >>
rect 5885 2195 5935 2245
<< nsubstratencontact >>
rect 6035 2195 6085 2245
<< nsubstratencontact >>
rect 6185 2195 6235 2245
<< nsubstratencontact >>
rect 6335 2195 6385 2245
<< nsubstratencontact >>
rect 6485 2195 6535 2245
<< nsubstratencontact >>
rect 6635 2195 6685 2245
<< nsubstratencontact >>
rect 6785 2195 6835 2245
<< nsubstratencontact >>
rect 6935 2195 6985 2245
<< nsubstratencontact >>
rect 7085 2195 7135 2245
<< nsubstratencontact >>
rect 7235 2195 7285 2245
<< nsubstratencontact >>
rect 7385 2195 7435 2245
<< nsubstratencontact >>
rect 7535 2195 7585 2245
<< nsubstratencontact >>
rect 7685 2195 7735 2245
<< nsubstratencontact >>
rect 7835 2195 7885 2245
<< nsubstratencontact >>
rect 7985 2195 8035 2245
<< nsubstratencontact >>
rect 8135 2195 8185 2245
<< ndcontact >>
rect 8675 2165 8725 2215
<< ndcontact >>
rect 8825 2165 8875 2215
<< ndcontact >>
rect 8975 2165 9025 2215
<< ndcontact >>
rect 9125 2165 9175 2215
<< ndcontact >>
rect 9275 2165 9325 2215
<< polycontact >>
rect 10025 2165 10075 2215
<< psubstratepcontact >>
rect 10535 2165 10585 2215
<< psubstratepcontact >>
rect 10685 2165 10735 2215
<< psubstratepcontact >>
rect 65 2015 115 2065
<< psubstratepcontact >>
rect 215 2015 265 2065
<< polycontact >>
rect 725 2015 775 2065
<< polycontact >>
rect 10025 2015 10075 2065
<< psubstratepcontact >>
rect 10535 2015 10585 2065
<< psubstratepcontact >>
rect 10685 2015 10735 2065
<< ndcontact >>
rect 905 1925 955 1975
<< ndcontact >>
rect 1055 1925 1105 1975
<< ndcontact >>
rect 1205 1925 1255 1975
<< ndcontact >>
rect 1355 1925 1405 1975
<< ndcontact >>
rect 1505 1925 1555 1975
<< ndcontact >>
rect 1655 1925 1705 1975
<< ndcontact >>
rect 9095 1925 9145 1975
<< ndcontact >>
rect 9245 1925 9295 1975
<< ndcontact >>
rect 9395 1925 9445 1975
<< ndcontact >>
rect 9545 1925 9595 1975
<< ndcontact >>
rect 9695 1925 9745 1975
<< ndcontact >>
rect 9845 1925 9895 1975
<< psubstratepcontact >>
rect 65 1865 115 1915
<< psubstratepcontact >>
rect 215 1865 265 1915
<< polycontact >>
rect 725 1865 775 1915
<< polycontact >>
rect 10025 1865 10075 1915
<< psubstratepcontact >>
rect 10535 1865 10585 1915
<< psubstratepcontact >>
rect 10685 1865 10735 1915
<< psubstratepcontact >>
rect 65 1715 115 1765
<< psubstratepcontact >>
rect 215 1715 265 1765
<< polycontact >>
rect 725 1715 775 1765
<< ndcontact >>
rect 1475 1685 1525 1735
<< ndcontact >>
rect 1625 1685 1675 1735
<< ndcontact >>
rect 1775 1685 1825 1735
<< ndcontact >>
rect 1925 1685 1975 1735
<< ndcontact >>
rect 2075 1685 2125 1735
<< ndcontact >>
rect 8675 1685 8725 1735
<< ndcontact >>
rect 8825 1685 8875 1735
<< ndcontact >>
rect 8975 1685 9025 1735
<< ndcontact >>
rect 9125 1685 9175 1735
<< ndcontact >>
rect 9275 1685 9325 1735
<< polycontact >>
rect 10025 1715 10075 1765
<< psubstratepcontact >>
rect 10535 1715 10585 1765
<< psubstratepcontact >>
rect 10685 1715 10735 1765
<< psubstratepcontact >>
rect 65 1565 115 1615
<< psubstratepcontact >>
rect 215 1565 265 1615
<< polycontact >>
rect 725 1565 775 1615
<< polycontact >>
rect 10025 1565 10075 1615
<< psubstratepcontact >>
rect 10535 1565 10585 1615
<< psubstratepcontact >>
rect 10685 1565 10735 1615
<< psubstratepcontact >>
rect 65 1415 115 1465
<< psubstratepcontact >>
rect 215 1415 265 1465
<< polycontact >>
rect 725 1415 775 1465
<< ndcontact >>
rect 905 1445 955 1495
<< ndcontact >>
rect 1055 1445 1105 1495
<< ndcontact >>
rect 1205 1445 1255 1495
<< ndcontact >>
rect 1355 1445 1405 1495
<< ndcontact >>
rect 1505 1445 1555 1495
<< ndcontact >>
rect 1655 1445 1705 1495
<< ndcontact >>
rect 9095 1445 9145 1495
<< ndcontact >>
rect 9245 1445 9295 1495
<< ndcontact >>
rect 9395 1445 9445 1495
<< ndcontact >>
rect 9545 1445 9595 1495
<< ndcontact >>
rect 9695 1445 9745 1495
<< ndcontact >>
rect 9845 1445 9895 1495
<< polycontact >>
rect 10025 1415 10075 1465
<< psubstratepcontact >>
rect 10535 1415 10585 1465
<< psubstratepcontact >>
rect 10685 1415 10735 1465
<< psubstratepcontact >>
rect 65 1265 115 1315
<< psubstratepcontact >>
rect 215 1265 265 1315
<< polycontact >>
rect 725 1265 775 1315
<< nsubstratencontact >>
rect 2585 1295 2635 1345
<< nsubstratencontact >>
rect 2735 1295 2785 1345
<< nsubstratencontact >>
rect 2885 1295 2935 1345
<< nsubstratencontact >>
rect 3035 1295 3085 1345
<< nsubstratencontact >>
rect 3185 1295 3235 1345
<< nsubstratencontact >>
rect 3335 1295 3385 1345
<< nsubstratencontact >>
rect 3485 1295 3535 1345
<< nsubstratencontact >>
rect 3635 1295 3685 1345
<< nsubstratencontact >>
rect 3785 1295 3835 1345
<< nsubstratencontact >>
rect 3935 1295 3985 1345
<< nsubstratencontact >>
rect 4085 1295 4135 1345
<< nsubstratencontact >>
rect 4235 1295 4285 1345
<< nsubstratencontact >>
rect 4385 1295 4435 1345
<< nsubstratencontact >>
rect 4535 1295 4585 1345
<< nsubstratencontact >>
rect 4685 1295 4735 1345
<< nsubstratencontact >>
rect 4835 1295 4885 1345
<< nsubstratencontact >>
rect 4985 1295 5035 1345
<< nsubstratencontact >>
rect 5135 1295 5185 1345
<< nsubstratencontact >>
rect 5285 1295 5335 1345
<< nsubstratencontact >>
rect 5435 1295 5485 1345
<< nsubstratencontact >>
rect 5585 1295 5635 1345
<< nsubstratencontact >>
rect 5735 1295 5785 1345
<< nsubstratencontact >>
rect 5885 1295 5935 1345
<< nsubstratencontact >>
rect 6035 1295 6085 1345
<< nsubstratencontact >>
rect 6185 1295 6235 1345
<< nsubstratencontact >>
rect 6335 1295 6385 1345
<< nsubstratencontact >>
rect 6485 1295 6535 1345
<< nsubstratencontact >>
rect 6635 1295 6685 1345
<< nsubstratencontact >>
rect 6785 1295 6835 1345
<< nsubstratencontact >>
rect 6935 1295 6985 1345
<< nsubstratencontact >>
rect 7085 1295 7135 1345
<< nsubstratencontact >>
rect 7235 1295 7285 1345
<< nsubstratencontact >>
rect 7385 1295 7435 1345
<< nsubstratencontact >>
rect 7535 1295 7585 1345
<< nsubstratencontact >>
rect 7685 1295 7735 1345
<< nsubstratencontact >>
rect 7835 1295 7885 1345
<< nsubstratencontact >>
rect 7985 1295 8035 1345
<< nsubstratencontact >>
rect 8135 1295 8185 1345
<< nsubstratencontact >>
rect 8285 1295 8335 1345
<< polycontact >>
rect 10025 1265 10075 1315
<< psubstratepcontact >>
rect 10535 1265 10585 1315
<< psubstratepcontact >>
rect 10685 1265 10735 1315
<< ndcontact >>
rect 1475 1205 1525 1255
<< ndcontact >>
rect 1625 1205 1675 1255
<< ndcontact >>
rect 1775 1205 1825 1255
<< ndcontact >>
rect 1925 1205 1975 1255
<< ndcontact >>
rect 2075 1205 2125 1255
<< ndcontact >>
rect 8675 1205 8725 1255
<< ndcontact >>
rect 8825 1205 8875 1255
<< ndcontact >>
rect 8975 1205 9025 1255
<< ndcontact >>
rect 9125 1205 9175 1255
<< ndcontact >>
rect 9275 1205 9325 1255
<< psubstratepcontact >>
rect 65 1115 115 1165
<< psubstratepcontact >>
rect 215 1115 265 1165
<< polycontact >>
rect 725 1115 775 1165
<< nsubstratencontact >>
rect 2585 1145 2635 1195
<< nsubstratencontact >>
rect 2735 1145 2785 1195
<< nsubstratencontact >>
rect 2885 1145 2935 1195
<< nsubstratencontact >>
rect 3035 1145 3085 1195
<< nsubstratencontact >>
rect 3185 1145 3235 1195
<< nsubstratencontact >>
rect 3335 1145 3385 1195
<< nsubstratencontact >>
rect 3485 1145 3535 1195
<< nsubstratencontact >>
rect 3635 1145 3685 1195
<< nsubstratencontact >>
rect 3785 1145 3835 1195
<< nsubstratencontact >>
rect 3935 1145 3985 1195
<< nsubstratencontact >>
rect 4085 1145 4135 1195
<< nsubstratencontact >>
rect 4235 1145 4285 1195
<< nsubstratencontact >>
rect 4385 1145 4435 1195
<< nsubstratencontact >>
rect 4535 1145 4585 1195
<< nsubstratencontact >>
rect 4685 1145 4735 1195
<< nsubstratencontact >>
rect 4835 1145 4885 1195
<< nsubstratencontact >>
rect 4985 1145 5035 1195
<< nsubstratencontact >>
rect 5135 1145 5185 1195
<< nsubstratencontact >>
rect 5285 1145 5335 1195
<< nsubstratencontact >>
rect 5435 1145 5485 1195
<< nsubstratencontact >>
rect 5585 1145 5635 1195
<< nsubstratencontact >>
rect 5735 1145 5785 1195
<< nsubstratencontact >>
rect 5885 1145 5935 1195
<< nsubstratencontact >>
rect 6035 1145 6085 1195
<< nsubstratencontact >>
rect 6185 1145 6235 1195
<< nsubstratencontact >>
rect 6335 1145 6385 1195
<< nsubstratencontact >>
rect 6485 1145 6535 1195
<< nsubstratencontact >>
rect 6635 1145 6685 1195
<< nsubstratencontact >>
rect 6785 1145 6835 1195
<< nsubstratencontact >>
rect 6935 1145 6985 1195
<< nsubstratencontact >>
rect 7085 1145 7135 1195
<< nsubstratencontact >>
rect 7235 1145 7285 1195
<< nsubstratencontact >>
rect 7385 1145 7435 1195
<< nsubstratencontact >>
rect 7535 1145 7585 1195
<< nsubstratencontact >>
rect 7685 1145 7735 1195
<< nsubstratencontact >>
rect 7835 1145 7885 1195
<< nsubstratencontact >>
rect 7985 1145 8035 1195
<< nsubstratencontact >>
rect 8135 1145 8185 1195
<< nsubstratencontact >>
rect 8285 1145 8335 1195
<< polycontact >>
rect 10025 1115 10075 1165
<< psubstratepcontact >>
rect 10535 1115 10585 1165
<< psubstratepcontact >>
rect 10685 1115 10735 1165
<< psubstratepcontact >>
rect 65 965 115 1015
<< psubstratepcontact >>
rect 215 965 265 1015
<< polycontact >>
rect 725 965 775 1015
<< ndcontact >>
rect 905 965 955 1015
<< ndcontact >>
rect 1055 965 1105 1015
<< ndcontact >>
rect 1205 965 1255 1015
<< ndcontact >>
rect 1355 965 1405 1015
<< ndcontact >>
rect 1505 965 1555 1015
<< ndcontact >>
rect 1655 965 1705 1015
<< ndcontact >>
rect 9095 965 9145 1015
<< ndcontact >>
rect 9245 965 9295 1015
<< ndcontact >>
rect 9395 965 9445 1015
<< ndcontact >>
rect 9545 965 9595 1015
<< ndcontact >>
rect 9695 965 9745 1015
<< ndcontact >>
rect 9845 965 9895 1015
<< polycontact >>
rect 10025 965 10075 1015
<< psubstratepcontact >>
rect 10535 965 10585 1015
<< psubstratepcontact >>
rect 10685 965 10735 1015
<< psubstratepcontact >>
rect 65 815 115 865
<< psubstratepcontact >>
rect 215 815 265 865
<< polycontact >>
rect 725 815 775 865
<< polycontact >>
rect 10025 815 10075 865
<< psubstratepcontact >>
rect 10535 815 10585 865
<< psubstratepcontact >>
rect 10685 815 10735 865
<< ndcontact >>
rect 1475 725 1525 775
<< ndcontact >>
rect 1625 725 1675 775
<< ndcontact >>
rect 1775 725 1825 775
<< ndcontact >>
rect 1925 725 1975 775
<< ndcontact >>
rect 2075 725 2125 775
<< ndcontact >>
rect 8675 725 8725 775
<< ndcontact >>
rect 8825 725 8875 775
<< ndcontact >>
rect 8975 725 9025 775
<< ndcontact >>
rect 9125 725 9175 775
<< ndcontact >>
rect 9275 725 9325 775
<< psubstratepcontact >>
rect 65 665 115 715
<< psubstratepcontact >>
rect 215 665 265 715
<< polycontact >>
rect 725 665 775 715
<< polycontact >>
rect 10025 665 10075 715
<< psubstratepcontact >>
rect 10535 665 10585 715
<< psubstratepcontact >>
rect 10685 665 10735 715
<< psubstratepcontact >>
rect 65 515 115 565
<< psubstratepcontact >>
rect 215 515 265 565
<< polycontact >>
rect 725 515 775 565
<< ndcontact >>
rect 905 485 955 535
<< ndcontact >>
rect 1055 485 1105 535
<< ndcontact >>
rect 1205 485 1255 535
<< ndcontact >>
rect 1355 485 1405 535
<< ndcontact >>
rect 1505 485 1555 535
<< ndcontact >>
rect 1655 485 1705 535
<< ndcontact >>
rect 1805 485 1855 535
<< ndcontact >>
rect 1955 485 2005 535
<< ndcontact >>
rect 8795 485 8845 535
<< ndcontact >>
rect 8945 485 8995 535
<< ndcontact >>
rect 9095 485 9145 535
<< ndcontact >>
rect 9245 485 9295 535
<< ndcontact >>
rect 9395 485 9445 535
<< ndcontact >>
rect 9545 485 9595 535
<< ndcontact >>
rect 9695 485 9745 535
<< ndcontact >>
rect 9845 485 9895 535
<< polycontact >>
rect 10025 515 10075 565
<< psubstratepcontact >>
rect 10535 515 10585 565
<< psubstratepcontact >>
rect 10685 515 10735 565
<< psubstratepcontact >>
rect 65 365 115 415
<< psubstratepcontact >>
rect 215 365 265 415
<< psubstratepcontact >>
rect 10535 365 10585 415
<< psubstratepcontact >>
rect 10685 365 10735 415
<< psubstratepcontact >>
rect 65 215 115 265
<< psubstratepcontact >>
rect 215 215 265 265
<< psubstratepcontact >>
rect 755 215 805 265
<< psubstratepcontact >>
rect 995 215 1045 265
<< psubstratepcontact >>
rect 1235 215 1285 265
<< psubstratepcontact >>
rect 1475 215 1525 265
<< psubstratepcontact >>
rect 1715 215 1765 265
<< psubstratepcontact >>
rect 1955 215 2005 265
<< psubstratepcontact >>
rect 2195 215 2245 265
<< psubstratepcontact >>
rect 2435 215 2485 265
<< psubstratepcontact >>
rect 2675 215 2725 265
<< psubstratepcontact >>
rect 2915 215 2965 265
<< psubstratepcontact >>
rect 3155 215 3205 265
<< psubstratepcontact >>
rect 3395 215 3445 265
<< psubstratepcontact >>
rect 3635 215 3685 265
<< psubstratepcontact >>
rect 3875 215 3925 265
<< psubstratepcontact >>
rect 4115 215 4165 265
<< psubstratepcontact >>
rect 4355 215 4405 265
<< psubstratepcontact >>
rect 4595 215 4645 265
<< psubstratepcontact >>
rect 4835 215 4885 265
<< psubstratepcontact >>
rect 5915 215 5965 265
<< psubstratepcontact >>
rect 6155 215 6205 265
<< psubstratepcontact >>
rect 6395 215 6445 265
<< psubstratepcontact >>
rect 6635 215 6685 265
<< psubstratepcontact >>
rect 6875 215 6925 265
<< psubstratepcontact >>
rect 7115 215 7165 265
<< psubstratepcontact >>
rect 7355 215 7405 265
<< psubstratepcontact >>
rect 7595 215 7645 265
<< psubstratepcontact >>
rect 7835 215 7885 265
<< psubstratepcontact >>
rect 8075 215 8125 265
<< psubstratepcontact >>
rect 8315 215 8365 265
<< psubstratepcontact >>
rect 8555 215 8605 265
<< psubstratepcontact >>
rect 8795 215 8845 265
<< psubstratepcontact >>
rect 9035 215 9085 265
<< psubstratepcontact >>
rect 9275 215 9325 265
<< psubstratepcontact >>
rect 9515 215 9565 265
<< psubstratepcontact >>
rect 9755 215 9805 265
<< psubstratepcontact >>
rect 9995 215 10045 265
<< psubstratepcontact >>
rect 10535 215 10585 265
<< psubstratepcontact >>
rect 10685 215 10735 265
<< psubstratepcontact >>
rect 65 65 115 115
<< psubstratepcontact >>
rect 215 65 265 115
<< psubstratepcontact >>
rect 755 65 805 115
<< psubstratepcontact >>
rect 995 65 1045 115
<< psubstratepcontact >>
rect 1235 65 1285 115
<< psubstratepcontact >>
rect 1475 65 1525 115
<< psubstratepcontact >>
rect 1715 65 1765 115
<< psubstratepcontact >>
rect 1955 65 2005 115
<< psubstratepcontact >>
rect 2195 65 2245 115
<< psubstratepcontact >>
rect 2435 65 2485 115
<< psubstratepcontact >>
rect 2675 65 2725 115
<< psubstratepcontact >>
rect 2915 65 2965 115
<< psubstratepcontact >>
rect 3155 65 3205 115
<< psubstratepcontact >>
rect 3395 65 3445 115
<< psubstratepcontact >>
rect 3635 65 3685 115
<< psubstratepcontact >>
rect 3875 65 3925 115
<< psubstratepcontact >>
rect 4115 65 4165 115
<< psubstratepcontact >>
rect 4355 65 4405 115
<< psubstratepcontact >>
rect 4595 65 4645 115
<< psubstratepcontact >>
rect 4835 65 4885 115
<< psubstratepcontact >>
rect 5915 65 5965 115
<< psubstratepcontact >>
rect 6155 65 6205 115
<< psubstratepcontact >>
rect 6395 65 6445 115
<< psubstratepcontact >>
rect 6635 65 6685 115
<< psubstratepcontact >>
rect 6875 65 6925 115
<< psubstratepcontact >>
rect 7115 65 7165 115
<< psubstratepcontact >>
rect 7355 65 7405 115
<< psubstratepcontact >>
rect 7595 65 7645 115
<< psubstratepcontact >>
rect 7835 65 7885 115
<< psubstratepcontact >>
rect 8075 65 8125 115
<< psubstratepcontact >>
rect 8315 65 8365 115
<< psubstratepcontact >>
rect 8555 65 8605 115
<< psubstratepcontact >>
rect 8795 65 8845 115
<< psubstratepcontact >>
rect 9035 65 9085 115
<< psubstratepcontact >>
rect 9275 65 9325 115
<< psubstratepcontact >>
rect 9515 65 9565 115
<< psubstratepcontact >>
rect 9755 65 9805 115
<< psubstratepcontact >>
rect 9995 65 10045 115
<< psubstratepcontact >>
rect 10535 65 10585 115
<< psubstratepcontact >>
rect 10685 65 10735 115
<< metal1 >>
rect 1350 23010 9450 31110
rect 1860 22710 8940 23010
rect 2160 22410 8640 22710
rect 2460 22110 8340 22410
rect 2760 21810 8040 22110
rect 3060 21510 7740 21810
rect 3360 21210 7440 21510
rect 3600 21120 7200 21210
rect 0 20520 3510 20850
rect 0 13470 330 20520
rect 540 19680 3450 20160
rect 540 14310 1080 19680
rect 3600 19530 4290 21120
rect 4470 20520 6330 20850
rect 4440 19680 6360 20160
rect 1230 18360 4950 19530
rect 1170 17730 3450 18210
rect 3600 17580 4290 18360
rect 4440 17730 4920 18210
rect 1230 16410 4950 17580
rect 1170 15780 3450 16260
rect 3600 15630 4290 16410
rect 4440 15780 4920 16260
rect 1230 14460 4950 15630
rect 540 13830 3450 14310
rect 0 13140 3510 13470
rect 0 12630 3510 12960
rect 0 11790 3510 12120
rect 0 11280 3510 11610
rect 0 4230 330 11280
rect 540 10440 3450 10920
rect 540 5070 1080 10440
rect 3600 10290 4290 14460
rect 5040 14310 5760 19680
rect 6510 19530 7200 21120
rect 7290 20520 10800 20850
rect 7350 19680 10260 20160
rect 5850 18360 9570 19530
rect 5880 17730 6360 18210
rect 6510 17580 7200 18360
rect 7350 17730 9630 18210
rect 5850 16410 9570 17580
rect 5880 15780 6360 16260
rect 6510 15630 7200 16410
rect 7350 15780 9630 16260
rect 5850 14460 9570 15630
rect 4440 13830 6360 14310
rect 4440 13140 6300 13470
rect 4440 12630 6300 12960
rect 4440 11790 4860 12120
rect 5250 11790 5550 12120
rect 5880 11790 6300 12120
rect 4440 11280 6300 11610
rect 4440 10440 6360 10920
rect 1230 9120 4650 10290
rect 1170 8490 3450 8970
rect 3600 8340 4290 9120
rect 4440 8490 4710 8970
rect 1230 7170 4650 8340
rect 1170 6540 3450 7020
rect 3600 6390 4290 7170
rect 4440 6540 4710 7020
rect 1230 5220 4650 6390
rect 540 4590 3450 5070
rect 0 3900 3480 4230
rect 0 3390 3510 3720
rect 0 330 330 3390
rect 3600 3000 4290 5220
rect 4830 5070 5970 10440
rect 6510 10290 7200 14460
rect 9720 14310 10260 19680
rect 7350 13830 10260 14310
rect 10470 13470 10800 20520
rect 7290 13140 10800 13470
rect 7290 12630 10800 12960
rect 7290 11790 10800 12120
rect 7290 11280 10800 11610
rect 7350 10440 10260 10920
rect 6150 9120 9570 10290
rect 6090 8490 6360 8970
rect 6510 8340 7200 9120
rect 7350 8490 9630 8970
rect 6150 7170 9570 8340
rect 6090 6540 6360 7020
rect 6510 6390 7200 7170
rect 7350 6540 9630 7020
rect 6150 5220 9570 6390
rect 4440 4590 6360 5070
rect 4440 3900 6360 4230
rect 4440 3390 6360 3720
rect 3510 2910 4290 3000
rect 3330 2820 4290 2910
rect 6510 3000 7200 5220
rect 9720 5070 10260 10440
rect 7350 4590 10260 5070
rect 10470 4230 10800 11280
rect 7320 3900 10800 4230
rect 7290 3390 10800 3720
rect 6510 2910 7290 3000
rect 6510 2820 7470 2910
rect 3150 2730 4380 2820
rect 6420 2730 7650 2820
rect 900 2610 2430 2730
rect 2970 2640 4560 2730
rect 6240 2640 7830 2730
rect 690 2370 1770 2490
rect 690 2010 1350 2370
rect 1890 2250 2430 2610
rect 2790 2550 4740 2640
rect 6060 2550 8010 2640
rect 8370 2610 9900 2730
rect 2610 2460 4890 2550
rect 5910 2460 8190 2550
rect 1440 2130 2430 2250
rect 2550 2130 8220 2460
rect 8370 2250 8910 2610
rect 9030 2370 10110 2490
rect 8370 2130 9360 2250
rect 690 1890 1770 2010
rect 690 1530 1350 1890
rect 1890 1770 2430 2130
rect 1440 1650 2430 1770
rect 690 1410 1770 1530
rect 1890 1410 2430 1650
rect 8370 1770 8910 2130
rect 9450 2010 10110 2370
rect 9030 1890 10110 2010
rect 8370 1650 9360 1770
rect 8370 1410 8910 1650
rect 9450 1530 10110 1890
rect 9030 1410 10110 1530
rect 690 1050 1350 1410
rect 1890 1290 8910 1410
rect 1440 1170 9360 1290
rect 690 930 1770 1050
rect 690 570 1350 930
rect 1890 810 8910 1170
rect 9450 1050 10110 1410
rect 9030 930 10110 1050
rect 1440 690 9360 810
rect 4050 630 6750 690
rect 690 330 2160 570
rect 4410 540 6390 630
rect 9450 570 10110 930
rect 4770 450 6030 540
rect 0 0 5100 330
rect 5250 0 5610 450
rect 8640 330 10110 570
rect 10470 330 10800 3390
rect 5760 0 10800 330
<< metal2 >>
rect 1410 23070 9390 31050
rect 0 20520 10800 20850
rect 0 19680 10800 20160
rect 0 18540 10800 19350
rect 0 17730 10800 18210
rect 0 16740 10800 17550
rect 0 15780 10800 16260
rect 5790 15750 6270 15780
rect 0 14790 10800 15600
rect 0 13830 10800 14310
rect 5790 13800 6270 13830
rect 0 13140 10800 13470
rect 0 12630 10800 12960
rect 0 11790 10800 12120
rect 0 11280 10800 11610
rect 0 10440 10800 10920
rect 0 9300 10800 10110
rect 0 8490 10800 8970
rect 0 7500 10800 8310
rect 0 6540 10800 7020
rect 0 5550 10800 6360
rect 0 4590 10800 5070
rect 0 3900 10800 4230
rect 0 3390 10800 3720
rect 0 1560 1350 2340
rect 8670 1560 10800 2340
rect 0 0 10800 330
<< via1 >>
rect 1775 30635 1825 30685
rect 2075 30635 2125 30685
rect 2375 30635 2425 30685
rect 2675 30635 2725 30685
rect 2975 30635 3025 30685
rect 3275 30635 3325 30685
rect 3575 30635 3625 30685
rect 3875 30635 3925 30685
rect 4175 30635 4225 30685
rect 4475 30635 4525 30685
rect 4775 30635 4825 30685
rect 5075 30635 5125 30685
rect 5375 30635 5425 30685
rect 5675 30635 5725 30685
rect 5975 30635 6025 30685
rect 6275 30635 6325 30685
rect 6575 30635 6625 30685
rect 6875 30635 6925 30685
rect 7175 30635 7225 30685
rect 7475 30635 7525 30685
rect 7775 30635 7825 30685
rect 8075 30635 8125 30685
rect 8375 30635 8425 30685
rect 8675 30635 8725 30685
rect 8975 30635 9025 30685
rect 1775 30335 1825 30385
rect 2075 30335 2125 30385
rect 2375 30335 2425 30385
rect 2675 30335 2725 30385
rect 2975 30335 3025 30385
rect 3275 30335 3325 30385
rect 3575 30335 3625 30385
rect 3875 30335 3925 30385
rect 4175 30335 4225 30385
rect 4475 30335 4525 30385
rect 4775 30335 4825 30385
rect 5075 30335 5125 30385
rect 5375 30335 5425 30385
rect 5675 30335 5725 30385
rect 5975 30335 6025 30385
rect 6275 30335 6325 30385
rect 6575 30335 6625 30385
rect 6875 30335 6925 30385
rect 7175 30335 7225 30385
rect 7475 30335 7525 30385
rect 7775 30335 7825 30385
rect 8075 30335 8125 30385
rect 8375 30335 8425 30385
rect 8675 30335 8725 30385
rect 8975 30335 9025 30385
rect 1775 30035 1825 30085
rect 2075 30035 2125 30085
rect 2375 30035 2425 30085
rect 2675 30035 2725 30085
rect 2975 30035 3025 30085
rect 3275 30035 3325 30085
rect 3575 30035 3625 30085
rect 3875 30035 3925 30085
rect 4175 30035 4225 30085
rect 4475 30035 4525 30085
rect 4775 30035 4825 30085
rect 5075 30035 5125 30085
rect 5375 30035 5425 30085
rect 5675 30035 5725 30085
rect 5975 30035 6025 30085
rect 6275 30035 6325 30085
rect 6575 30035 6625 30085
rect 6875 30035 6925 30085
rect 7175 30035 7225 30085
rect 7475 30035 7525 30085
rect 7775 30035 7825 30085
rect 8075 30035 8125 30085
rect 8375 30035 8425 30085
rect 8675 30035 8725 30085
rect 8975 30035 9025 30085
rect 1775 29735 1825 29785
rect 2075 29735 2125 29785
rect 2375 29735 2425 29785
rect 2675 29735 2725 29785
rect 2975 29735 3025 29785
rect 3275 29735 3325 29785
rect 3575 29735 3625 29785
rect 3875 29735 3925 29785
rect 4175 29735 4225 29785
rect 4475 29735 4525 29785
rect 4775 29735 4825 29785
rect 5075 29735 5125 29785
rect 5375 29735 5425 29785
rect 5675 29735 5725 29785
rect 5975 29735 6025 29785
rect 6275 29735 6325 29785
rect 6575 29735 6625 29785
rect 6875 29735 6925 29785
rect 7175 29735 7225 29785
rect 7475 29735 7525 29785
rect 7775 29735 7825 29785
rect 8075 29735 8125 29785
rect 8375 29735 8425 29785
rect 8675 29735 8725 29785
rect 8975 29735 9025 29785
rect 1775 29435 1825 29485
rect 2075 29435 2125 29485
rect 2375 29435 2425 29485
rect 2675 29435 2725 29485
rect 2975 29435 3025 29485
rect 3275 29435 3325 29485
rect 3575 29435 3625 29485
rect 3875 29435 3925 29485
rect 4175 29435 4225 29485
rect 4475 29435 4525 29485
rect 4775 29435 4825 29485
rect 5075 29435 5125 29485
rect 5375 29435 5425 29485
rect 5675 29435 5725 29485
rect 5975 29435 6025 29485
rect 6275 29435 6325 29485
rect 6575 29435 6625 29485
rect 6875 29435 6925 29485
rect 7175 29435 7225 29485
rect 7475 29435 7525 29485
rect 7775 29435 7825 29485
rect 8075 29435 8125 29485
rect 8375 29435 8425 29485
rect 8675 29435 8725 29485
rect 8975 29435 9025 29485
rect 1775 29135 1825 29185
rect 2075 29135 2125 29185
rect 2375 29135 2425 29185
rect 2675 29135 2725 29185
rect 2975 29135 3025 29185
rect 3275 29135 3325 29185
rect 3575 29135 3625 29185
rect 3875 29135 3925 29185
rect 4175 29135 4225 29185
rect 4475 29135 4525 29185
rect 4775 29135 4825 29185
rect 5075 29135 5125 29185
rect 5375 29135 5425 29185
rect 5675 29135 5725 29185
rect 5975 29135 6025 29185
rect 6275 29135 6325 29185
rect 6575 29135 6625 29185
rect 6875 29135 6925 29185
rect 7175 29135 7225 29185
rect 7475 29135 7525 29185
rect 7775 29135 7825 29185
rect 8075 29135 8125 29185
rect 8375 29135 8425 29185
rect 8675 29135 8725 29185
rect 8975 29135 9025 29185
rect 1775 28835 1825 28885
rect 2075 28835 2125 28885
rect 2375 28835 2425 28885
rect 2675 28835 2725 28885
rect 2975 28835 3025 28885
rect 3275 28835 3325 28885
rect 3575 28835 3625 28885
rect 3875 28835 3925 28885
rect 4175 28835 4225 28885
rect 4475 28835 4525 28885
rect 4775 28835 4825 28885
rect 5075 28835 5125 28885
rect 5375 28835 5425 28885
rect 5675 28835 5725 28885
rect 5975 28835 6025 28885
rect 6275 28835 6325 28885
rect 6575 28835 6625 28885
rect 6875 28835 6925 28885
rect 7175 28835 7225 28885
rect 7475 28835 7525 28885
rect 7775 28835 7825 28885
rect 8075 28835 8125 28885
rect 8375 28835 8425 28885
rect 8675 28835 8725 28885
rect 8975 28835 9025 28885
rect 1775 28535 1825 28585
rect 2075 28535 2125 28585
rect 2375 28535 2425 28585
rect 2675 28535 2725 28585
rect 2975 28535 3025 28585
rect 3275 28535 3325 28585
rect 3575 28535 3625 28585
rect 3875 28535 3925 28585
rect 4175 28535 4225 28585
rect 4475 28535 4525 28585
rect 4775 28535 4825 28585
rect 5075 28535 5125 28585
rect 5375 28535 5425 28585
rect 5675 28535 5725 28585
rect 5975 28535 6025 28585
rect 6275 28535 6325 28585
rect 6575 28535 6625 28585
rect 6875 28535 6925 28585
rect 7175 28535 7225 28585
rect 7475 28535 7525 28585
rect 7775 28535 7825 28585
rect 8075 28535 8125 28585
rect 8375 28535 8425 28585
rect 8675 28535 8725 28585
rect 8975 28535 9025 28585
rect 1775 28235 1825 28285
rect 2075 28235 2125 28285
rect 2375 28235 2425 28285
rect 2675 28235 2725 28285
rect 2975 28235 3025 28285
rect 3275 28235 3325 28285
rect 3575 28235 3625 28285
rect 3875 28235 3925 28285
rect 4175 28235 4225 28285
rect 4475 28235 4525 28285
rect 4775 28235 4825 28285
rect 5075 28235 5125 28285
rect 5375 28235 5425 28285
rect 5675 28235 5725 28285
rect 5975 28235 6025 28285
rect 6275 28235 6325 28285
rect 6575 28235 6625 28285
rect 6875 28235 6925 28285
rect 7175 28235 7225 28285
rect 7475 28235 7525 28285
rect 7775 28235 7825 28285
rect 8075 28235 8125 28285
rect 8375 28235 8425 28285
rect 8675 28235 8725 28285
rect 8975 28235 9025 28285
rect 1775 27935 1825 27985
rect 2075 27935 2125 27985
rect 2375 27935 2425 27985
rect 2675 27935 2725 27985
rect 2975 27935 3025 27985
rect 3275 27935 3325 27985
rect 3575 27935 3625 27985
rect 3875 27935 3925 27985
rect 4175 27935 4225 27985
rect 4475 27935 4525 27985
rect 4775 27935 4825 27985
rect 5075 27935 5125 27985
rect 5375 27935 5425 27985
rect 5675 27935 5725 27985
rect 5975 27935 6025 27985
rect 6275 27935 6325 27985
rect 6575 27935 6625 27985
rect 6875 27935 6925 27985
rect 7175 27935 7225 27985
rect 7475 27935 7525 27985
rect 7775 27935 7825 27985
rect 8075 27935 8125 27985
rect 8375 27935 8425 27985
rect 8675 27935 8725 27985
rect 8975 27935 9025 27985
rect 1775 27635 1825 27685
rect 2075 27635 2125 27685
rect 2375 27635 2425 27685
rect 2675 27635 2725 27685
rect 2975 27635 3025 27685
rect 3275 27635 3325 27685
rect 3575 27635 3625 27685
rect 3875 27635 3925 27685
rect 4175 27635 4225 27685
rect 4475 27635 4525 27685
rect 4775 27635 4825 27685
rect 5075 27635 5125 27685
rect 5375 27635 5425 27685
rect 5675 27635 5725 27685
rect 5975 27635 6025 27685
rect 6275 27635 6325 27685
rect 6575 27635 6625 27685
rect 6875 27635 6925 27685
rect 7175 27635 7225 27685
rect 7475 27635 7525 27685
rect 7775 27635 7825 27685
rect 8075 27635 8125 27685
rect 8375 27635 8425 27685
rect 8675 27635 8725 27685
rect 8975 27635 9025 27685
rect 1775 27335 1825 27385
rect 2075 27335 2125 27385
rect 2375 27335 2425 27385
rect 2675 27335 2725 27385
rect 2975 27335 3025 27385
rect 3275 27335 3325 27385
rect 3575 27335 3625 27385
rect 3875 27335 3925 27385
rect 4175 27335 4225 27385
rect 4475 27335 4525 27385
rect 4775 27335 4825 27385
rect 5075 27335 5125 27385
rect 5375 27335 5425 27385
rect 5675 27335 5725 27385
rect 5975 27335 6025 27385
rect 6275 27335 6325 27385
rect 6575 27335 6625 27385
rect 6875 27335 6925 27385
rect 7175 27335 7225 27385
rect 7475 27335 7525 27385
rect 7775 27335 7825 27385
rect 8075 27335 8125 27385
rect 8375 27335 8425 27385
rect 8675 27335 8725 27385
rect 8975 27335 9025 27385
rect 1775 27035 1825 27085
rect 2075 27035 2125 27085
rect 2375 27035 2425 27085
rect 2675 27035 2725 27085
rect 2975 27035 3025 27085
rect 3275 27035 3325 27085
rect 3575 27035 3625 27085
rect 3875 27035 3925 27085
rect 4175 27035 4225 27085
rect 4475 27035 4525 27085
rect 4775 27035 4825 27085
rect 5075 27035 5125 27085
rect 5375 27035 5425 27085
rect 5675 27035 5725 27085
rect 5975 27035 6025 27085
rect 6275 27035 6325 27085
rect 6575 27035 6625 27085
rect 6875 27035 6925 27085
rect 7175 27035 7225 27085
rect 7475 27035 7525 27085
rect 7775 27035 7825 27085
rect 8075 27035 8125 27085
rect 8375 27035 8425 27085
rect 8675 27035 8725 27085
rect 8975 27035 9025 27085
rect 1775 26735 1825 26785
rect 2075 26735 2125 26785
rect 2375 26735 2425 26785
rect 2675 26735 2725 26785
rect 2975 26735 3025 26785
rect 3275 26735 3325 26785
rect 3575 26735 3625 26785
rect 3875 26735 3925 26785
rect 4175 26735 4225 26785
rect 4475 26735 4525 26785
rect 4775 26735 4825 26785
rect 5075 26735 5125 26785
rect 5375 26735 5425 26785
rect 5675 26735 5725 26785
rect 5975 26735 6025 26785
rect 6275 26735 6325 26785
rect 6575 26735 6625 26785
rect 6875 26735 6925 26785
rect 7175 26735 7225 26785
rect 7475 26735 7525 26785
rect 7775 26735 7825 26785
rect 8075 26735 8125 26785
rect 8375 26735 8425 26785
rect 8675 26735 8725 26785
rect 8975 26735 9025 26785
rect 1775 26435 1825 26485
rect 2075 26435 2125 26485
rect 2375 26435 2425 26485
rect 2675 26435 2725 26485
rect 2975 26435 3025 26485
rect 3275 26435 3325 26485
rect 3575 26435 3625 26485
rect 3875 26435 3925 26485
rect 4175 26435 4225 26485
rect 4475 26435 4525 26485
rect 4775 26435 4825 26485
rect 5075 26435 5125 26485
rect 5375 26435 5425 26485
rect 5675 26435 5725 26485
rect 5975 26435 6025 26485
rect 6275 26435 6325 26485
rect 6575 26435 6625 26485
rect 6875 26435 6925 26485
rect 7175 26435 7225 26485
rect 7475 26435 7525 26485
rect 7775 26435 7825 26485
rect 8075 26435 8125 26485
rect 8375 26435 8425 26485
rect 8675 26435 8725 26485
rect 8975 26435 9025 26485
rect 1775 26135 1825 26185
rect 2075 26135 2125 26185
rect 2375 26135 2425 26185
rect 2675 26135 2725 26185
rect 2975 26135 3025 26185
rect 3275 26135 3325 26185
rect 3575 26135 3625 26185
rect 3875 26135 3925 26185
rect 4175 26135 4225 26185
rect 4475 26135 4525 26185
rect 4775 26135 4825 26185
rect 5075 26135 5125 26185
rect 5375 26135 5425 26185
rect 5675 26135 5725 26185
rect 5975 26135 6025 26185
rect 6275 26135 6325 26185
rect 6575 26135 6625 26185
rect 6875 26135 6925 26185
rect 7175 26135 7225 26185
rect 7475 26135 7525 26185
rect 7775 26135 7825 26185
rect 8075 26135 8125 26185
rect 8375 26135 8425 26185
rect 8675 26135 8725 26185
rect 8975 26135 9025 26185
rect 1775 25835 1825 25885
rect 2075 25835 2125 25885
rect 2375 25835 2425 25885
rect 2675 25835 2725 25885
rect 2975 25835 3025 25885
rect 3275 25835 3325 25885
rect 3575 25835 3625 25885
rect 3875 25835 3925 25885
rect 4175 25835 4225 25885
rect 4475 25835 4525 25885
rect 4775 25835 4825 25885
rect 5075 25835 5125 25885
rect 5375 25835 5425 25885
rect 5675 25835 5725 25885
rect 5975 25835 6025 25885
rect 6275 25835 6325 25885
rect 6575 25835 6625 25885
rect 6875 25835 6925 25885
rect 7175 25835 7225 25885
rect 7475 25835 7525 25885
rect 7775 25835 7825 25885
rect 8075 25835 8125 25885
rect 8375 25835 8425 25885
rect 8675 25835 8725 25885
rect 8975 25835 9025 25885
rect 1775 25535 1825 25585
rect 2075 25535 2125 25585
rect 2375 25535 2425 25585
rect 2675 25535 2725 25585
rect 2975 25535 3025 25585
rect 3275 25535 3325 25585
rect 3575 25535 3625 25585
rect 3875 25535 3925 25585
rect 4175 25535 4225 25585
rect 4475 25535 4525 25585
rect 4775 25535 4825 25585
rect 5075 25535 5125 25585
rect 5375 25535 5425 25585
rect 5675 25535 5725 25585
rect 5975 25535 6025 25585
rect 6275 25535 6325 25585
rect 6575 25535 6625 25585
rect 6875 25535 6925 25585
rect 7175 25535 7225 25585
rect 7475 25535 7525 25585
rect 7775 25535 7825 25585
rect 8075 25535 8125 25585
rect 8375 25535 8425 25585
rect 8675 25535 8725 25585
rect 8975 25535 9025 25585
rect 1775 25235 1825 25285
rect 2075 25235 2125 25285
rect 2375 25235 2425 25285
rect 2675 25235 2725 25285
rect 2975 25235 3025 25285
rect 3275 25235 3325 25285
rect 3575 25235 3625 25285
rect 3875 25235 3925 25285
rect 4175 25235 4225 25285
rect 4475 25235 4525 25285
rect 4775 25235 4825 25285
rect 5075 25235 5125 25285
rect 5375 25235 5425 25285
rect 5675 25235 5725 25285
rect 5975 25235 6025 25285
rect 6275 25235 6325 25285
rect 6575 25235 6625 25285
rect 6875 25235 6925 25285
rect 7175 25235 7225 25285
rect 7475 25235 7525 25285
rect 7775 25235 7825 25285
rect 8075 25235 8125 25285
rect 8375 25235 8425 25285
rect 8675 25235 8725 25285
rect 8975 25235 9025 25285
rect 1775 24935 1825 24985
rect 2075 24935 2125 24985
rect 2375 24935 2425 24985
rect 2675 24935 2725 24985
rect 2975 24935 3025 24985
rect 3275 24935 3325 24985
rect 3575 24935 3625 24985
rect 3875 24935 3925 24985
rect 4175 24935 4225 24985
rect 4475 24935 4525 24985
rect 4775 24935 4825 24985
rect 5075 24935 5125 24985
rect 5375 24935 5425 24985
rect 5675 24935 5725 24985
rect 5975 24935 6025 24985
rect 6275 24935 6325 24985
rect 6575 24935 6625 24985
rect 6875 24935 6925 24985
rect 7175 24935 7225 24985
rect 7475 24935 7525 24985
rect 7775 24935 7825 24985
rect 8075 24935 8125 24985
rect 8375 24935 8425 24985
rect 8675 24935 8725 24985
rect 8975 24935 9025 24985
rect 1775 24635 1825 24685
rect 2075 24635 2125 24685
rect 2375 24635 2425 24685
rect 2675 24635 2725 24685
rect 2975 24635 3025 24685
rect 3275 24635 3325 24685
rect 3575 24635 3625 24685
rect 3875 24635 3925 24685
rect 4175 24635 4225 24685
rect 4475 24635 4525 24685
rect 4775 24635 4825 24685
rect 5075 24635 5125 24685
rect 5375 24635 5425 24685
rect 5675 24635 5725 24685
rect 5975 24635 6025 24685
rect 6275 24635 6325 24685
rect 6575 24635 6625 24685
rect 6875 24635 6925 24685
rect 7175 24635 7225 24685
rect 7475 24635 7525 24685
rect 7775 24635 7825 24685
rect 8075 24635 8125 24685
rect 8375 24635 8425 24685
rect 8675 24635 8725 24685
rect 8975 24635 9025 24685
rect 1775 24335 1825 24385
rect 2075 24335 2125 24385
rect 2375 24335 2425 24385
rect 2675 24335 2725 24385
rect 2975 24335 3025 24385
rect 3275 24335 3325 24385
rect 3575 24335 3625 24385
rect 3875 24335 3925 24385
rect 4175 24335 4225 24385
rect 4475 24335 4525 24385
rect 4775 24335 4825 24385
rect 5075 24335 5125 24385
rect 5375 24335 5425 24385
rect 5675 24335 5725 24385
rect 5975 24335 6025 24385
rect 6275 24335 6325 24385
rect 6575 24335 6625 24385
rect 6875 24335 6925 24385
rect 7175 24335 7225 24385
rect 7475 24335 7525 24385
rect 7775 24335 7825 24385
rect 8075 24335 8125 24385
rect 8375 24335 8425 24385
rect 8675 24335 8725 24385
rect 8975 24335 9025 24385
rect 1775 24035 1825 24085
rect 2075 24035 2125 24085
rect 2375 24035 2425 24085
rect 2675 24035 2725 24085
rect 2975 24035 3025 24085
rect 3275 24035 3325 24085
rect 3575 24035 3625 24085
rect 3875 24035 3925 24085
rect 4175 24035 4225 24085
rect 4475 24035 4525 24085
rect 4775 24035 4825 24085
rect 5075 24035 5125 24085
rect 5375 24035 5425 24085
rect 5675 24035 5725 24085
rect 5975 24035 6025 24085
rect 6275 24035 6325 24085
rect 6575 24035 6625 24085
rect 6875 24035 6925 24085
rect 7175 24035 7225 24085
rect 7475 24035 7525 24085
rect 7775 24035 7825 24085
rect 8075 24035 8125 24085
rect 8375 24035 8425 24085
rect 8675 24035 8725 24085
rect 8975 24035 9025 24085
rect 1775 23735 1825 23785
rect 2075 23735 2125 23785
rect 2375 23735 2425 23785
rect 2675 23735 2725 23785
rect 2975 23735 3025 23785
rect 3275 23735 3325 23785
rect 3575 23735 3625 23785
rect 3875 23735 3925 23785
rect 4175 23735 4225 23785
rect 4475 23735 4525 23785
rect 4775 23735 4825 23785
rect 5075 23735 5125 23785
rect 5375 23735 5425 23785
rect 5675 23735 5725 23785
rect 5975 23735 6025 23785
rect 6275 23735 6325 23785
rect 6575 23735 6625 23785
rect 6875 23735 6925 23785
rect 7175 23735 7225 23785
rect 7475 23735 7525 23785
rect 7775 23735 7825 23785
rect 8075 23735 8125 23785
rect 8375 23735 8425 23785
rect 8675 23735 8725 23785
rect 8975 23735 9025 23785
rect 1775 23435 1825 23485
rect 2075 23435 2125 23485
rect 2375 23435 2425 23485
rect 2675 23435 2725 23485
rect 2975 23435 3025 23485
rect 3275 23435 3325 23485
rect 3575 23435 3625 23485
rect 3875 23435 3925 23485
rect 4175 23435 4225 23485
rect 4475 23435 4525 23485
rect 4775 23435 4825 23485
rect 5075 23435 5125 23485
rect 5375 23435 5425 23485
rect 5675 23435 5725 23485
rect 5975 23435 6025 23485
rect 6275 23435 6325 23485
rect 6575 23435 6625 23485
rect 6875 23435 6925 23485
rect 7175 23435 7225 23485
rect 7475 23435 7525 23485
rect 7775 23435 7825 23485
rect 8075 23435 8125 23485
rect 8375 23435 8425 23485
rect 8675 23435 8725 23485
rect 8975 23435 9025 23485
rect 155 20735 205 20785
rect 395 20735 445 20785
rect 635 20735 685 20785
rect 875 20735 925 20785
rect 1115 20735 1165 20785
rect 1355 20735 1405 20785
rect 1595 20735 1645 20785
rect 1835 20735 1885 20785
rect 2075 20735 2125 20785
rect 2315 20735 2365 20785
rect 2555 20735 2605 20785
rect 2795 20735 2845 20785
rect 3035 20735 3085 20785
rect 3275 20735 3325 20785
rect 4655 20735 4705 20785
rect 4895 20735 4945 20785
rect 5135 20735 5185 20785
rect 5375 20735 5425 20785
rect 5615 20735 5665 20785
rect 5855 20735 5905 20785
rect 6095 20735 6145 20785
rect 7475 20735 7525 20785
rect 7715 20735 7765 20785
rect 7955 20735 8005 20785
rect 8195 20735 8245 20785
rect 8435 20735 8485 20785
rect 8675 20735 8725 20785
rect 8915 20735 8965 20785
rect 9155 20735 9205 20785
rect 9395 20735 9445 20785
rect 9635 20735 9685 20785
rect 9875 20735 9925 20785
rect 10115 20735 10165 20785
rect 10355 20735 10405 20785
rect 10595 20735 10645 20785
rect 155 20585 205 20635
rect 395 20585 445 20635
rect 635 20585 685 20635
rect 875 20585 925 20635
rect 1115 20585 1165 20635
rect 1355 20585 1405 20635
rect 1595 20585 1645 20635
rect 1835 20585 1885 20635
rect 2075 20585 2125 20635
rect 2315 20585 2365 20635
rect 2555 20585 2605 20635
rect 2795 20585 2845 20635
rect 3035 20585 3085 20635
rect 3275 20585 3325 20635
rect 4655 20585 4705 20635
rect 4895 20585 4945 20635
rect 5135 20585 5185 20635
rect 5375 20585 5425 20635
rect 5615 20585 5665 20635
rect 5855 20585 5905 20635
rect 6095 20585 6145 20635
rect 7475 20585 7525 20635
rect 7715 20585 7765 20635
rect 7955 20585 8005 20635
rect 8195 20585 8245 20635
rect 8435 20585 8485 20635
rect 8675 20585 8725 20635
rect 8915 20585 8965 20635
rect 9155 20585 9205 20635
rect 9395 20585 9445 20635
rect 9635 20585 9685 20635
rect 9875 20585 9925 20635
rect 10115 20585 10165 20635
rect 10355 20585 10405 20635
rect 10595 20585 10645 20635
rect 605 20045 655 20095
rect 755 20045 805 20095
rect 1055 20045 1105 20095
rect 1385 20045 1435 20095
rect 1685 20045 1735 20095
rect 1985 20045 2035 20095
rect 2285 20045 2335 20095
rect 2585 20045 2635 20095
rect 2885 20045 2935 20095
rect 3185 20045 3235 20095
rect 4655 20045 4705 20095
rect 5315 20045 5365 20095
rect 5465 20045 5515 20095
rect 6095 20045 6145 20095
rect 7565 20045 7615 20095
rect 7865 20045 7915 20095
rect 8165 20045 8215 20095
rect 8465 20045 8515 20095
rect 8765 20045 8815 20095
rect 9065 20045 9115 20095
rect 9365 20045 9415 20095
rect 9665 20045 9715 20095
rect 9965 20045 10045 20095
rect 10145 20045 10195 20095
rect 605 19895 655 19945
rect 755 19895 805 19945
rect 1055 19895 1105 19945
rect 1385 19895 1435 19945
rect 1685 19895 1735 19945
rect 1985 19895 2035 19945
rect 2285 19895 2335 19945
rect 2585 19895 2635 19945
rect 2885 19895 2935 19945
rect 3185 19895 3235 19945
rect 4655 19895 4705 19945
rect 5315 19895 5365 19945
rect 5465 19895 5515 19945
rect 6095 19895 6145 19945
rect 7565 19895 7615 19945
rect 7865 19895 7915 19945
rect 8165 19895 8215 19945
rect 8465 19895 8515 19945
rect 8765 19895 8815 19945
rect 9065 19895 9115 19945
rect 9365 19895 9415 19945
rect 9665 19895 9715 19945
rect 9995 19895 10045 19945
rect 10145 19895 10195 19945
rect 605 19745 655 19795
rect 755 19745 805 19795
rect 1055 19745 1105 19795
rect 1385 19745 1435 19795
rect 1685 19745 1735 19795
rect 1985 19745 2035 19795
rect 2285 19745 2335 19795
rect 2585 19745 2635 19795
rect 2885 19745 2935 19795
rect 3185 19745 3235 19795
rect 4655 19745 4705 19795
rect 5315 19745 5365 19795
rect 5465 19745 5515 19795
rect 6095 19745 6145 19795
rect 7565 19745 7615 19795
rect 7865 19745 7915 19795
rect 8165 19745 8215 19795
rect 8465 19745 8515 19795
rect 8765 19745 8815 19795
rect 9065 19745 9115 19795
rect 9365 19745 9415 19795
rect 9665 19745 9715 19795
rect 9995 19745 10045 19795
rect 10145 19745 10195 19795
rect 65 19265 115 19315
rect 215 19265 265 19315
rect 10535 19265 10585 19315
rect 10685 19265 10735 19315
rect 65 19025 115 19075
rect 215 19025 265 19075
rect 10535 19025 10585 19075
rect 10685 19025 10735 19075
rect 65 18785 115 18835
rect 215 18785 265 18835
rect 10535 18785 10585 18835
rect 10685 18785 10735 18835
rect 605 18095 655 18145
rect 755 18095 805 18145
rect 1385 18095 1435 18145
rect 1685 18095 1735 18145
rect 1985 18095 2035 18145
rect 2285 18095 2335 18145
rect 2585 18095 2635 18145
rect 2885 18095 2935 18145
rect 3185 18095 3235 18145
rect 4655 18095 4705 18145
rect 5315 18095 5365 18145
rect 5465 18095 5515 18145
rect 6095 18095 6145 18145
rect 7565 18095 7615 18145
rect 7865 18095 7915 18145
rect 8165 18095 8215 18145
rect 8465 18095 8515 18145
rect 8765 18095 8815 18145
rect 9065 18095 9115 18145
rect 9365 18095 9415 18145
rect 9995 18095 10045 18145
rect 10145 18095 10195 18145
rect 605 17945 655 17995
rect 755 17945 805 17995
rect 1385 17945 1435 17995
rect 1685 17945 1735 17995
rect 1985 17945 2035 17995
rect 2285 17945 2335 17995
rect 2585 17945 2635 17995
rect 2885 17945 2935 17995
rect 3185 17945 3235 17995
rect 4655 17945 4705 17995
rect 5315 17945 5365 17995
rect 5465 17945 5515 17995
rect 6095 17945 6145 17995
rect 7565 17945 7615 17995
rect 7865 17945 7915 17995
rect 8165 17945 8215 17995
rect 8465 17945 8515 17995
rect 8765 17945 8815 17995
rect 9065 17945 9115 17995
rect 9365 17945 9415 17995
rect 9995 17945 10045 17995
rect 10145 17945 10195 17995
rect 605 17795 655 17845
rect 755 17795 805 17845
rect 1385 17795 1435 17845
rect 1685 17795 1735 17845
rect 1985 17795 2035 17845
rect 2285 17795 2335 17845
rect 2585 17795 2635 17845
rect 2885 17795 2935 17845
rect 3185 17795 3235 17845
rect 4655 17795 4705 17845
rect 5315 17795 5365 17845
rect 5465 17795 5515 17845
rect 6095 17795 6145 17845
rect 7565 17795 7615 17845
rect 7865 17795 7915 17845
rect 8165 17795 8215 17845
rect 8465 17795 8515 17845
rect 8765 17795 8815 17845
rect 9065 17795 9115 17845
rect 9365 17795 9415 17845
rect 9995 17795 10045 17845
rect 10145 17795 10195 17845
rect 65 17345 115 17395
rect 215 17345 265 17395
rect 10535 17345 10585 17395
rect 10685 17345 10735 17395
rect 65 17105 115 17155
rect 215 17105 265 17155
rect 10535 17105 10585 17155
rect 10685 17105 10735 17155
rect 65 16865 115 16915
rect 215 16865 265 16915
rect 10535 16865 10585 16915
rect 10685 16865 10735 16915
rect 605 16145 655 16195
rect 755 16145 805 16195
rect 1385 16145 1435 16195
rect 1685 16145 1735 16195
rect 1985 16145 2035 16195
rect 2285 16145 2335 16195
rect 2585 16145 2635 16195
rect 2885 16145 2935 16195
rect 3185 16145 3235 16195
rect 4655 16145 4705 16195
rect 5315 16145 5365 16195
rect 5465 16145 5515 16195
rect 6095 16145 6145 16195
rect 7565 16145 7615 16195
rect 7865 16145 7915 16195
rect 8165 16145 8215 16195
rect 8465 16145 8515 16195
rect 8765 16145 8815 16195
rect 9065 16145 9115 16195
rect 9365 16145 9415 16195
rect 9995 16145 10045 16195
rect 10145 16145 10195 16195
rect 605 15995 655 16045
rect 755 15995 805 16045
rect 1385 15995 1435 16045
rect 1685 15995 1735 16045
rect 1985 15995 2035 16045
rect 2285 15995 2335 16045
rect 2585 15995 2635 16045
rect 2885 15995 2935 16045
rect 3185 15995 3235 16045
rect 4655 15995 4705 16045
rect 5315 15995 5365 16045
rect 5465 15995 5515 16045
rect 6095 15995 6145 16045
rect 7565 15995 7615 16045
rect 7865 15995 7915 16045
rect 8165 15995 8215 16045
rect 8465 15995 8515 16045
rect 8765 15995 8815 16045
rect 9065 15995 9115 16045
rect 9365 15995 9415 16045
rect 9995 15995 10045 16045
rect 10145 15995 10195 16045
rect 605 15845 655 15895
rect 755 15845 805 15895
rect 1385 15845 1435 15895
rect 1685 15845 1735 15895
rect 1985 15845 2035 15895
rect 2285 15845 2335 15895
rect 2585 15845 2635 15895
rect 2885 15845 2935 15895
rect 3185 15845 3235 15895
rect 4655 15845 4705 15895
rect 5315 15845 5365 15895
rect 5465 15845 5515 15895
rect 6095 15845 6145 15895
rect 7565 15845 7615 15895
rect 7865 15845 7915 15895
rect 8165 15845 8215 15895
rect 8465 15845 8515 15895
rect 8765 15845 8815 15895
rect 9065 15845 9115 15895
rect 9365 15845 9415 15895
rect 9995 15845 10045 15895
rect 10145 15845 10195 15895
rect 65 15395 115 15445
rect 215 15395 265 15445
rect 10535 15395 10585 15445
rect 10685 15395 10735 15445
rect 65 15155 115 15205
rect 215 15155 265 15205
rect 10535 15155 10585 15205
rect 10685 15155 10735 15205
rect 65 14915 115 14965
rect 215 14915 265 14965
rect 10535 14915 10585 14965
rect 10685 14915 10735 14965
rect 605 14195 655 14245
rect 755 14195 805 14245
rect 1385 14195 1435 14245
rect 1685 14195 1735 14245
rect 1985 14195 2035 14245
rect 2285 14195 2335 14245
rect 2585 14195 2635 14245
rect 2885 14195 2935 14245
rect 3185 14195 3235 14245
rect 4655 14195 4705 14245
rect 5315 14195 5365 14245
rect 5465 14195 5515 14245
rect 6095 14195 6145 14245
rect 7565 14195 7615 14245
rect 7865 14195 7915 14245
rect 8165 14195 8215 14245
rect 8465 14195 8515 14245
rect 8765 14195 8815 14245
rect 9065 14195 9115 14245
rect 9365 14195 9415 14245
rect 9995 14195 10045 14245
rect 10145 14195 10195 14245
rect 605 14045 655 14095
rect 755 14045 805 14095
rect 1385 14045 1435 14095
rect 1685 14045 1735 14095
rect 1985 14045 2035 14095
rect 2285 14045 2335 14095
rect 2585 14045 2635 14095
rect 2885 14045 2935 14095
rect 3185 14045 3235 14095
rect 4655 14045 4705 14095
rect 5315 14045 5365 14095
rect 5465 14045 5515 14095
rect 6095 14045 6145 14095
rect 7565 14045 7615 14095
rect 7865 14045 7915 14095
rect 8165 14045 8215 14095
rect 8465 14045 8515 14095
rect 8765 14045 8815 14095
rect 9065 14045 9115 14095
rect 9365 14045 9415 14095
rect 9995 14045 10045 14095
rect 10145 14045 10195 14095
rect 605 13895 655 13945
rect 755 13895 805 13945
rect 1385 13895 1435 13945
rect 1685 13895 1735 13945
rect 1985 13895 2035 13945
rect 2285 13895 2335 13945
rect 2585 13895 2635 13945
rect 2885 13895 2935 13945
rect 3185 13895 3235 13945
rect 4655 13895 4705 13945
rect 5315 13895 5365 13945
rect 5465 13895 5515 13945
rect 6095 13895 6145 13945
rect 7565 13895 7615 13945
rect 7865 13895 7915 13945
rect 8165 13895 8215 13945
rect 8465 13895 8515 13945
rect 8765 13895 8815 13945
rect 9065 13895 9115 13945
rect 9365 13895 9415 13945
rect 9995 13895 10045 13945
rect 10145 13895 10195 13945
rect 155 13355 205 13405
rect 395 13355 445 13405
rect 635 13355 685 13405
rect 1355 13355 1405 13405
rect 1595 13355 1645 13405
rect 1835 13355 1885 13405
rect 2075 13355 2125 13405
rect 2315 13355 2365 13405
rect 2555 13355 2605 13405
rect 2795 13355 2845 13405
rect 3035 13355 3085 13405
rect 3275 13355 3325 13405
rect 4625 13355 4675 13405
rect 5315 13355 5365 13405
rect 6065 13355 6115 13405
rect 7475 13355 7525 13405
rect 7715 13355 7765 13405
rect 7955 13355 8005 13405
rect 8195 13355 8245 13405
rect 8435 13355 8485 13405
rect 8675 13355 8725 13405
rect 8915 13355 8965 13405
rect 9155 13355 9205 13405
rect 9395 13355 9445 13405
rect 10115 13355 10165 13405
rect 10355 13355 10405 13405
rect 10595 13355 10645 13405
rect 155 13205 205 13255
rect 395 13205 445 13255
rect 635 13205 685 13255
rect 1355 13205 1405 13255
rect 1595 13205 1645 13255
rect 1835 13205 1885 13255
rect 2075 13205 2125 13255
rect 2315 13205 2365 13255
rect 2555 13205 2605 13255
rect 2795 13205 2845 13255
rect 3035 13205 3085 13255
rect 3275 13205 3325 13255
rect 4625 13205 4675 13255
rect 5315 13205 5365 13255
rect 6065 13205 6115 13255
rect 7475 13205 7525 13255
rect 7715 13205 7765 13255
rect 7955 13205 8005 13255
rect 8195 13205 8245 13255
rect 8435 13205 8485 13255
rect 8675 13205 8725 13255
rect 8915 13205 8965 13255
rect 9155 13205 9205 13255
rect 9395 13205 9445 13255
rect 10115 13205 10165 13255
rect 10355 13205 10405 13255
rect 10595 13205 10645 13255
rect 155 12845 205 12895
rect 395 12845 445 12895
rect 635 12845 685 12895
rect 1355 12845 1405 12895
rect 1595 12845 1645 12895
rect 1835 12845 1885 12895
rect 2075 12845 2125 12895
rect 2315 12845 2365 12895
rect 2555 12845 2605 12895
rect 2795 12845 2845 12895
rect 3035 12845 3085 12895
rect 3275 12845 3325 12895
rect 4625 12845 4675 12895
rect 5315 12845 5365 12895
rect 6065 12845 6115 12895
rect 7475 12845 7525 12895
rect 7715 12845 7765 12895
rect 7955 12845 8005 12895
rect 8195 12845 8245 12895
rect 8435 12845 8485 12895
rect 8675 12845 8725 12895
rect 8915 12845 8965 12895
rect 9155 12845 9205 12895
rect 9395 12845 9445 12895
rect 10115 12845 10165 12895
rect 10355 12845 10405 12895
rect 10595 12845 10645 12895
rect 155 12695 205 12745
rect 395 12695 445 12745
rect 635 12695 685 12745
rect 1355 12695 1405 12745
rect 1595 12695 1645 12745
rect 1835 12695 1885 12745
rect 2075 12695 2125 12745
rect 2315 12695 2365 12745
rect 2555 12695 2605 12745
rect 2795 12695 2845 12745
rect 3035 12695 3085 12745
rect 3275 12695 3325 12745
rect 4625 12695 4675 12745
rect 5315 12695 5365 12745
rect 6065 12695 6115 12745
rect 7475 12695 7525 12745
rect 7715 12695 7765 12745
rect 7955 12695 8005 12745
rect 8195 12695 8245 12745
rect 8435 12695 8485 12745
rect 8675 12695 8725 12745
rect 8915 12695 8965 12745
rect 9155 12695 9205 12745
rect 9395 12695 9445 12745
rect 10115 12695 10165 12745
rect 10355 12695 10405 12745
rect 10595 12695 10645 12745
rect 155 12005 205 12055
rect 395 12005 445 12055
rect 635 12005 685 12055
rect 875 12005 925 12055
rect 1115 12005 1165 12055
rect 1355 12005 1405 12055
rect 1595 12005 1645 12055
rect 1835 12005 1885 12055
rect 2075 12005 2125 12055
rect 2315 12005 2365 12055
rect 2555 12005 2605 12055
rect 2795 12005 2845 12055
rect 3035 12005 3085 12055
rect 3275 12005 3325 12055
rect 4625 12005 4675 12055
rect 5315 12005 5365 12055
rect 6065 12005 6115 12055
rect 7475 12005 7525 12055
rect 7715 12005 7765 12055
rect 7955 12005 8005 12055
rect 8195 12005 8245 12055
rect 8435 12005 8485 12055
rect 8675 12005 8725 12055
rect 8915 12005 8965 12055
rect 9155 12005 9205 12055
rect 9395 12005 9445 12055
rect 9635 12005 9685 12055
rect 9875 12005 9925 12055
rect 10115 12005 10165 12055
rect 10355 12005 10405 12055
rect 10595 12005 10645 12055
rect 155 11855 205 11905
rect 395 11855 445 11905
rect 635 11855 685 11905
rect 875 11855 925 11905
rect 1115 11855 1165 11905
rect 1355 11855 1405 11905
rect 1595 11855 1645 11905
rect 1835 11855 1885 11905
rect 2075 11855 2125 11905
rect 2315 11855 2365 11905
rect 2555 11855 2605 11905
rect 2795 11855 2845 11905
rect 3035 11855 3085 11905
rect 3275 11855 3325 11905
rect 4625 11855 4675 11905
rect 5315 11855 5365 11905
rect 6065 11855 6115 11905
rect 7475 11855 7525 11905
rect 7715 11855 7765 11905
rect 7955 11855 8005 11905
rect 8195 11855 8245 11905
rect 8435 11855 8485 11905
rect 8675 11855 8725 11905
rect 8915 11855 8965 11905
rect 9155 11855 9205 11905
rect 9395 11855 9445 11905
rect 9635 11855 9685 11905
rect 9875 11855 9925 11905
rect 10115 11855 10165 11905
rect 10355 11855 10405 11905
rect 10595 11855 10645 11905
rect 155 11495 205 11545
rect 395 11495 445 11545
rect 635 11495 685 11545
rect 875 11495 925 11545
rect 1115 11495 1165 11545
rect 1355 11495 1405 11545
rect 1595 11495 1645 11545
rect 1835 11495 1885 11545
rect 2075 11495 2125 11545
rect 2315 11495 2365 11545
rect 2555 11495 2605 11545
rect 2795 11495 2845 11545
rect 3035 11495 3085 11545
rect 3275 11495 3325 11545
rect 4625 11495 4675 11545
rect 5315 11495 5365 11545
rect 6065 11495 6115 11545
rect 7475 11495 7525 11545
rect 7715 11495 7765 11545
rect 7955 11495 8005 11545
rect 8195 11495 8245 11545
rect 8435 11495 8485 11545
rect 8675 11495 8725 11545
rect 8915 11495 8965 11545
rect 9155 11495 9205 11545
rect 9395 11495 9445 11545
rect 9635 11495 9685 11545
rect 9875 11495 9925 11545
rect 10115 11495 10165 11545
rect 10355 11495 10405 11545
rect 10595 11495 10645 11545
rect 155 11345 205 11395
rect 395 11345 445 11395
rect 635 11345 685 11395
rect 875 11345 925 11395
rect 1115 11345 1165 11395
rect 1355 11345 1405 11395
rect 1595 11345 1645 11395
rect 1835 11345 1885 11395
rect 2075 11345 2125 11395
rect 2315 11345 2365 11395
rect 2555 11345 2605 11395
rect 2795 11345 2845 11395
rect 3035 11345 3085 11395
rect 3275 11345 3325 11395
rect 4625 11345 4675 11395
rect 5315 11345 5365 11395
rect 6065 11345 6115 11395
rect 7475 11345 7525 11395
rect 7715 11345 7765 11395
rect 7955 11345 8005 11395
rect 8195 11345 8245 11395
rect 8435 11345 8485 11395
rect 8675 11345 8725 11395
rect 8915 11345 8965 11395
rect 9155 11345 9205 11395
rect 9395 11345 9445 11395
rect 9635 11345 9685 11395
rect 9875 11345 9925 11395
rect 10115 11345 10165 11395
rect 10355 11345 10405 11395
rect 10595 11345 10645 11395
rect 605 10805 655 10855
rect 755 10805 805 10855
rect 1385 10805 1435 10855
rect 1685 10805 1735 10855
rect 1985 10805 2035 10855
rect 2285 10805 2335 10855
rect 2585 10805 2635 10855
rect 2885 10805 2935 10855
rect 3185 10805 3235 10855
rect 4475 10805 4525 10855
rect 5315 10805 5365 10855
rect 5465 10805 5515 10855
rect 6275 10805 6325 10855
rect 7565 10805 7615 10855
rect 7865 10805 7915 10855
rect 8165 10805 8215 10855
rect 8465 10805 8515 10855
rect 8765 10805 8815 10855
rect 9065 10805 9115 10855
rect 9365 10805 9415 10855
rect 9995 10805 10045 10855
rect 10145 10805 10195 10855
rect 605 10655 655 10705
rect 755 10655 805 10705
rect 1385 10655 1435 10705
rect 1685 10655 1735 10705
rect 1985 10655 2035 10705
rect 2285 10655 2335 10705
rect 2585 10655 2635 10705
rect 2885 10655 2935 10705
rect 3185 10655 3235 10705
rect 4475 10655 4525 10705
rect 5315 10655 5365 10705
rect 5465 10655 5515 10705
rect 6275 10655 6325 10705
rect 7565 10655 7615 10705
rect 7865 10655 7915 10705
rect 8165 10655 8215 10705
rect 8465 10655 8515 10705
rect 8765 10655 8815 10705
rect 9065 10655 9115 10705
rect 9365 10655 9415 10705
rect 9995 10655 10045 10705
rect 10145 10655 10195 10705
rect 605 10505 655 10555
rect 755 10505 805 10555
rect 1385 10505 1435 10555
rect 1685 10505 1735 10555
rect 1985 10505 2035 10555
rect 2285 10505 2335 10555
rect 2585 10505 2635 10555
rect 2885 10505 2935 10555
rect 3185 10505 3235 10555
rect 4475 10505 4525 10555
rect 5315 10505 5365 10555
rect 5465 10505 5515 10555
rect 6275 10505 6325 10555
rect 7565 10505 7615 10555
rect 7865 10505 7915 10555
rect 8165 10505 8215 10555
rect 8465 10505 8515 10555
rect 8765 10505 8815 10555
rect 9065 10505 9115 10555
rect 9365 10505 9415 10555
rect 9995 10505 10045 10555
rect 10145 10505 10195 10555
rect 65 10025 115 10075
rect 215 10025 265 10075
rect 10535 10025 10585 10075
rect 10685 10025 10735 10075
rect 65 9785 115 9835
rect 215 9785 265 9835
rect 10535 9785 10585 9835
rect 10685 9785 10735 9835
rect 65 9545 115 9595
rect 215 9545 265 9595
rect 10535 9545 10585 9595
rect 10685 9545 10735 9595
rect 605 8855 655 8905
rect 755 8855 805 8905
rect 1385 8855 1435 8905
rect 1685 8855 1735 8905
rect 1985 8855 2035 8905
rect 2285 8855 2335 8905
rect 2585 8855 2635 8905
rect 2885 8855 2935 8905
rect 3185 8855 3235 8905
rect 4475 8855 4525 8905
rect 5315 8855 5365 8905
rect 5465 8855 5515 8905
rect 6275 8855 6325 8905
rect 7565 8855 7615 8905
rect 7865 8855 7915 8905
rect 8165 8855 8215 8905
rect 8465 8855 8515 8905
rect 8765 8855 8815 8905
rect 9065 8855 9115 8905
rect 9365 8855 9415 8905
rect 9995 8855 10045 8905
rect 10145 8855 10195 8905
rect 605 8705 655 8755
rect 755 8705 805 8755
rect 1385 8705 1435 8755
rect 1685 8705 1735 8755
rect 1985 8705 2035 8755
rect 2285 8705 2335 8755
rect 2585 8705 2635 8755
rect 2885 8705 2935 8755
rect 3185 8705 3235 8755
rect 4475 8705 4525 8755
rect 5315 8705 5365 8755
rect 5465 8705 5515 8755
rect 6275 8705 6325 8755
rect 7565 8705 7615 8755
rect 7865 8705 7915 8755
rect 8165 8705 8215 8755
rect 8465 8705 8515 8755
rect 8765 8705 8815 8755
rect 9065 8705 9115 8755
rect 9365 8705 9415 8755
rect 9995 8705 10045 8755
rect 10145 8705 10195 8755
rect 605 8555 655 8605
rect 755 8555 805 8605
rect 1385 8555 1435 8605
rect 1685 8555 1735 8605
rect 1985 8555 2035 8605
rect 2285 8555 2335 8605
rect 2585 8555 2635 8605
rect 2885 8555 2935 8605
rect 3185 8555 3235 8605
rect 4475 8555 4525 8605
rect 5315 8555 5365 8605
rect 5465 8555 5515 8605
rect 6275 8555 6325 8605
rect 7565 8555 7615 8605
rect 7865 8555 7915 8605
rect 8165 8555 8215 8605
rect 8465 8555 8515 8605
rect 8765 8555 8815 8605
rect 9065 8555 9115 8605
rect 9365 8555 9415 8605
rect 9995 8555 10045 8605
rect 10145 8555 10195 8605
rect 65 8105 115 8155
rect 215 8105 265 8155
rect 10535 8105 10585 8155
rect 10685 8105 10735 8155
rect 65 7865 115 7915
rect 215 7865 265 7915
rect 10535 7865 10585 7915
rect 10685 7865 10735 7915
rect 65 7625 115 7675
rect 215 7625 265 7675
rect 10535 7625 10585 7675
rect 10685 7625 10735 7675
rect 605 6905 655 6955
rect 755 6905 805 6955
rect 1385 6905 1435 6955
rect 1685 6905 1735 6955
rect 1985 6905 2035 6955
rect 2285 6905 2335 6955
rect 2585 6905 2635 6955
rect 2885 6905 2935 6955
rect 3185 6905 3235 6955
rect 4475 6905 4525 6955
rect 5315 6905 5365 6955
rect 5465 6905 5515 6955
rect 6275 6905 6325 6955
rect 7565 6905 7615 6955
rect 7865 6905 7915 6955
rect 8165 6905 8215 6955
rect 8465 6905 8515 6955
rect 8765 6905 8815 6955
rect 9065 6905 9115 6955
rect 9365 6905 9415 6955
rect 9995 6905 10045 6955
rect 10145 6905 10195 6955
rect 605 6755 655 6805
rect 755 6755 805 6805
rect 1385 6755 1435 6805
rect 1685 6755 1735 6805
rect 1985 6755 2035 6805
rect 2285 6755 2335 6805
rect 2585 6755 2635 6805
rect 2885 6755 2935 6805
rect 3185 6755 3235 6805
rect 4475 6755 4525 6805
rect 5315 6755 5365 6805
rect 5465 6755 5515 6805
rect 6275 6755 6325 6805
rect 7565 6755 7615 6805
rect 7865 6755 7915 6805
rect 8165 6755 8215 6805
rect 8465 6755 8515 6805
rect 8765 6755 8815 6805
rect 9065 6755 9115 6805
rect 9365 6755 9415 6805
rect 9995 6755 10045 6805
rect 10145 6755 10195 6805
rect 605 6605 655 6655
rect 755 6605 805 6655
rect 1385 6605 1435 6655
rect 1685 6605 1735 6655
rect 1985 6605 2035 6655
rect 2285 6605 2335 6655
rect 2585 6605 2635 6655
rect 2885 6605 2935 6655
rect 3185 6605 3235 6655
rect 4475 6605 4525 6655
rect 5315 6605 5365 6655
rect 5465 6605 5515 6655
rect 6275 6605 6325 6655
rect 7565 6605 7615 6655
rect 7865 6605 7915 6655
rect 8165 6605 8215 6655
rect 8465 6605 8515 6655
rect 8765 6605 8815 6655
rect 9065 6605 9115 6655
rect 9365 6605 9415 6655
rect 9995 6605 10045 6655
rect 10145 6605 10195 6655
rect 65 6155 115 6205
rect 215 6155 265 6205
rect 10535 6155 10585 6205
rect 10685 6155 10735 6205
rect 65 5915 115 5965
rect 215 5915 265 5965
rect 10535 5915 10585 5965
rect 10685 5915 10735 5965
rect 65 5675 115 5725
rect 215 5675 265 5725
rect 10535 5675 10585 5725
rect 10685 5675 10735 5725
rect 605 4955 655 5005
rect 755 4955 805 5005
rect 1385 4955 1435 5005
rect 1685 4955 1735 5005
rect 1985 4955 2035 5005
rect 2285 4955 2335 5005
rect 2585 4955 2635 5005
rect 2885 4955 2935 5005
rect 3185 4955 3235 5005
rect 4475 4955 4525 5005
rect 5315 4955 5365 5005
rect 5465 4955 5515 5005
rect 6275 4955 6325 5005
rect 7565 4955 7615 5005
rect 7865 4955 7915 5005
rect 8165 4955 8215 5005
rect 8465 4955 8515 5005
rect 8765 4955 8815 5005
rect 9065 4955 9115 5005
rect 9365 4955 9415 5005
rect 9995 4955 10045 5005
rect 10145 4955 10195 5005
rect 605 4805 655 4855
rect 755 4805 805 4855
rect 1385 4805 1435 4855
rect 1685 4805 1735 4855
rect 1985 4805 2035 4855
rect 2285 4805 2335 4855
rect 2585 4805 2635 4855
rect 2885 4805 2935 4855
rect 3185 4805 3235 4855
rect 4475 4805 4525 4855
rect 5315 4805 5365 4855
rect 5465 4805 5515 4855
rect 6275 4805 6325 4855
rect 7565 4805 7615 4855
rect 7865 4805 7915 4855
rect 8165 4805 8215 4855
rect 8465 4805 8515 4855
rect 8765 4805 8815 4855
rect 9065 4805 9115 4855
rect 9365 4805 9415 4855
rect 9995 4805 10045 4855
rect 10145 4805 10195 4855
rect 605 4655 655 4705
rect 755 4655 805 4705
rect 1385 4655 1435 4705
rect 1685 4655 1735 4705
rect 1985 4655 2035 4705
rect 2285 4655 2335 4705
rect 2585 4655 2635 4705
rect 2885 4655 2935 4705
rect 3185 4655 3235 4705
rect 4475 4655 4525 4705
rect 5315 4655 5365 4705
rect 5465 4655 5515 4705
rect 6275 4655 6325 4705
rect 7565 4655 7615 4705
rect 7865 4655 7915 4705
rect 8165 4655 8215 4705
rect 8465 4655 8515 4705
rect 8765 4655 8815 4705
rect 9065 4655 9115 4705
rect 9365 4655 9415 4705
rect 9995 4655 10045 4705
rect 10145 4655 10195 4705
rect 155 4115 205 4165
rect 395 4115 445 4165
rect 635 4115 685 4165
rect 1355 4115 1405 4165
rect 1595 4115 1645 4165
rect 1835 4115 1885 4165
rect 2075 4115 2125 4165
rect 2315 4115 2365 4165
rect 2555 4115 2605 4165
rect 2795 4115 2845 4165
rect 3035 4115 3085 4165
rect 3275 4115 3325 4165
rect 4475 4115 4525 4165
rect 5435 4115 5485 4165
rect 6275 4115 6325 4165
rect 7475 4115 7525 4165
rect 7715 4115 7765 4165
rect 7955 4115 8005 4165
rect 8195 4115 8245 4165
rect 8435 4115 8485 4165
rect 8675 4115 8725 4165
rect 8915 4115 8965 4165
rect 9155 4115 9205 4165
rect 9395 4115 9445 4165
rect 10115 4115 10165 4165
rect 10355 4115 10405 4165
rect 10595 4115 10645 4165
rect 155 3965 205 4015
rect 395 3965 445 4015
rect 635 3965 685 4015
rect 1355 3965 1405 4015
rect 1595 3965 1645 4015
rect 1835 3965 1885 4015
rect 2075 3965 2125 4015
rect 2315 3965 2365 4015
rect 2555 3965 2605 4015
rect 2795 3965 2845 4015
rect 3035 3965 3085 4015
rect 3275 3965 3325 4015
rect 4475 3965 4525 4015
rect 5435 3965 5485 4015
rect 6275 3965 6325 4015
rect 7475 3965 7525 4015
rect 7715 3965 7765 4015
rect 7955 3965 8005 4015
rect 8195 3965 8245 4015
rect 8435 3965 8485 4015
rect 8675 3965 8725 4015
rect 8915 3965 8965 4015
rect 9155 3965 9205 4015
rect 9395 3965 9445 4015
rect 10115 3965 10165 4015
rect 10355 3965 10405 4015
rect 10595 3965 10645 4015
rect 155 3605 205 3655
rect 395 3605 445 3655
rect 635 3605 685 3655
rect 1355 3605 1405 3655
rect 1595 3605 1645 3655
rect 1835 3605 1885 3655
rect 2075 3605 2125 3655
rect 2315 3605 2365 3655
rect 2555 3605 2605 3655
rect 2795 3605 2845 3655
rect 3035 3605 3085 3655
rect 3275 3605 3325 3655
rect 4475 3605 4525 3655
rect 5435 3605 5485 3655
rect 6275 3605 6325 3655
rect 7475 3605 7525 3655
rect 7715 3605 7765 3655
rect 7955 3605 8005 3655
rect 8195 3605 8245 3655
rect 8435 3605 8485 3655
rect 8675 3605 8725 3655
rect 8915 3605 8965 3655
rect 9155 3605 9205 3655
rect 9395 3605 9445 3655
rect 10115 3605 10165 3655
rect 10355 3605 10405 3655
rect 10595 3605 10645 3655
rect 155 3455 205 3505
rect 395 3455 445 3505
rect 635 3455 685 3505
rect 1355 3455 1405 3505
rect 1595 3455 1645 3505
rect 1835 3455 1885 3505
rect 2075 3455 2125 3505
rect 2315 3455 2365 3505
rect 2555 3455 2605 3505
rect 2795 3455 2845 3505
rect 3035 3455 3085 3505
rect 3275 3455 3325 3505
rect 4475 3455 4525 3505
rect 5435 3455 5485 3505
rect 6275 3455 6325 3505
rect 7475 3455 7525 3505
rect 7715 3455 7765 3505
rect 7955 3455 8005 3505
rect 8195 3455 8245 3505
rect 8435 3455 8485 3505
rect 8675 3455 8725 3505
rect 8915 3455 8965 3505
rect 9155 3455 9205 3505
rect 9395 3455 9445 3505
rect 10115 3455 10165 3505
rect 10355 3455 10405 3505
rect 10595 3455 10645 3505
rect 65 2225 115 2275
rect 215 2225 265 2275
rect 725 2225 775 2275
rect 875 2225 925 2275
rect 1025 2225 1075 2275
rect 1175 2225 1225 2275
rect 9575 2225 9625 2275
rect 9725 2225 9775 2275
rect 9875 2225 9925 2275
rect 10025 2225 10075 2275
rect 10535 2225 10585 2275
rect 10685 2225 10735 2275
rect 65 2075 115 2125
rect 215 2075 265 2125
rect 725 2075 775 2125
rect 875 2075 925 2125
rect 1025 2075 1075 2125
rect 1175 2075 1225 2125
rect 9575 2075 9625 2125
rect 9725 2075 9775 2125
rect 9875 2075 9925 2125
rect 10025 2075 10075 2125
rect 10535 2075 10585 2125
rect 10685 2075 10735 2125
rect 65 1925 115 1975
rect 215 1925 265 1975
rect 725 1925 775 1975
rect 875 1925 925 1975
rect 1025 1925 1075 1975
rect 1175 1925 1225 1975
rect 9575 1925 9625 1975
rect 9725 1925 9775 1975
rect 9875 1925 9925 1975
rect 10025 1925 10075 1975
rect 10535 1925 10585 1975
rect 10685 1925 10735 1975
rect 65 1775 115 1825
rect 215 1775 265 1825
rect 725 1775 775 1825
rect 875 1775 925 1825
rect 1025 1775 1075 1825
rect 1175 1775 1225 1825
rect 9575 1775 9625 1825
rect 9725 1775 9775 1825
rect 9875 1775 9925 1825
rect 10025 1775 10075 1825
rect 10535 1775 10585 1825
rect 10685 1775 10735 1825
rect 65 1625 115 1675
rect 215 1625 265 1675
rect 725 1625 775 1675
rect 875 1625 925 1675
rect 1025 1625 1075 1675
rect 1175 1625 1225 1675
rect 9575 1625 9625 1675
rect 9725 1625 9775 1675
rect 9875 1625 9925 1675
rect 10025 1625 10075 1675
rect 10535 1625 10585 1675
rect 10685 1625 10735 1675
rect 95 215 145 265
rect 875 215 925 265
rect 1115 215 1165 265
rect 1355 215 1405 265
rect 1595 215 1645 265
rect 1835 215 1885 265
rect 2075 215 2125 265
rect 2315 215 2365 265
rect 2555 215 2605 265
rect 2795 215 2845 265
rect 3035 215 3085 265
rect 3275 215 3325 265
rect 3515 215 3565 265
rect 3755 215 3805 265
rect 3995 215 4045 265
rect 4235 215 4285 265
rect 4475 215 4525 265
rect 4715 215 4765 265
rect 4955 215 5005 265
rect 5795 215 5845 265
rect 6035 215 6085 265
rect 6275 215 6325 265
rect 6515 215 6565 265
rect 6755 215 6805 265
rect 6995 215 7045 265
rect 7235 215 7285 265
rect 7475 215 7525 265
rect 7715 215 7765 265
rect 7955 215 8005 265
rect 8195 215 8245 265
rect 8435 215 8485 265
rect 8675 215 8725 265
rect 8915 215 8965 265
rect 9155 215 9205 265
rect 9395 215 9445 265
rect 9635 215 9685 265
rect 9875 215 9925 265
rect 10655 215 10705 265
rect 95 65 145 115
rect 875 65 925 115
rect 1115 65 1165 115
rect 1355 65 1405 115
rect 1595 65 1645 115
rect 1835 65 1885 115
rect 2075 65 2125 115
rect 2315 65 2365 115
rect 2555 65 2605 115
rect 2795 65 2845 115
rect 3035 65 3085 115
rect 3275 65 3325 115
rect 3515 65 3565 115
rect 3755 65 3805 115
rect 3995 65 4045 115
rect 4235 65 4285 115
rect 4475 65 4525 115
rect 4715 65 4765 115
rect 4955 65 5005 115
rect 5795 65 5845 115
rect 6035 65 6085 115
rect 6275 65 6325 115
rect 6515 65 6565 115
rect 6755 65 6805 115
rect 6995 65 7045 115
rect 7235 65 7285 115
rect 7475 65 7525 115
rect 7715 65 7765 115
rect 7955 65 8005 115
rect 8195 65 8245 115
rect 8435 65 8485 115
rect 8675 65 8725 115
rect 8915 65 8965 115
rect 9155 65 9205 115
rect 9395 65 9445 115
rect 9635 65 9685 115
rect 9875 65 9925 115
rect 10655 65 10705 115
<< metal3 >>
rect 1530 30810 9270 30930
rect 1530 23310 1650 30810
rect 9150 23310 9270 30810
rect 1530 23190 9270 23310
rect 690 0 1170 20850
rect 1650 0 2130 20850
rect 2610 0 3090 20850
rect 3570 0 4050 20850
rect 4530 0 5010 20850
rect 5790 0 6270 20850
rect 6750 0 7230 20850
rect 7710 0 8190 20850
rect 8670 0 9150 20850
rect 9630 0 10110 20850
<< via2 >>
rect 1925 30485 1975 30535
rect 2225 30485 2275 30535
rect 2525 30485 2575 30535
rect 2825 30485 2875 30535
rect 3125 30485 3175 30535
rect 3425 30485 3475 30535
rect 3725 30485 3775 30535
rect 4025 30485 4075 30535
rect 4325 30485 4375 30535
rect 4625 30485 4675 30535
rect 4925 30485 4975 30535
rect 5225 30485 5275 30535
rect 5525 30485 5575 30535
rect 5825 30485 5875 30535
rect 6125 30485 6175 30535
rect 6425 30485 6475 30535
rect 6725 30485 6775 30535
rect 7025 30485 7075 30535
rect 7325 30485 7375 30535
rect 7625 30485 7675 30535
rect 7925 30485 7975 30535
rect 8225 30485 8275 30535
rect 8525 30485 8575 30535
rect 8825 30485 8875 30535
rect 1925 30185 1975 30235
rect 2225 30185 2275 30235
rect 2525 30185 2575 30235
rect 2825 30185 2875 30235
rect 3125 30185 3175 30235
rect 3425 30185 3475 30235
rect 3725 30185 3775 30235
rect 4025 30185 4075 30235
rect 4325 30185 4375 30235
rect 4625 30185 4675 30235
rect 4925 30185 4975 30235
rect 5225 30185 5275 30235
rect 5525 30185 5575 30235
rect 5825 30185 5875 30235
rect 6125 30185 6175 30235
rect 6425 30185 6475 30235
rect 6725 30185 6775 30235
rect 7025 30185 7075 30235
rect 7325 30185 7375 30235
rect 7625 30185 7675 30235
rect 7925 30185 7975 30235
rect 8225 30185 8275 30235
rect 8525 30185 8575 30235
rect 8825 30185 8875 30235
rect 1925 29885 1975 29935
rect 2225 29885 2275 29935
rect 2525 29885 2575 29935
rect 2825 29885 2875 29935
rect 3125 29885 3175 29935
rect 3425 29885 3475 29935
rect 3725 29885 3775 29935
rect 4025 29885 4075 29935
rect 4325 29885 4375 29935
rect 4625 29885 4675 29935
rect 4925 29885 4975 29935
rect 5225 29885 5275 29935
rect 5525 29885 5575 29935
rect 5825 29885 5875 29935
rect 6125 29885 6175 29935
rect 6425 29885 6475 29935
rect 6725 29885 6775 29935
rect 7025 29885 7075 29935
rect 7325 29885 7375 29935
rect 7625 29885 7675 29935
rect 7925 29885 7975 29935
rect 8225 29885 8275 29935
rect 8525 29885 8575 29935
rect 8825 29885 8875 29935
rect 1925 29585 1975 29635
rect 2225 29585 2275 29635
rect 2525 29585 2575 29635
rect 2825 29585 2875 29635
rect 3125 29585 3175 29635
rect 3425 29585 3475 29635
rect 3725 29585 3775 29635
rect 4025 29585 4075 29635
rect 4325 29585 4375 29635
rect 4625 29585 4675 29635
rect 4925 29585 4975 29635
rect 5225 29585 5275 29635
rect 5525 29585 5575 29635
rect 5825 29585 5875 29635
rect 6125 29585 6175 29635
rect 6425 29585 6475 29635
rect 6725 29585 6775 29635
rect 7025 29585 7075 29635
rect 7325 29585 7375 29635
rect 7625 29585 7675 29635
rect 7925 29585 7975 29635
rect 8225 29585 8275 29635
rect 8525 29585 8575 29635
rect 8825 29585 8875 29635
rect 1925 29285 1975 29335
rect 2225 29285 2275 29335
rect 2525 29285 2575 29335
rect 2825 29285 2875 29335
rect 3125 29285 3175 29335
rect 3425 29285 3475 29335
rect 3725 29285 3775 29335
rect 4025 29285 4075 29335
rect 4325 29285 4375 29335
rect 4625 29285 4675 29335
rect 4925 29285 4975 29335
rect 5225 29285 5275 29335
rect 5525 29285 5575 29335
rect 5825 29285 5875 29335
rect 6125 29285 6175 29335
rect 6425 29285 6475 29335
rect 6725 29285 6775 29335
rect 7025 29285 7075 29335
rect 7325 29285 7375 29335
rect 7625 29285 7675 29335
rect 7925 29285 7975 29335
rect 8225 29285 8275 29335
rect 8525 29285 8575 29335
rect 8825 29285 8875 29335
rect 1925 28985 1975 29035
rect 2225 28985 2275 29035
rect 2525 28985 2575 29035
rect 2825 28985 2875 29035
rect 3125 28985 3175 29035
rect 3425 28985 3475 29035
rect 3725 28985 3775 29035
rect 4025 28985 4075 29035
rect 4325 28985 4375 29035
rect 4625 28985 4675 29035
rect 4925 28985 4975 29035
rect 5225 28985 5275 29035
rect 5525 28985 5575 29035
rect 5825 28985 5875 29035
rect 6125 28985 6175 29035
rect 6425 28985 6475 29035
rect 6725 28985 6775 29035
rect 7025 28985 7075 29035
rect 7325 28985 7375 29035
rect 7625 28985 7675 29035
rect 7925 28985 7975 29035
rect 8225 28985 8275 29035
rect 8525 28985 8575 29035
rect 8825 28985 8875 29035
rect 1925 28685 1975 28735
rect 2225 28685 2275 28735
rect 2525 28685 2575 28735
rect 2825 28685 2875 28735
rect 3125 28685 3175 28735
rect 3425 28685 3475 28735
rect 3725 28685 3775 28735
rect 4025 28685 4075 28735
rect 4325 28685 4375 28735
rect 4625 28685 4675 28735
rect 4925 28685 4975 28735
rect 5225 28685 5275 28735
rect 5525 28685 5575 28735
rect 5825 28685 5875 28735
rect 6125 28685 6175 28735
rect 6425 28685 6475 28735
rect 6725 28685 6775 28735
rect 7025 28685 7075 28735
rect 7325 28685 7375 28735
rect 7625 28685 7675 28735
rect 7925 28685 7975 28735
rect 8225 28685 8275 28735
rect 8525 28685 8575 28735
rect 8825 28685 8875 28735
rect 1925 28385 1975 28435
rect 2225 28385 2275 28435
rect 2525 28385 2575 28435
rect 2825 28385 2875 28435
rect 3125 28385 3175 28435
rect 3425 28385 3475 28435
rect 3725 28385 3775 28435
rect 4025 28385 4075 28435
rect 4325 28385 4375 28435
rect 4625 28385 4675 28435
rect 4925 28385 4975 28435
rect 5225 28385 5275 28435
rect 5525 28385 5575 28435
rect 5825 28385 5875 28435
rect 6125 28385 6175 28435
rect 6425 28385 6475 28435
rect 6725 28385 6775 28435
rect 7025 28385 7075 28435
rect 7325 28385 7375 28435
rect 7625 28385 7675 28435
rect 7925 28385 7975 28435
rect 8225 28385 8275 28435
rect 8525 28385 8575 28435
rect 8825 28385 8875 28435
rect 1925 28085 1975 28135
rect 2225 28085 2275 28135
rect 2525 28085 2575 28135
rect 2825 28085 2875 28135
rect 3125 28085 3175 28135
rect 3425 28085 3475 28135
rect 3725 28085 3775 28135
rect 4025 28085 4075 28135
rect 4325 28085 4375 28135
rect 4625 28085 4675 28135
rect 4925 28085 4975 28135
rect 5225 28085 5275 28135
rect 5525 28085 5575 28135
rect 5825 28085 5875 28135
rect 6125 28085 6175 28135
rect 6425 28085 6475 28135
rect 6725 28085 6775 28135
rect 7025 28085 7075 28135
rect 7325 28085 7375 28135
rect 7625 28085 7675 28135
rect 7925 28085 7975 28135
rect 8225 28085 8275 28135
rect 8525 28085 8575 28135
rect 8825 28085 8875 28135
rect 1925 27785 1975 27835
rect 2225 27785 2275 27835
rect 2525 27785 2575 27835
rect 2825 27785 2875 27835
rect 3125 27785 3175 27835
rect 3425 27785 3475 27835
rect 3725 27785 3775 27835
rect 4025 27785 4075 27835
rect 4325 27785 4375 27835
rect 4625 27785 4675 27835
rect 4925 27785 4975 27835
rect 5225 27785 5275 27835
rect 5525 27785 5575 27835
rect 5825 27785 5875 27835
rect 6125 27785 6175 27835
rect 6425 27785 6475 27835
rect 6725 27785 6775 27835
rect 7025 27785 7075 27835
rect 7325 27785 7375 27835
rect 7625 27785 7675 27835
rect 7925 27785 7975 27835
rect 8225 27785 8275 27835
rect 8525 27785 8575 27835
rect 8825 27785 8875 27835
rect 1925 27485 1975 27535
rect 2225 27485 2275 27535
rect 2525 27485 2575 27535
rect 2825 27485 2875 27535
rect 3125 27485 3175 27535
rect 3425 27485 3475 27535
rect 3725 27485 3775 27535
rect 4025 27485 4075 27535
rect 4325 27485 4375 27535
rect 4625 27485 4675 27535
rect 4925 27485 4975 27535
rect 5225 27485 5275 27535
rect 5525 27485 5575 27535
rect 5825 27485 5875 27535
rect 6125 27485 6175 27535
rect 6425 27485 6475 27535
rect 6725 27485 6775 27535
rect 7025 27485 7075 27535
rect 7325 27485 7375 27535
rect 7625 27485 7675 27535
rect 7925 27485 7975 27535
rect 8225 27485 8275 27535
rect 8525 27485 8575 27535
rect 8825 27485 8875 27535
rect 1925 27185 1975 27235
rect 2225 27185 2275 27235
rect 2525 27185 2575 27235
rect 2825 27185 2875 27235
rect 3125 27185 3175 27235
rect 3425 27185 3475 27235
rect 3725 27185 3775 27235
rect 4025 27185 4075 27235
rect 4325 27185 4375 27235
rect 4625 27185 4675 27235
rect 4925 27185 4975 27235
rect 5225 27185 5275 27235
rect 5525 27185 5575 27235
rect 5825 27185 5875 27235
rect 6125 27185 6175 27235
rect 6425 27185 6475 27235
rect 6725 27185 6775 27235
rect 7025 27185 7075 27235
rect 7325 27185 7375 27235
rect 7625 27185 7675 27235
rect 7925 27185 7975 27235
rect 8225 27185 8275 27235
rect 8525 27185 8575 27235
rect 8825 27185 8875 27235
rect 1925 26885 1975 26935
rect 2225 26885 2275 26935
rect 2525 26885 2575 26935
rect 2825 26885 2875 26935
rect 3125 26885 3175 26935
rect 3425 26885 3475 26935
rect 3725 26885 3775 26935
rect 4025 26885 4075 26935
rect 4325 26885 4375 26935
rect 4625 26885 4675 26935
rect 4925 26885 4975 26935
rect 5225 26885 5275 26935
rect 5525 26885 5575 26935
rect 5825 26885 5875 26935
rect 6125 26885 6175 26935
rect 6425 26885 6475 26935
rect 6725 26885 6775 26935
rect 7025 26885 7075 26935
rect 7325 26885 7375 26935
rect 7625 26885 7675 26935
rect 7925 26885 7975 26935
rect 8225 26885 8275 26935
rect 8525 26885 8575 26935
rect 8825 26885 8875 26935
rect 1925 26585 1975 26635
rect 2225 26585 2275 26635
rect 2525 26585 2575 26635
rect 2825 26585 2875 26635
rect 3125 26585 3175 26635
rect 3425 26585 3475 26635
rect 3725 26585 3775 26635
rect 4025 26585 4075 26635
rect 4325 26585 4375 26635
rect 4625 26585 4675 26635
rect 4925 26585 4975 26635
rect 5225 26585 5275 26635
rect 5525 26585 5575 26635
rect 5825 26585 5875 26635
rect 6125 26585 6175 26635
rect 6425 26585 6475 26635
rect 6725 26585 6775 26635
rect 7025 26585 7075 26635
rect 7325 26585 7375 26635
rect 7625 26585 7675 26635
rect 7925 26585 7975 26635
rect 8225 26585 8275 26635
rect 8525 26585 8575 26635
rect 8825 26585 8875 26635
rect 1925 26285 1975 26335
rect 2225 26285 2275 26335
rect 2525 26285 2575 26335
rect 2825 26285 2875 26335
rect 3125 26285 3175 26335
rect 3425 26285 3475 26335
rect 3725 26285 3775 26335
rect 4025 26285 4075 26335
rect 4325 26285 4375 26335
rect 4625 26285 4675 26335
rect 4925 26285 4975 26335
rect 5225 26285 5275 26335
rect 5525 26285 5575 26335
rect 5825 26285 5875 26335
rect 6125 26285 6175 26335
rect 6425 26285 6475 26335
rect 6725 26285 6775 26335
rect 7025 26285 7075 26335
rect 7325 26285 7375 26335
rect 7625 26285 7675 26335
rect 7925 26285 7975 26335
rect 8225 26285 8275 26335
rect 8525 26285 8575 26335
rect 8825 26285 8875 26335
rect 1925 25985 1975 26035
rect 2225 25985 2275 26035
rect 2525 25985 2575 26035
rect 2825 25985 2875 26035
rect 3125 25985 3175 26035
rect 3425 25985 3475 26035
rect 3725 25985 3775 26035
rect 4025 25985 4075 26035
rect 4325 25985 4375 26035
rect 4625 25985 4675 26035
rect 4925 25985 4975 26035
rect 5225 25985 5275 26035
rect 5525 25985 5575 26035
rect 5825 25985 5875 26035
rect 6125 25985 6175 26035
rect 6425 25985 6475 26035
rect 6725 25985 6775 26035
rect 7025 25985 7075 26035
rect 7325 25985 7375 26035
rect 7625 25985 7675 26035
rect 7925 25985 7975 26035
rect 8225 25985 8275 26035
rect 8525 25985 8575 26035
rect 8825 25985 8875 26035
rect 1925 25685 1975 25735
rect 2225 25685 2275 25735
rect 2525 25685 2575 25735
rect 2825 25685 2875 25735
rect 3125 25685 3175 25735
rect 3425 25685 3475 25735
rect 3725 25685 3775 25735
rect 4025 25685 4075 25735
rect 4325 25685 4375 25735
rect 4625 25685 4675 25735
rect 4925 25685 4975 25735
rect 5225 25685 5275 25735
rect 5525 25685 5575 25735
rect 5825 25685 5875 25735
rect 6125 25685 6175 25735
rect 6425 25685 6475 25735
rect 6725 25685 6775 25735
rect 7025 25685 7075 25735
rect 7325 25685 7375 25735
rect 7625 25685 7675 25735
rect 7925 25685 7975 25735
rect 8225 25685 8275 25735
rect 8525 25685 8575 25735
rect 8825 25685 8875 25735
rect 1925 25385 1975 25435
rect 2225 25385 2275 25435
rect 2525 25385 2575 25435
rect 2825 25385 2875 25435
rect 3125 25385 3175 25435
rect 3425 25385 3475 25435
rect 3725 25385 3775 25435
rect 4025 25385 4075 25435
rect 4325 25385 4375 25435
rect 4625 25385 4675 25435
rect 4925 25385 4975 25435
rect 5225 25385 5275 25435
rect 5525 25385 5575 25435
rect 5825 25385 5875 25435
rect 6125 25385 6175 25435
rect 6425 25385 6475 25435
rect 6725 25385 6775 25435
rect 7025 25385 7075 25435
rect 7325 25385 7375 25435
rect 7625 25385 7675 25435
rect 7925 25385 7975 25435
rect 8225 25385 8275 25435
rect 8525 25385 8575 25435
rect 8825 25385 8875 25435
rect 1925 25085 1975 25135
rect 2225 25085 2275 25135
rect 2525 25085 2575 25135
rect 2825 25085 2875 25135
rect 3125 25085 3175 25135
rect 3425 25085 3475 25135
rect 3725 25085 3775 25135
rect 4025 25085 4075 25135
rect 4325 25085 4375 25135
rect 4625 25085 4675 25135
rect 4925 25085 4975 25135
rect 5225 25085 5275 25135
rect 5525 25085 5575 25135
rect 5825 25085 5875 25135
rect 6125 25085 6175 25135
rect 6425 25085 6475 25135
rect 6725 25085 6775 25135
rect 7025 25085 7075 25135
rect 7325 25085 7375 25135
rect 7625 25085 7675 25135
rect 7925 25085 7975 25135
rect 8225 25085 8275 25135
rect 8525 25085 8575 25135
rect 8825 25085 8875 25135
rect 1925 24785 1975 24835
rect 2225 24785 2275 24835
rect 2525 24785 2575 24835
rect 2825 24785 2875 24835
rect 3125 24785 3175 24835
rect 3425 24785 3475 24835
rect 3725 24785 3775 24835
rect 4025 24785 4075 24835
rect 4325 24785 4375 24835
rect 4625 24785 4675 24835
rect 4925 24785 4975 24835
rect 5225 24785 5275 24835
rect 5525 24785 5575 24835
rect 5825 24785 5875 24835
rect 6125 24785 6175 24835
rect 6425 24785 6475 24835
rect 6725 24785 6775 24835
rect 7025 24785 7075 24835
rect 7325 24785 7375 24835
rect 7625 24785 7675 24835
rect 7925 24785 7975 24835
rect 8225 24785 8275 24835
rect 8525 24785 8575 24835
rect 8825 24785 8875 24835
rect 1925 24485 1975 24535
rect 2225 24485 2275 24535
rect 2525 24485 2575 24535
rect 2825 24485 2875 24535
rect 3125 24485 3175 24535
rect 3425 24485 3475 24535
rect 3725 24485 3775 24535
rect 4025 24485 4075 24535
rect 4325 24485 4375 24535
rect 4625 24485 4675 24535
rect 4925 24485 4975 24535
rect 5225 24485 5275 24535
rect 5525 24485 5575 24535
rect 5825 24485 5875 24535
rect 6125 24485 6175 24535
rect 6425 24485 6475 24535
rect 6725 24485 6775 24535
rect 7025 24485 7075 24535
rect 7325 24485 7375 24535
rect 7625 24485 7675 24535
rect 7925 24485 7975 24535
rect 8225 24485 8275 24535
rect 8525 24485 8575 24535
rect 8825 24485 8875 24535
rect 1925 24185 1975 24235
rect 2225 24185 2275 24235
rect 2525 24185 2575 24235
rect 2825 24185 2875 24235
rect 3125 24185 3175 24235
rect 3425 24185 3475 24235
rect 3725 24185 3775 24235
rect 4025 24185 4075 24235
rect 4325 24185 4375 24235
rect 4625 24185 4675 24235
rect 4925 24185 4975 24235
rect 5225 24185 5275 24235
rect 5525 24185 5575 24235
rect 5825 24185 5875 24235
rect 6125 24185 6175 24235
rect 6425 24185 6475 24235
rect 6725 24185 6775 24235
rect 7025 24185 7075 24235
rect 7325 24185 7375 24235
rect 7625 24185 7675 24235
rect 7925 24185 7975 24235
rect 8225 24185 8275 24235
rect 8525 24185 8575 24235
rect 8825 24185 8875 24235
rect 1925 23885 1975 23935
rect 2225 23885 2275 23935
rect 2525 23885 2575 23935
rect 2825 23885 2875 23935
rect 3125 23885 3175 23935
rect 3425 23885 3475 23935
rect 3725 23885 3775 23935
rect 4025 23885 4075 23935
rect 4325 23885 4375 23935
rect 4625 23885 4675 23935
rect 4925 23885 4975 23935
rect 5225 23885 5275 23935
rect 5525 23885 5575 23935
rect 5825 23885 5875 23935
rect 6125 23885 6175 23935
rect 6425 23885 6475 23935
rect 6725 23885 6775 23935
rect 7025 23885 7075 23935
rect 7325 23885 7375 23935
rect 7625 23885 7675 23935
rect 7925 23885 7975 23935
rect 8225 23885 8275 23935
rect 8525 23885 8575 23935
rect 8825 23885 8875 23935
rect 1925 23585 1975 23635
rect 2225 23585 2275 23635
rect 2525 23585 2575 23635
rect 2825 23585 2875 23635
rect 3125 23585 3175 23635
rect 3425 23585 3475 23635
rect 3725 23585 3775 23635
rect 4025 23585 4075 23635
rect 4325 23585 4375 23635
rect 4625 23585 4675 23635
rect 4925 23585 4975 23635
rect 5225 23585 5275 23635
rect 5525 23585 5575 23635
rect 5825 23585 5875 23635
rect 6125 23585 6175 23635
rect 6425 23585 6475 23635
rect 6725 23585 6775 23635
rect 7025 23585 7075 23635
rect 7325 23585 7375 23635
rect 7625 23585 7675 23635
rect 7925 23585 7975 23635
rect 8225 23585 8275 23635
rect 8525 23585 8575 23635
rect 8825 23585 8875 23635
rect 755 20735 805 20785
rect 905 20735 955 20785
rect 1055 20735 1105 20785
rect 2675 20735 2725 20785
rect 2825 20735 2875 20785
rect 2975 20735 3025 20785
rect 4595 20735 4645 20785
rect 4745 20735 4795 20785
rect 4895 20735 4945 20785
rect 6815 20735 6865 20785
rect 6965 20735 7015 20785
rect 7115 20735 7165 20785
rect 8735 20735 8785 20785
rect 8885 20735 8935 20785
rect 9035 20735 9085 20785
rect 755 20585 805 20635
rect 905 20585 955 20635
rect 1055 20585 1105 20635
rect 2675 20585 2725 20635
rect 2825 20585 2875 20635
rect 2975 20585 3025 20635
rect 4595 20585 4645 20635
rect 4745 20585 4795 20635
rect 4895 20585 4945 20635
rect 6815 20585 6865 20635
rect 6965 20585 7015 20635
rect 7115 20585 7165 20635
rect 8735 20585 8785 20635
rect 8885 20585 8935 20635
rect 9035 20585 9085 20635
rect 1715 20045 1765 20095
rect 1865 20045 1915 20095
rect 2015 20045 2065 20095
rect 3635 20045 3685 20095
rect 3785 20045 3835 20095
rect 3935 20045 3985 20095
rect 5855 20045 5905 20095
rect 6005 20045 6055 20095
rect 6155 20045 6205 20095
rect 7775 20045 7825 20095
rect 7925 20045 7975 20095
rect 8075 20045 8125 20095
rect 9695 20045 9745 20095
rect 9845 20045 9895 20095
rect 9995 20045 10045 20095
rect 1715 19895 1765 19945
rect 1865 19895 1915 19945
rect 2015 19895 2065 19945
rect 3635 19895 3685 19945
rect 3785 19895 3835 19945
rect 3935 19895 3985 19945
rect 5855 19895 5905 19945
rect 6005 19895 6055 19945
rect 6155 19895 6205 19945
rect 7775 19895 7825 19945
rect 7925 19895 7975 19945
rect 8075 19895 8125 19945
rect 9695 19895 9745 19945
rect 9845 19895 9895 19945
rect 9995 19895 10045 19945
rect 1715 19745 1765 19795
rect 1865 19745 1915 19795
rect 2015 19745 2065 19795
rect 3635 19745 3685 19795
rect 3785 19745 3835 19795
rect 3935 19745 3985 19795
rect 5855 19745 5905 19795
rect 6005 19745 6055 19795
rect 6155 19745 6205 19795
rect 7775 19745 7825 19795
rect 7925 19745 7975 19795
rect 8075 19745 8125 19795
rect 9695 19745 9745 19795
rect 9845 19745 9895 19795
rect 9995 19745 10045 19795
rect 755 19205 805 19255
rect 905 19205 955 19255
rect 1055 19205 1105 19255
rect 2675 19205 2725 19255
rect 2825 19205 2875 19255
rect 2975 19205 3025 19255
rect 4595 19205 4645 19255
rect 4745 19205 4795 19255
rect 4895 19205 4945 19255
rect 6815 19205 6865 19255
rect 6965 19205 7015 19255
rect 7115 19205 7165 19255
rect 8735 19205 8785 19255
rect 8885 19205 8935 19255
rect 9035 19205 9085 19255
rect 755 19055 805 19105
rect 905 19055 955 19105
rect 1055 19055 1105 19105
rect 2675 19055 2725 19105
rect 2825 19055 2875 19105
rect 2975 19055 3025 19105
rect 4595 19055 4645 19105
rect 4745 19055 4795 19105
rect 4895 19055 4945 19105
rect 6815 19055 6865 19105
rect 6965 19055 7015 19105
rect 7115 19055 7165 19105
rect 8735 19055 8785 19105
rect 8885 19055 8935 19105
rect 9035 19055 9085 19105
rect 755 18905 805 18955
rect 905 18905 955 18955
rect 1055 18905 1105 18955
rect 2675 18905 2725 18955
rect 2825 18905 2875 18955
rect 2975 18905 3025 18955
rect 4595 18905 4645 18955
rect 4745 18905 4795 18955
rect 4895 18905 4945 18955
rect 6815 18905 6865 18955
rect 6965 18905 7015 18955
rect 7115 18905 7165 18955
rect 8735 18905 8785 18955
rect 8885 18905 8935 18955
rect 9035 18905 9085 18955
rect 755 18755 805 18805
rect 905 18755 955 18805
rect 1055 18755 1105 18805
rect 2675 18755 2725 18805
rect 2825 18755 2875 18805
rect 2975 18755 3025 18805
rect 4595 18755 4645 18805
rect 4745 18755 4795 18805
rect 4895 18755 4945 18805
rect 6815 18755 6865 18805
rect 6965 18755 7015 18805
rect 7115 18755 7165 18805
rect 8735 18755 8785 18805
rect 8885 18755 8935 18805
rect 9035 18755 9085 18805
rect 755 18605 805 18655
rect 905 18605 955 18655
rect 1055 18605 1105 18655
rect 2675 18605 2725 18655
rect 2825 18605 2875 18655
rect 2975 18605 3025 18655
rect 4595 18605 4645 18655
rect 4745 18605 4795 18655
rect 4895 18605 4945 18655
rect 6815 18605 6865 18655
rect 6965 18605 7015 18655
rect 7115 18605 7165 18655
rect 8735 18605 8785 18655
rect 8885 18605 8935 18655
rect 9035 18605 9085 18655
rect 1715 18095 1765 18145
rect 1865 18095 1915 18145
rect 2015 18095 2065 18145
rect 3635 18095 3685 18145
rect 3785 18095 3835 18145
rect 3935 18095 3985 18145
rect 5855 18095 5905 18145
rect 6005 18095 6055 18145
rect 6155 18095 6205 18145
rect 7775 18095 7825 18145
rect 7925 18095 7975 18145
rect 8075 18095 8125 18145
rect 9695 18095 9745 18145
rect 9845 18095 9895 18145
rect 9995 18095 10045 18145
rect 1715 17945 1765 17995
rect 1865 17945 1915 17995
rect 2015 17945 2065 17995
rect 3635 17945 3685 17995
rect 3785 17945 3835 17995
rect 3935 17945 3985 17995
rect 5855 17945 5905 17995
rect 6005 17945 6055 17995
rect 6155 17945 6205 17995
rect 7775 17945 7825 17995
rect 7925 17945 7975 17995
rect 8075 17945 8125 17995
rect 9695 17945 9745 17995
rect 9845 17945 9895 17995
rect 9995 17945 10045 17995
rect 1715 17795 1765 17845
rect 1865 17795 1915 17845
rect 2015 17795 2065 17845
rect 3635 17795 3685 17845
rect 3785 17795 3835 17845
rect 3935 17795 3985 17845
rect 5855 17795 5905 17845
rect 6005 17795 6055 17845
rect 6155 17795 6205 17845
rect 7775 17795 7825 17845
rect 7925 17795 7975 17845
rect 8075 17795 8125 17845
rect 9695 17795 9745 17845
rect 9845 17795 9895 17845
rect 9995 17795 10045 17845
rect 755 17405 805 17455
rect 905 17405 955 17455
rect 1055 17405 1105 17455
rect 2675 17405 2725 17455
rect 2825 17405 2875 17455
rect 2975 17405 3025 17455
rect 4595 17405 4645 17455
rect 4745 17405 4795 17455
rect 4895 17405 4945 17455
rect 6815 17405 6865 17455
rect 6965 17405 7015 17455
rect 7115 17405 7165 17455
rect 8735 17405 8785 17455
rect 8885 17405 8935 17455
rect 9035 17405 9085 17455
rect 755 17255 805 17305
rect 905 17255 955 17305
rect 1055 17255 1105 17305
rect 2675 17255 2725 17305
rect 2825 17255 2875 17305
rect 2975 17255 3025 17305
rect 4595 17255 4645 17305
rect 4745 17255 4795 17305
rect 4895 17255 4945 17305
rect 6815 17255 6865 17305
rect 6965 17255 7015 17305
rect 7115 17255 7165 17305
rect 8735 17255 8785 17305
rect 8885 17255 8935 17305
rect 9035 17255 9085 17305
rect 755 17105 805 17155
rect 905 17105 955 17155
rect 1055 17105 1105 17155
rect 2675 17105 2725 17155
rect 2825 17105 2875 17155
rect 2975 17105 3025 17155
rect 4595 17105 4645 17155
rect 4745 17105 4795 17155
rect 4895 17105 4945 17155
rect 6815 17105 6865 17155
rect 6965 17105 7015 17155
rect 7115 17105 7165 17155
rect 8735 17105 8785 17155
rect 8885 17105 8935 17155
rect 9035 17105 9085 17155
rect 755 16955 805 17005
rect 905 16955 955 17005
rect 1055 16955 1105 17005
rect 2675 16955 2725 17005
rect 2825 16955 2875 17005
rect 2975 16955 3025 17005
rect 4595 16955 4645 17005
rect 4745 16955 4795 17005
rect 4895 16955 4945 17005
rect 6815 16955 6865 17005
rect 6965 16955 7015 17005
rect 7115 16955 7165 17005
rect 8735 16955 8785 17005
rect 8885 16955 8935 17005
rect 9035 16955 9085 17005
rect 755 16805 805 16855
rect 905 16805 955 16855
rect 1055 16805 1105 16855
rect 2675 16805 2725 16855
rect 2825 16805 2875 16855
rect 2975 16805 3025 16855
rect 4595 16805 4645 16855
rect 4745 16805 4795 16855
rect 4895 16805 4945 16855
rect 6815 16805 6865 16855
rect 6965 16805 7015 16855
rect 7115 16805 7165 16855
rect 8735 16805 8785 16855
rect 8885 16805 8935 16855
rect 9035 16805 9085 16855
rect 1715 16145 1765 16195
rect 1865 16145 1915 16195
rect 2015 16145 2065 16195
rect 3635 16145 3685 16195
rect 3785 16145 3835 16195
rect 3935 16145 3985 16195
rect 5855 16115 5905 16165
rect 6005 16115 6055 16165
rect 6155 16115 6205 16165
rect 7775 16145 7825 16195
rect 7925 16145 7975 16195
rect 8075 16145 8125 16195
rect 9695 16145 9745 16195
rect 9845 16145 9895 16195
rect 9995 16145 10045 16195
rect 1715 15995 1765 16045
rect 1865 15995 1915 16045
rect 2015 15995 2065 16045
rect 3635 15995 3685 16045
rect 3785 15995 3835 16045
rect 3935 15995 3985 16045
rect 5855 15965 5905 16015
rect 6005 15965 6055 16015
rect 6155 15965 6205 16015
rect 7775 15995 7825 16045
rect 7925 15995 7975 16045
rect 8075 15995 8125 16045
rect 9695 15995 9745 16045
rect 9845 15995 9895 16045
rect 9995 15995 10045 16045
rect 1715 15845 1765 15895
rect 1865 15845 1915 15895
rect 2015 15845 2065 15895
rect 3635 15845 3685 15895
rect 3785 15845 3835 15895
rect 3935 15845 3985 15895
rect 5855 15815 5905 15865
rect 6005 15815 6055 15865
rect 6155 15815 6205 15865
rect 7775 15845 7825 15895
rect 7925 15845 7975 15895
rect 8075 15845 8125 15895
rect 9695 15845 9745 15895
rect 9845 15845 9895 15895
rect 9995 15845 10045 15895
rect 755 15455 805 15505
rect 905 15455 955 15505
rect 1055 15455 1105 15505
rect 2675 15455 2725 15505
rect 2825 15455 2875 15505
rect 2975 15455 3025 15505
rect 4595 15455 4645 15505
rect 4745 15455 4795 15505
rect 4895 15455 4945 15505
rect 6815 15455 6865 15505
rect 6965 15455 7015 15505
rect 7115 15455 7165 15505
rect 8735 15455 8785 15505
rect 8885 15455 8935 15505
rect 9035 15455 9085 15505
rect 755 15305 805 15355
rect 905 15305 955 15355
rect 1055 15305 1105 15355
rect 2675 15305 2725 15355
rect 2825 15305 2875 15355
rect 2975 15305 3025 15355
rect 4595 15305 4645 15355
rect 4745 15305 4795 15355
rect 4895 15305 4945 15355
rect 6815 15305 6865 15355
rect 6965 15305 7015 15355
rect 7115 15305 7165 15355
rect 8735 15305 8785 15355
rect 8885 15305 8935 15355
rect 9035 15305 9085 15355
rect 755 15155 805 15205
rect 905 15155 955 15205
rect 1055 15155 1105 15205
rect 2675 15155 2725 15205
rect 2825 15155 2875 15205
rect 2975 15155 3025 15205
rect 4595 15155 4645 15205
rect 4745 15155 4795 15205
rect 4895 15155 4945 15205
rect 6815 15155 6865 15205
rect 6965 15155 7015 15205
rect 7115 15155 7165 15205
rect 8735 15155 8785 15205
rect 8885 15155 8935 15205
rect 9035 15155 9085 15205
rect 755 15005 805 15055
rect 905 15005 955 15055
rect 1055 15005 1105 15055
rect 2675 15005 2725 15055
rect 2825 15005 2875 15055
rect 2975 15005 3025 15055
rect 4595 15005 4645 15055
rect 4745 15005 4795 15055
rect 4895 15005 4945 15055
rect 6815 15005 6865 15055
rect 6965 15005 7015 15055
rect 7115 15005 7165 15055
rect 8735 15005 8785 15055
rect 8885 15005 8935 15055
rect 9035 15005 9085 15055
rect 755 14855 805 14905
rect 905 14855 955 14905
rect 1055 14855 1105 14905
rect 2675 14855 2725 14905
rect 2825 14855 2875 14905
rect 2975 14855 3025 14905
rect 4595 14855 4645 14905
rect 4745 14855 4795 14905
rect 4895 14855 4945 14905
rect 6815 14855 6865 14905
rect 6965 14855 7015 14905
rect 7115 14855 7165 14905
rect 8735 14855 8785 14905
rect 8885 14855 8935 14905
rect 9035 14855 9085 14905
rect 1715 14195 1765 14245
rect 1865 14195 1915 14245
rect 2015 14195 2065 14245
rect 3635 14195 3685 14245
rect 3785 14195 3835 14245
rect 3935 14195 3985 14245
rect 5855 14165 5905 14215
rect 6005 14165 6055 14215
rect 6155 14165 6205 14215
rect 7775 14195 7825 14245
rect 7925 14195 7975 14245
rect 8075 14195 8125 14245
rect 9695 14195 9745 14245
rect 9845 14195 9895 14245
rect 9995 14195 10045 14245
rect 1715 14045 1765 14095
rect 1865 14045 1915 14095
rect 2015 14045 2065 14095
rect 3635 14045 3685 14095
rect 3785 14045 3835 14095
rect 3935 14045 3985 14095
rect 5855 14015 5905 14065
rect 6005 14015 6055 14065
rect 6155 14015 6205 14065
rect 7775 14045 7825 14095
rect 7925 14045 7975 14095
rect 8075 14045 8125 14095
rect 9695 14045 9745 14095
rect 9845 14045 9895 14095
rect 9995 14045 10045 14095
rect 1715 13895 1765 13945
rect 1865 13895 1915 13945
rect 2015 13895 2065 13945
rect 3635 13895 3685 13945
rect 3785 13895 3835 13945
rect 3935 13895 3985 13945
rect 5855 13865 5905 13915
rect 6005 13865 6055 13915
rect 6155 13865 6205 13915
rect 7775 13895 7825 13945
rect 7925 13895 7975 13945
rect 8075 13895 8125 13945
rect 9695 13895 9745 13945
rect 9845 13895 9895 13945
rect 9995 13895 10045 13945
rect 755 13355 805 13405
rect 905 13355 955 13405
rect 1055 13355 1105 13405
rect 2675 13355 2725 13405
rect 2825 13355 2875 13405
rect 2975 13355 3025 13405
rect 4595 13355 4645 13405
rect 4745 13355 4795 13405
rect 4895 13355 4945 13405
rect 6815 13355 6865 13405
rect 6965 13355 7015 13405
rect 7115 13355 7165 13405
rect 8735 13355 8785 13405
rect 8885 13355 8935 13405
rect 9035 13355 9085 13405
rect 755 13205 805 13255
rect 905 13205 955 13255
rect 1055 13205 1105 13255
rect 2675 13205 2725 13255
rect 2825 13205 2875 13255
rect 2975 13205 3025 13255
rect 4595 13205 4645 13255
rect 4745 13205 4795 13255
rect 4895 13205 4945 13255
rect 6815 13205 6865 13255
rect 6965 13205 7015 13255
rect 7115 13205 7165 13255
rect 8735 13205 8785 13255
rect 8885 13205 8935 13255
rect 9035 13205 9085 13255
rect 1715 12845 1765 12895
rect 1865 12845 1915 12895
rect 2015 12845 2065 12895
rect 3635 12845 3685 12895
rect 3785 12845 3835 12895
rect 3935 12845 3985 12895
rect 5855 12845 5905 12895
rect 6005 12845 6055 12895
rect 6155 12845 6205 12895
rect 7775 12845 7825 12895
rect 7925 12845 7975 12895
rect 8075 12845 8125 12895
rect 9695 12845 9745 12895
rect 9845 12845 9895 12895
rect 9995 12845 10045 12895
rect 1715 12695 1765 12745
rect 1865 12695 1915 12745
rect 2015 12695 2065 12745
rect 3635 12695 3685 12745
rect 3785 12695 3835 12745
rect 3935 12695 3985 12745
rect 5855 12695 5905 12745
rect 6005 12695 6055 12745
rect 6155 12695 6205 12745
rect 7775 12695 7825 12745
rect 7925 12695 7975 12745
rect 8075 12695 8125 12745
rect 9695 12695 9745 12745
rect 9845 12695 9895 12745
rect 9995 12695 10045 12745
rect 755 12005 805 12055
rect 905 12005 955 12055
rect 1055 12005 1105 12055
rect 2675 12005 2725 12055
rect 2825 12005 2875 12055
rect 2975 12005 3025 12055
rect 4595 12005 4645 12055
rect 4745 12005 4795 12055
rect 4895 12005 4945 12055
rect 6815 12005 6865 12055
rect 6965 12005 7015 12055
rect 7115 12005 7165 12055
rect 8735 12005 8785 12055
rect 8885 12005 8935 12055
rect 9035 12005 9085 12055
rect 755 11855 805 11905
rect 905 11855 955 11905
rect 1055 11855 1105 11905
rect 2675 11855 2725 11905
rect 2825 11855 2875 11905
rect 2975 11855 3025 11905
rect 4595 11855 4645 11905
rect 4745 11855 4795 11905
rect 4895 11855 4945 11905
rect 6815 11855 6865 11905
rect 6965 11855 7015 11905
rect 7115 11855 7165 11905
rect 8735 11855 8785 11905
rect 8885 11855 8935 11905
rect 9035 11855 9085 11905
rect 1715 11495 1765 11545
rect 1865 11495 1915 11545
rect 2015 11495 2065 11545
rect 3635 11495 3685 11545
rect 3785 11495 3835 11545
rect 3935 11495 3985 11545
rect 5855 11495 5905 11545
rect 6005 11495 6055 11545
rect 6155 11495 6205 11545
rect 7775 11495 7825 11545
rect 7925 11495 7975 11545
rect 8075 11495 8125 11545
rect 9695 11495 9745 11545
rect 9845 11495 9895 11545
rect 9995 11495 10045 11545
rect 1715 11345 1765 11395
rect 1865 11345 1915 11395
rect 2015 11345 2065 11395
rect 3635 11345 3685 11395
rect 3785 11345 3835 11395
rect 3935 11345 3985 11395
rect 5855 11345 5905 11395
rect 6005 11345 6055 11395
rect 6155 11345 6205 11395
rect 7775 11345 7825 11395
rect 7925 11345 7975 11395
rect 8075 11345 8125 11395
rect 9695 11345 9745 11395
rect 9845 11345 9895 11395
rect 9995 11345 10045 11395
rect 755 10805 805 10855
rect 905 10805 955 10855
rect 1055 10805 1105 10855
rect 2675 10805 2725 10855
rect 2825 10805 2875 10855
rect 2975 10805 3025 10855
rect 4595 10805 4645 10855
rect 4745 10805 4795 10855
rect 4895 10805 4945 10855
rect 6815 10805 6865 10855
rect 6965 10805 7015 10855
rect 7115 10805 7165 10855
rect 8735 10805 8785 10855
rect 8885 10805 8935 10855
rect 9035 10805 9085 10855
rect 755 10655 805 10705
rect 905 10655 955 10705
rect 1055 10655 1105 10705
rect 2675 10655 2725 10705
rect 2825 10655 2875 10705
rect 2975 10655 3025 10705
rect 4595 10655 4645 10705
rect 4745 10655 4795 10705
rect 4895 10655 4945 10705
rect 6815 10655 6865 10705
rect 6965 10655 7015 10705
rect 7115 10655 7165 10705
rect 8735 10655 8785 10705
rect 8885 10655 8935 10705
rect 9035 10655 9085 10705
rect 755 10505 805 10555
rect 905 10505 955 10555
rect 1055 10505 1105 10555
rect 2675 10505 2725 10555
rect 2825 10505 2875 10555
rect 2975 10505 3025 10555
rect 4595 10505 4645 10555
rect 4745 10505 4795 10555
rect 4895 10505 4945 10555
rect 6815 10505 6865 10555
rect 6965 10505 7015 10555
rect 7115 10505 7165 10555
rect 8735 10505 8785 10555
rect 8885 10505 8935 10555
rect 9035 10505 9085 10555
rect 1715 9965 1765 10015
rect 1865 9965 1915 10015
rect 2015 9965 2065 10015
rect 3635 9965 3685 10015
rect 3785 9965 3835 10015
rect 3935 9965 3985 10015
rect 5855 9965 5905 10015
rect 6005 9965 6055 10015
rect 6155 9965 6205 10015
rect 7775 9965 7825 10015
rect 7925 9965 7975 10015
rect 8075 9965 8125 10015
rect 9695 9965 9745 10015
rect 9845 9965 9895 10015
rect 9995 9965 10045 10015
rect 1715 9815 1765 9865
rect 1865 9815 1915 9865
rect 2015 9815 2065 9865
rect 3635 9815 3685 9865
rect 3785 9815 3835 9865
rect 3935 9815 3985 9865
rect 5855 9815 5905 9865
rect 6005 9815 6055 9865
rect 6155 9815 6205 9865
rect 7775 9815 7825 9865
rect 7925 9815 7975 9865
rect 8075 9815 8125 9865
rect 9695 9815 9745 9865
rect 9845 9815 9895 9865
rect 9995 9815 10045 9865
rect 1715 9665 1765 9715
rect 1865 9665 1915 9715
rect 2015 9665 2065 9715
rect 3635 9665 3685 9715
rect 3785 9665 3835 9715
rect 3935 9665 3985 9715
rect 5855 9665 5905 9715
rect 6005 9665 6055 9715
rect 6155 9665 6205 9715
rect 7775 9665 7825 9715
rect 7925 9665 7975 9715
rect 8075 9665 8125 9715
rect 9695 9665 9745 9715
rect 9845 9665 9895 9715
rect 9995 9665 10045 9715
rect 1715 9515 1765 9565
rect 1865 9515 1915 9565
rect 2015 9515 2065 9565
rect 3635 9515 3685 9565
rect 3785 9515 3835 9565
rect 3935 9515 3985 9565
rect 5855 9515 5905 9565
rect 6005 9515 6055 9565
rect 6155 9515 6205 9565
rect 7775 9515 7825 9565
rect 7925 9515 7975 9565
rect 8075 9515 8125 9565
rect 9695 9515 9745 9565
rect 9845 9515 9895 9565
rect 9995 9515 10045 9565
rect 1715 9365 1765 9415
rect 1865 9365 1915 9415
rect 2015 9365 2065 9415
rect 3635 9365 3685 9415
rect 3785 9365 3835 9415
rect 3935 9365 3985 9415
rect 5855 9365 5905 9415
rect 6005 9365 6055 9415
rect 6155 9365 6205 9415
rect 7775 9365 7825 9415
rect 7925 9365 7975 9415
rect 8075 9365 8125 9415
rect 9695 9365 9745 9415
rect 9845 9365 9895 9415
rect 9995 9365 10045 9415
rect 755 8855 805 8905
rect 905 8855 955 8905
rect 1055 8855 1105 8905
rect 2675 8855 2725 8905
rect 2825 8855 2875 8905
rect 2975 8855 3025 8905
rect 4595 8855 4645 8905
rect 4745 8855 4795 8905
rect 4895 8855 4945 8905
rect 6815 8855 6865 8905
rect 6965 8855 7015 8905
rect 7115 8855 7165 8905
rect 8735 8855 8785 8905
rect 8885 8855 8935 8905
rect 9035 8855 9085 8905
rect 755 8705 805 8755
rect 905 8705 955 8755
rect 1055 8705 1105 8755
rect 2675 8705 2725 8755
rect 2825 8705 2875 8755
rect 2975 8705 3025 8755
rect 4595 8705 4645 8755
rect 4745 8705 4795 8755
rect 4895 8705 4945 8755
rect 6815 8705 6865 8755
rect 6965 8705 7015 8755
rect 7115 8705 7165 8755
rect 8735 8705 8785 8755
rect 8885 8705 8935 8755
rect 9035 8705 9085 8755
rect 755 8555 805 8605
rect 905 8555 955 8605
rect 1055 8555 1105 8605
rect 2675 8555 2725 8605
rect 2825 8555 2875 8605
rect 2975 8555 3025 8605
rect 4595 8555 4645 8605
rect 4745 8555 4795 8605
rect 4895 8555 4945 8605
rect 6815 8555 6865 8605
rect 6965 8555 7015 8605
rect 7115 8555 7165 8605
rect 8735 8555 8785 8605
rect 8885 8555 8935 8605
rect 9035 8555 9085 8605
rect 1715 8165 1765 8215
rect 1865 8165 1915 8215
rect 2015 8165 2065 8215
rect 3635 8165 3685 8215
rect 3785 8165 3835 8215
rect 3935 8165 3985 8215
rect 5855 8165 5905 8215
rect 6005 8165 6055 8215
rect 6155 8165 6205 8215
rect 7775 8165 7825 8215
rect 7925 8165 7975 8215
rect 8075 8165 8125 8215
rect 9695 8165 9745 8215
rect 9845 8165 9895 8215
rect 9995 8165 10045 8215
rect 1715 8015 1765 8065
rect 1865 8015 1915 8065
rect 2015 8015 2065 8065
rect 3635 8015 3685 8065
rect 3785 8015 3835 8065
rect 3935 8015 3985 8065
rect 5855 8015 5905 8065
rect 6005 8015 6055 8065
rect 6155 8015 6205 8065
rect 7775 8015 7825 8065
rect 7925 8015 7975 8065
rect 8075 8015 8125 8065
rect 9695 8015 9745 8065
rect 9845 8015 9895 8065
rect 9995 8015 10045 8065
rect 1715 7865 1765 7915
rect 1865 7865 1915 7915
rect 2015 7865 2065 7915
rect 3635 7865 3685 7915
rect 3785 7865 3835 7915
rect 3935 7865 3985 7915
rect 5855 7865 5905 7915
rect 6005 7865 6055 7915
rect 6155 7865 6205 7915
rect 7775 7865 7825 7915
rect 7925 7865 7975 7915
rect 8075 7865 8125 7915
rect 9695 7865 9745 7915
rect 9845 7865 9895 7915
rect 9995 7865 10045 7915
rect 1715 7715 1765 7765
rect 1865 7715 1915 7765
rect 2015 7715 2065 7765
rect 3635 7715 3685 7765
rect 3785 7715 3835 7765
rect 3935 7715 3985 7765
rect 5855 7715 5905 7765
rect 6005 7715 6055 7765
rect 6155 7715 6205 7765
rect 7775 7715 7825 7765
rect 7925 7715 7975 7765
rect 8075 7715 8125 7765
rect 9695 7715 9745 7765
rect 9845 7715 9895 7765
rect 9995 7715 10045 7765
rect 1715 7565 1765 7615
rect 1865 7565 1915 7615
rect 2015 7565 2065 7615
rect 3635 7565 3685 7615
rect 3785 7565 3835 7615
rect 3935 7565 3985 7615
rect 5855 7565 5905 7615
rect 6005 7565 6055 7615
rect 6155 7565 6205 7615
rect 7775 7565 7825 7615
rect 7925 7565 7975 7615
rect 8075 7565 8125 7615
rect 9695 7565 9745 7615
rect 9845 7565 9895 7615
rect 9995 7565 10045 7615
rect 755 6905 805 6955
rect 905 6905 955 6955
rect 1055 6905 1105 6955
rect 2675 6905 2725 6955
rect 2825 6905 2875 6955
rect 2975 6905 3025 6955
rect 4595 6905 4645 6955
rect 4745 6905 4795 6955
rect 4895 6905 4945 6955
rect 6815 6905 6865 6955
rect 6965 6905 7015 6955
rect 7115 6905 7165 6955
rect 8735 6905 8785 6955
rect 8885 6905 8935 6955
rect 9035 6905 9085 6955
rect 755 6755 805 6805
rect 905 6755 955 6805
rect 1055 6755 1105 6805
rect 2675 6755 2725 6805
rect 2825 6755 2875 6805
rect 2975 6755 3025 6805
rect 4595 6755 4645 6805
rect 4745 6755 4795 6805
rect 4895 6755 4945 6805
rect 6815 6755 6865 6805
rect 6965 6755 7015 6805
rect 7115 6755 7165 6805
rect 8735 6755 8785 6805
rect 8885 6755 8935 6805
rect 9035 6755 9085 6805
rect 755 6605 805 6655
rect 905 6605 955 6655
rect 1055 6605 1105 6655
rect 2675 6605 2725 6655
rect 2825 6605 2875 6655
rect 2975 6605 3025 6655
rect 4595 6605 4645 6655
rect 4745 6605 4795 6655
rect 4895 6605 4945 6655
rect 6815 6605 6865 6655
rect 6965 6605 7015 6655
rect 7115 6605 7165 6655
rect 8735 6605 8785 6655
rect 8885 6605 8935 6655
rect 9035 6605 9085 6655
rect 1715 6215 1765 6265
rect 1865 6215 1915 6265
rect 2015 6215 2065 6265
rect 3635 6215 3685 6265
rect 3785 6215 3835 6265
rect 3935 6215 3985 6265
rect 5855 6215 5905 6265
rect 6005 6215 6055 6265
rect 6155 6215 6205 6265
rect 7775 6215 7825 6265
rect 7925 6215 7975 6265
rect 8075 6215 8125 6265
rect 9695 6215 9745 6265
rect 9845 6215 9895 6265
rect 9995 6215 10045 6265
rect 1715 6065 1765 6115
rect 1865 6065 1915 6115
rect 2015 6065 2065 6115
rect 3635 6065 3685 6115
rect 3785 6065 3835 6115
rect 3935 6065 3985 6115
rect 5855 6065 5905 6115
rect 6005 6065 6055 6115
rect 6155 6065 6205 6115
rect 7775 6065 7825 6115
rect 7925 6065 7975 6115
rect 8075 6065 8125 6115
rect 9695 6065 9745 6115
rect 9845 6065 9895 6115
rect 9995 6065 10045 6115
rect 1715 5915 1765 5965
rect 1865 5915 1915 5965
rect 2015 5915 2065 5965
rect 3635 5915 3685 5965
rect 3785 5915 3835 5965
rect 3935 5915 3985 5965
rect 5855 5915 5905 5965
rect 6005 5915 6055 5965
rect 6155 5915 6205 5965
rect 7775 5915 7825 5965
rect 7925 5915 7975 5965
rect 8075 5915 8125 5965
rect 9695 5915 9745 5965
rect 9845 5915 9895 5965
rect 9995 5915 10045 5965
rect 1715 5765 1765 5815
rect 1865 5765 1915 5815
rect 2015 5765 2065 5815
rect 3635 5765 3685 5815
rect 3785 5765 3835 5815
rect 3935 5765 3985 5815
rect 5855 5765 5905 5815
rect 6005 5765 6055 5815
rect 6155 5765 6205 5815
rect 7775 5765 7825 5815
rect 7925 5765 7975 5815
rect 8075 5765 8125 5815
rect 9695 5765 9745 5815
rect 9845 5765 9895 5815
rect 9995 5765 10045 5815
rect 1715 5615 1765 5665
rect 1865 5615 1915 5665
rect 2015 5615 2065 5665
rect 3635 5615 3685 5665
rect 3785 5615 3835 5665
rect 3935 5615 3985 5665
rect 5855 5615 5905 5665
rect 6005 5615 6055 5665
rect 6155 5615 6205 5665
rect 7775 5615 7825 5665
rect 7925 5615 7975 5665
rect 8075 5615 8125 5665
rect 9695 5615 9745 5665
rect 9845 5615 9895 5665
rect 9995 5615 10045 5665
rect 755 4955 805 5005
rect 905 4955 955 5005
rect 1055 4955 1105 5005
rect 2675 4955 2725 5005
rect 2825 4955 2875 5005
rect 2975 4955 3025 5005
rect 4595 4955 4645 5005
rect 4745 4955 4795 5005
rect 4895 4955 4945 5005
rect 6815 4955 6865 5005
rect 6965 4955 7015 5005
rect 7115 4955 7165 5005
rect 8735 4955 8785 5005
rect 8885 4955 8935 5005
rect 9035 4955 9085 5005
rect 755 4805 805 4855
rect 905 4805 955 4855
rect 1055 4805 1105 4855
rect 2675 4805 2725 4855
rect 2825 4805 2875 4855
rect 2975 4805 3025 4855
rect 4595 4805 4645 4855
rect 4745 4805 4795 4855
rect 4895 4805 4945 4855
rect 6815 4805 6865 4855
rect 6965 4805 7015 4855
rect 7115 4805 7165 4855
rect 8735 4805 8785 4855
rect 8885 4805 8935 4855
rect 9035 4805 9085 4855
rect 755 4655 805 4705
rect 905 4655 955 4705
rect 1055 4655 1105 4705
rect 2675 4655 2725 4705
rect 2825 4655 2875 4705
rect 2975 4655 3025 4705
rect 4595 4655 4645 4705
rect 4745 4655 4795 4705
rect 4895 4655 4945 4705
rect 6815 4655 6865 4705
rect 6965 4655 7015 4705
rect 7115 4655 7165 4705
rect 8735 4655 8785 4705
rect 8885 4655 8935 4705
rect 9035 4655 9085 4705
rect 1715 4115 1765 4165
rect 1865 4115 1915 4165
rect 2015 4115 2065 4165
rect 3635 4115 3685 4165
rect 3785 4115 3835 4165
rect 3935 4115 3985 4165
rect 5855 4115 5905 4165
rect 6005 4115 6055 4165
rect 6155 4115 6205 4165
rect 7775 4115 7825 4165
rect 7925 4115 7975 4165
rect 8075 4115 8125 4165
rect 9695 4115 9745 4165
rect 9845 4115 9895 4165
rect 9995 4115 10045 4165
rect 1715 3965 1765 4015
rect 1865 3965 1915 4015
rect 2015 3965 2065 4015
rect 3635 3965 3685 4015
rect 3785 3965 3835 4015
rect 3935 3965 3985 4015
rect 5855 3965 5905 4015
rect 6005 3965 6055 4015
rect 6155 3965 6205 4015
rect 7775 3965 7825 4015
rect 7925 3965 7975 4015
rect 8075 3965 8125 4015
rect 9695 3965 9745 4015
rect 9845 3965 9895 4015
rect 9995 3965 10045 4015
rect 755 3605 805 3655
rect 905 3605 955 3655
rect 1055 3605 1105 3655
rect 2675 3605 2725 3655
rect 2825 3605 2875 3655
rect 2975 3605 3025 3655
rect 4595 3605 4645 3655
rect 4745 3605 4795 3655
rect 4895 3605 4945 3655
rect 6815 3605 6865 3655
rect 6965 3605 7015 3655
rect 7115 3605 7165 3655
rect 8735 3605 8785 3655
rect 8885 3605 8935 3655
rect 9035 3605 9085 3655
rect 755 3455 805 3505
rect 905 3455 955 3505
rect 1055 3455 1105 3505
rect 2675 3455 2725 3505
rect 2825 3455 2875 3505
rect 2975 3455 3025 3505
rect 4595 3455 4645 3505
rect 4745 3455 4795 3505
rect 4895 3455 4945 3505
rect 6815 3455 6865 3505
rect 6965 3455 7015 3505
rect 7115 3455 7165 3505
rect 8735 3455 8785 3505
rect 8885 3455 8935 3505
rect 9035 3455 9085 3505
rect 755 2225 805 2275
rect 905 2225 955 2275
rect 1055 2225 1105 2275
rect 8735 2225 8785 2275
rect 8885 2225 8935 2275
rect 9035 2225 9085 2275
rect 755 2075 805 2125
rect 905 2075 955 2125
rect 1055 2075 1105 2125
rect 8735 2075 8785 2125
rect 8885 2075 8935 2125
rect 9035 2075 9085 2125
rect 755 1925 805 1975
rect 905 1925 955 1975
rect 1055 1925 1105 1975
rect 8735 1925 8785 1975
rect 8885 1925 8935 1975
rect 9035 1925 9085 1975
rect 755 1775 805 1825
rect 905 1775 955 1825
rect 1055 1775 1105 1825
rect 8735 1775 8785 1825
rect 8885 1775 8935 1825
rect 9035 1775 9085 1825
rect 755 1625 805 1675
rect 905 1625 955 1675
rect 1055 1625 1105 1675
rect 8735 1625 8785 1675
rect 8885 1625 8935 1675
rect 9035 1625 9085 1675
rect 755 215 805 265
rect 905 215 955 265
rect 1055 215 1105 265
rect 2675 215 2725 265
rect 2825 215 2875 265
rect 2975 215 3025 265
rect 4595 215 4645 265
rect 4745 215 4795 265
rect 4895 215 4945 265
rect 6815 215 6865 265
rect 6965 215 7015 265
rect 7115 215 7165 265
rect 8735 215 8785 265
rect 8885 215 8935 265
rect 9035 215 9085 265
rect 755 65 805 115
rect 905 65 955 115
rect 1055 65 1105 115
rect 2675 65 2725 115
rect 2825 65 2875 115
rect 2975 65 3025 115
rect 4595 65 4645 115
rect 4745 65 4795 115
rect 4895 65 4945 115
rect 6815 65 6865 115
rect 6965 65 7015 115
rect 7115 65 7165 115
rect 8735 65 8785 115
rect 8885 65 8935 115
rect 9035 65 9085 115
<< pad >>
rect 1655 23315 9145 30805
<< metal3 >>
rect 1655 23315 9145 30805
<< pseudo_rnwell >>
rect 2400 1410 2430 2130
rect 8370 1410 8400 2130
<< rnwell >>
rect 2430 1410 8370 2130
<< labels >>
flabel metal1 s 4350 21330 4350 21330 2 FreeSans 400 0 0 0 pad
port 1 ne
flabel metal1 s 5340 120 5340 120 2 FreeSans 400 0 0 0 xpad
port 2 ne
flabel metal2 s 10200 3570 10200 3570 2 FreeSans 400 0 0 0 vss
flabel metal2 s 10200 13290 10200 13290 2 FreeSans 400 0 0 0 vss
port 7 ne
flabel metal2 s 10200 11970 10200 11970 2 FreeSans 400 0 0 0 vss
flabel metal2 s 10080 10740 10080 10740 2 FreeSans 400 0 0 0 vss
flabel metal2 s 10200 11430 10200 11430 2 FreeSans 400 0 0 0 vdd
flabel metal2 s 10200 12780 10200 12780 2 FreeSans 400 0 0 0 vdd
flabel metal2 s 10080 13980 10080 13980 2 FreeSans 400 0 0 0 vdd
port 6 ne
flabel rnwell s 5040 1710 5040 1710 2 FreeSans 400 0 0 0 r0_body
flabel nwell s -60 3930 -60 3930 2 FreeSans 400 0 0 0 vdd
flabel metal2 s 8520 150 8520 150 2 FreeSans 400 0 0 0 vss
<< checkpaint >>
rect -100 -70 10900 31120
<< end >>
