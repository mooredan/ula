magic
tech amic5n
timestamp 1609902395
<< checkpaint >>
rect 224000 257200 501000 501000
rect 224400 -1000 501000 257200
<< metal1 >>
rect 0 0 500000 500000
<< end >>
