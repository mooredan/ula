`celldefine
module decap5 ();
endmodule
`endcelldefine
