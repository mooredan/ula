`celldefine
module buf_b (z, a);
  output z;
  input  a;

  buf G1 (z, a);
endmodule
`endcelldefine
