* Output transition times
.include mag/pad_nwellres.cir
.include mag/inv_e.cir
.include mag/nand2_c.cir
.include mag/nor2_c.cir
.include mag/subc_2.cir

.lib device_models/AMI_C5N.lib TT
.lib device_models/AMI_C5N_rmodels.lib NOM 

.temp 25

.param VDD_VAL=5

* power supply
vvdd vdd 0 DC VDD_VAL
vvss vss 0 DC 0

* what sort of pre driver is needed here
* target is around 7-10ns rise/fall at the
* output of the big driver fets 80% of VDD
*  
* predriver needs to be function of break-before-make
* and fast going into tri-state
* vpd  pd  0 DC 0 PULSE(0 3 10n 4.8n 4.8n 80n 220n)
* vnpu npu 0 DC 0 PULSE(0 3 10n 4.8n 4.8n 80n 220n)


* .subckt pad_nwellres pad xpad anpu apd tri ntri vdd vss
xdut                   pad xpad a    a   vss vdd  vdd vss pad_nwellres



* vnpd  npd 0 DC 0 PULSE(0 {VDD_VAL} 10n 4.8n 4.8n 80n 220n)
* va    a 0 DC 0 PULSE(0 {VDD_VAL} 10n 4.8n 4.8n 80n 220n)
va    a 0 DC 0 PULSE(0 {VDD_VAL} 10n 4.8n 4.8n 45.2n 100n)


* npu and pd are the gate connections to the
* driver FETs
*
* these need to turn into gates for tristate
*
* MP11 npu a  vdd vdd  pfet w=6.0u   l=0.6u
* MN11 npu a  vss vss  nfet w=3.0u   l=0.6u
*
*
* MP10 pd a  vdd vdd  pfet w=7.5u   l=0.6u
* MN10 pd a  vss vss  nfet w=2.7u   l=0.6u

*.subckt inv_c z a vdd vss
* XNPU npu a vdd vss inv_e
* XPD   pd a vdd vss inv_e




* output load
cpad pad vgnd 50p
vvgnd vgnd 0 DC 0

* add small load to core side of the
* input series resistor


.save all

.tran 0.1n 900n

.control
destroy all
run

setplot tran1
plot v(xdut.npu) v(pad)
plot  v(xdut.pd)  v(pad)

let vdd_max = maximum(v(vdd))
let vol = vdd_max * 0.1
let voh = vdd_max * 0.9

print vdd_max
print vol
print voh


meas tran nputlh TRIG v(xdut.npu) VAL=vol RISE=1 TARG v(xdut.npu) VAL=voh RISE=1
meas tran nputhl TRIG v(xdut.npu) VAL=voh FALL=2 TARG v(xdut.npu) VAL=vol FALL=2
meas tran padtlh TRIG v(pad) VAL=vol RISE=2 TARG v(pad) VAL=voh RISE=2

meas tran pdtlh TRIG v(xdut.pd) VAL=vol RISE=1 TARG v(xdut.pd) VAL=voh RISE=1
meas tran pdthl TRIG v(xdut.pd) VAL=voh FALL=2 TARG v(xdut.pd) VAL=vol FALL=2
meas tran padthl TRIG v(pad) VAL=voh FALL=1 TARG v(pad) VAL=vol FALL=1

.endc

.end
