magic
tech scmos
timestamp 1591539050
<< nwell >>
rect -1 29 43 81
<< nselect >>
rect 15 2 29 25
<< pselect >>
rect 12 33 33 77
<< ntransistor >>
rect 21 4 23 23
<< ptransistor >>
rect 20 35 22 75
<< ndiffusion >>
rect 17 4 21 23
rect 23 4 27 23
<< pdiffusion >>
rect 14 35 20 75
rect 22 35 31 75
<< polysilicon >>
rect 20 75 22 77
rect 20 33 22 35
rect 21 23 23 30
rect 21 2 23 4
<< metal1 >>
rect 5 76 37 79
rect 6 69 9 73
rect 33 69 36 73
rect 6 62 9 66
rect 33 62 36 66
rect 6 55 9 59
rect 33 55 36 59
rect 6 48 9 52
rect 33 48 36 52
rect 6 41 9 45
rect 33 41 36 45
rect 6 34 9 38
rect 33 34 36 38
rect 6 27 9 31
rect 33 27 36 31
rect 6 20 9 24
rect 33 20 36 24
rect 6 13 9 17
rect 33 13 36 17
rect 6 6 9 10
rect 33 6 36 10
rect 5 0 37 3
rect -2 -10 2 -3
rect 5 -10 9 -3
rect 12 -10 16 -3
rect 19 -10 23 -3
rect 26 -10 30 -3
rect 33 -10 37 -3
rect 40 -10 44 -3
<< bb >>
rect 0 0 42 79
<< labels >>
rlabel metal1 5 0 5 0 2 Gnd
port 3 ne
rlabel nwell 5 30 5 30 2 Vdd
rlabel metal1 5 76 5 76 2 Vdd
port 2 ne
<< end >>
