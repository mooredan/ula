* Transient analysis of 

.include cell.cir

.lib ../../device_models/AMI_C5N.lib TT

.param VDD_VAL=5.0
.param FREQ=50.0Meg
.param PER={1 / FREQ}
.param pwrtime = 5e-9
.param TT=50p
.param CA=1f
.param CB=1f
.param CZ=1f

.csparam v_vdd = {VDD_VAL}
.csparam t_per = {PER}
.csparam pwrt = {pwrtime}

* power supply
Vvdd vdd 0 DC {VDD_VAL} PWL( 0 0  {pwrtime / 3}  0  {pwrtime * 2 / 3} {VDD_VAL})
Vvss vss 0 DC 0

* input a
Va   a_s 0 DC 0 PWL (                  0      0 
+                    {pwrtime + PER *  2}          0
+                    {pwrtime + PER *  2 + TT}  {VDD_VAL}
+                    {pwrtime + PER *  3}       {VDD_VAL} 
+                    {pwrtime + PER *  3 + TT}     0
+                    {pwrtime + PER *  4}          0
+                    {pwrtime + PER *  4 + TT}  {VDD_VAL}
+                   )
Ra_s a_s a 100
Ca   a   0 {CA} 


* input b
Vb   b_s 0 DC 0 PWL (                  0      0 
+                    {pwrtime + PER *  1}          0
+                    {pwrtime + PER *  1 + TT}  {VDD_VAL}
+                    {pwrtime + PER *  4}       {VDD_VAL} 
+                    {pwrtime + PER *  4 + TT}     0
+                    {pwrtime + PER *  5}          0
+                    {pwrtime + PER *  5 + TT}  {VDD_VAL}
+                    {pwrtime + PER *  6}       {VDD_VAL} 
+                    {pwrtime + PER *  6 + TT}     0
+                   )

Rb_s b_s b 100
Cb   b   0 {CA} 

* DUT
Xdut z a b vdd vss and2_b

* output load
Cz z 0 {CZ} 


* sweep transition time from : ~30ps  to: ~1.3 ns
*
*              cck (pF)         rise (ps)
*              ===========================
*              0.001               30.8 
*              0.5                 79.2
*              1.0                146.8 
*              2.5                355.8  
*              5.0                702.2
*             10.0               1395.2
*
* sweep output load     from : 10 fF   to: 2 pF  - seven loads

.control
  let vol  = $&v_vdd * 0.20
  set vol  = "$&vol"

  let voh  = $&v_vdd * 0.80
  set voh  = "$&voh"

  let vmid = $&v_vdd * 0.50
  set vmid = "$&vmid"

  let idx1 = 0
  set idx1 = "$&idx1"

  let t_per = $&t_per
  set t_per = "$&t_per"

  let ptime = $&pwrt
  set ptime = "$&ptime"

  foreach in_load 10e-15 500e-15 1e-12 3e-12 5e-12
  * foreach in_load 1e-15

     let idx2 = 0
     set idx2 = "$&idx2"

     foreach out_load 10e-15 50e-15 100e-15 250e-15 500e-15
     * foreach out_load 0.010e-12

      destroy all

      alter ca $in_load
      alter cb $in_load
      alter cz $out_load

      * run
      let tstop = ptime + $t_per * 7 
      set tstop = "$&tstop"
      tran 10p $tstop

      * echo in_load: $in_load
      * echo out_load: $out_load

      ************************************************************************************
      * a rising to z rising 
      ************************************************************************************
      meas tran tt__a_rise1 TRIG v(a) VAL=vol RISE=1 TARG v(a) VAL=voh RISE=1 
      meas tran tt__z_rise1 TRIG v(z) VAL=vol RISE=1 TARG v(z) VAL=voh RISE=1 
      meas tran td__a_rise1__z_rise1 TRIG v(a) VAL=vmid RISE=1 TARG v(z) VAL=vmid RISE=1

      let dtime = td__a_rise1__z_rise1
      set dtime = "$&dtime"
      let ittime = tt__a_rise1
      set ittime = "$&ittime"
      let ttime = tt__z_rise1
      set ttime = "$&ttime"
      echo delay: a_rise__z_rise $idx1 $idx2 in_rise: $ittime  out_load: $out_load  time: $dtime
      echo trans: a_rise__z_rise $idx1 $idx2 in_rise: $ittime  out_load: $out_load  time: $ttime



      ************************************************************************************
      * a falling to z falling 
      ************************************************************************************
      meas tran tt__a_fall1 TRIG v(a) VAL=voh FALL=1 TARG v(a) VAL=vol FALL=1 
      meas tran tt__z_fall1 TRIG v(z) VAL=voh FALL=1 TARG v(z) VAL=vol FALL=1 
      meas tran td__a_fall1__z_fall1 TRIG v(a) VAL=vmid FALL=1 TARG v(z) VAL=vmid FALL=1

      let dtime = td__a_fall1__z_fall1
      set dtime = "$&dtime"
      let ittime = tt__a_fall1
      set ittime = "$&ittime"
      let ttime = tt__z_fall1
      set ttime = "$&ttime"
      echo delay: a_fall__z_fall $idx1 $idx2 in_fall: $ittime  out_load: $out_load  time: $dtime
      echo trans: a_fall__z_fall $idx1 $idx2 in_fall: $ittime  out_load: $out_load  time: $ttime


      ************************************************************************************
      * b rising to z rising 
      ************************************************************************************
      meas tran tt__b_rise2 TRIG v(b) VAL=vol RISE=2 TARG v(b) VAL=voh RISE=2 
      meas tran tt__z_rise2 TRIG v(z) VAL=vol RISE=2 TARG v(z) VAL=voh RISE=2 
      meas tran td__b_rise2__z_rise2 TRIG v(b) VAL=vmid RISE=2 TARG v(z) VAL=vmid RISE=2

      let dtime = td__b_rise2__z_rise2
      set dtime = "$&dtime"
      let ittime = tt__b_rise2
      set ittime = "$&ittime"
      let ttime = tt__z_rise2
      set ttime = "$&ttime"
      echo delay: b_rise__z_rise $idx1 $idx2 in_rise: $ittime  out_load: $out_load  time: $dtime
      echo trans: b_rise__z_rise $idx1 $idx2 in_rise: $ittime  out_load: $out_load  time: $ttime


      ************************************************************************************
      * b falling to z falling
      ************************************************************************************
      meas tran tt__b_fall2 TRIG v(b) VAL=voh FALL=2 TARG v(b) VAL=vol FALL=2 
      meas tran tt__z_fall2 TRIG v(z) VAL=voh FALL=2 TARG v(z) VAL=vol FALL=2 
      meas tran td__b_fall2__z_fall2 TRIG v(b) VAL=vmid FALL=2 TARG v(z) VAL=vmid FALL=2

      let dtime = td__b_fall2__z_fall2
      set dtime = "$&dtime"
      let ittime = tt__b_fall2
      set ittime = "$&ittime"
      let ttime = tt__z_fall2
      set ttime = "$&ttime"
      echo delay: b_fall__z_fall $idx1 $idx2 in_fall: $ittime  out_load: $out_load  time: $dtime
      echo trans: b_fall__z_fall $idx1 $idx2 in_fall: $ittime  out_load: $out_load  time: $ttime


      let idx2 = idx2 + 1
      set idx2 = "$&idx2"

    end
    let idx1 = idx1 + 1
    set idx1 = "$&idx1"
  end

* setplot tran1
* plot v(vdd) v(a) v(b) v(z)
* plot v(a)
* plot v(z)

  ***********************************
  * Do input capacitance measurements
  ***********************************
  let vmid = $&v_vdd * 0.5
  set vmid = "$&vmid"
  
  alter ca 0
  alter cb 0
  alter cz 0
  
  * alter vvdd  dc 5.0
  alter vvdd  dc $&v_vdd
  alter va    dc $vmid
  alter vb    dc $vmid
  
  let idx = 70
  set idx = "$&idx"
  
  ***********************************
  * set up and measure input pin a
  ***********************************
  alter va ac 1.0
  
  ac dec 10 1 100e6
  
  let freq = real(frequency[$idx])
  set freq = "$&freq"
  
  let a_cap = '1.0 / (imag(v(a)[$idx] / i(va)[$idx]) * 2 * pi * real(frequency[$idx]))'
  set a_cap = "$&a_cap"
  echo incap: pin: a cap: $a_cap  freq: $freq
  
  ***********************************
  * set up and measure input pin b
  ***********************************
  alter va ac 0.0
  alter vb ac 1.0
  
  ac dec 10 1 100e6
  
  let freq = real(frequency[$idx])
  set freq = "$&freq"
  
  let b_cap = '1.0 / (imag(v(b)[$idx] / i(vb)[$idx]) * 2 * pi * real(frequency[$idx]))'
  set b_cap = "$&b_cap"
  echo incap: pin: b cap: $b_cap  freq: $freq

  quit 0
.endc

.end
