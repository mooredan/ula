magic
tech amic5n
timestamp 1608317705
<< nwell >>
rect 3480 900 5250 2430
<< ntransistor >>
rect 4230 120 4290 720
<< ptransistor >>
rect 4200 1080 4260 2250
rect 4470 1080 4530 2250
<< ndiffusion >>
rect 4110 120 4230 720
rect 4290 120 4410 720
<< pdiffusion >>
rect 4020 1080 4200 2250
rect 4260 1080 4470 2250
rect 4530 1080 4740 2250
<< polysilicon >>
rect 4200 2250 4260 2310
rect 4470 2250 4530 2310
rect 4200 1020 4260 1080
rect 4470 1020 4530 1080
rect 4230 720 4290 900
rect 4230 60 4290 120
<< metal1 >>
rect 3600 2280 5130 2370
rect 3600 1860 3930 1980
rect 4830 1860 5130 1980
rect 3600 1650 3930 1770
rect 4830 1650 5130 1770
rect 3600 1440 3930 1560
rect 4830 1440 5130 1560
rect 3600 1230 3930 1350
rect 4830 1230 5130 1350
rect 3600 1020 3930 1140
rect 4830 1020 5130 1140
rect 3600 810 3930 930
rect 4830 810 5130 930
rect 3600 600 3870 720
rect 4800 600 5130 720
rect 3600 390 3870 510
rect 4800 390 5130 510
rect 3600 180 3870 300
rect 4800 180 5130 300
rect 3600 0 5130 90
<< labels >>
flabel metal1  3600 0 3600 0 2 FreeSans 400 0 0 0 Gnd
port 3 ne
flabel nwell  3600 900 3600 900 2 FreeSans 400 0 0 0 Vdd
flabel metal1  3600 2280 3600 2280 2 FreeSans 400 0 0 0 Vdd
port 2 ne
<< checkpaint >>
rect -10 -10 5260 2440
<< end >>
