magic
tech amic5n
timestamp 1621863012
<< error_s >>
rect 45 985 75 1005
rect 125 985 155 1005
rect 45 955 155 985
rect 245 985 275 1005
rect 325 985 365 1005
rect 245 955 365 985
rect 425 985 465 1005
rect 425 955 505 985
use subc_2  subc_2_0 ~/projects/ula/mag
timestamp 1621863012
transform 1 0 0 0 1 0
box -105 -45 305 2455
use inv_c  inv_c_0
timestamp 1621863012
transform 1 0 200 0 1 0
box -105 -45 495 2455
<< end >>
