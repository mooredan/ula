* Human Body Model
* from Kang's book
.subckt hbm out

* Simple HBM/MM circuit
*
.param level=1.0
+ nom_voltage={level * 2000} 
+ td=1n
+ tr=1p

Cc n1 0 100p
S1 n1 n2 n5 0 SW OFF
Ls n2 n3 5u
Rs n3 out 1500
Cs n3 out 1p
Ct out 0 10p

.model SW SW(Ron=1 Roff=1G Vt=0.5)
.ic v(n1)={nom_voltage} v(n2)=0 v(out)=0 

* very fast switching on 
V1 n5 0 DC 0 PULSE(0 1 {td} {tr} 1 1 2)

.ends hbm
