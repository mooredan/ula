magic
tech scmos
magscale 1 2
timestamp 1570494029
<< error_s >>
rect 2400 1940 2406 1942
rect 2404 1936 2406 1940
rect 2400 1934 2406 1936
rect 2422 1940 2430 1942
rect 2422 1936 2424 1940
rect 2428 1936 2430 1940
rect 2422 1934 2430 1936
rect 2446 1940 2454 1942
rect 2446 1936 2448 1940
rect 2452 1936 2454 1940
rect 2446 1934 2454 1936
rect 2470 1940 2478 1942
rect 2470 1936 2472 1940
rect 2476 1936 2478 1940
rect 2470 1934 2478 1936
rect 2494 1940 2502 1942
rect 2494 1936 2496 1940
rect 2500 1936 2502 1940
rect 2494 1934 2502 1936
rect 2710 1940 2718 1942
rect 2710 1936 2712 1940
rect 2716 1936 2718 1940
rect 2710 1934 2718 1936
rect 2734 1940 2742 1942
rect 2734 1936 2736 1940
rect 2740 1936 2742 1940
rect 2734 1934 2742 1936
rect 2758 1940 2766 1942
rect 2758 1936 2760 1940
rect 2764 1936 2766 1940
rect 2758 1934 2766 1936
rect 2782 1940 2790 1942
rect 2782 1936 2784 1940
rect 2788 1936 2790 1940
rect 2782 1934 2790 1936
rect 2806 1940 2814 1942
rect 2806 1936 2808 1940
rect 2812 1936 2814 1940
rect 2806 1934 2814 1936
rect 2830 1940 2838 1942
rect 2830 1936 2832 1940
rect 2836 1936 2838 1940
rect 2830 1934 2838 1936
rect 2854 1940 2862 1942
rect 2854 1936 2856 1940
rect 2860 1936 2862 1940
rect 2854 1934 2862 1936
rect 2878 1940 2886 1942
rect 2878 1936 2880 1940
rect 2884 1936 2886 1940
rect 2878 1934 2886 1936
rect 2902 1940 2910 1942
rect 2902 1936 2904 1940
rect 2908 1936 2910 1940
rect 2902 1934 2910 1936
rect 2926 1940 2934 1942
rect 2926 1936 2928 1940
rect 2932 1936 2934 1940
rect 2926 1934 2934 1936
rect 2950 1940 2958 1942
rect 2950 1936 2952 1940
rect 2956 1936 2958 1940
rect 2950 1934 2958 1936
rect 2974 1940 2982 1942
rect 2974 1936 2976 1940
rect 2980 1936 2982 1940
rect 2974 1934 2982 1936
rect 2998 1940 3006 1942
rect 2998 1936 3000 1940
rect 3004 1936 3006 1940
rect 2998 1934 3006 1936
rect 3022 1940 3030 1942
rect 3022 1936 3024 1940
rect 3028 1936 3030 1940
rect 3022 1934 3030 1936
rect 3046 1940 3054 1942
rect 3046 1936 3048 1940
rect 3052 1936 3054 1940
rect 3046 1934 3054 1936
rect 3070 1940 3078 1942
rect 3070 1936 3072 1940
rect 3076 1936 3078 1940
rect 3070 1934 3078 1936
rect 3094 1940 3102 1942
rect 3094 1936 3096 1940
rect 3100 1936 3102 1940
rect 3094 1934 3102 1936
rect 3310 1940 3318 1942
rect 3310 1936 3312 1940
rect 3316 1936 3318 1940
rect 3310 1934 3318 1936
rect 3334 1940 3342 1942
rect 3334 1936 3336 1940
rect 3340 1936 3342 1940
rect 3334 1934 3342 1936
rect 3358 1940 3366 1942
rect 3358 1936 3360 1940
rect 3364 1936 3366 1940
rect 3358 1934 3366 1936
rect 3382 1940 3390 1942
rect 3382 1936 3384 1940
rect 3388 1936 3390 1940
rect 3382 1934 3390 1936
rect 3406 1940 3414 1942
rect 3406 1936 3408 1940
rect 3412 1936 3414 1940
rect 3406 1934 3414 1936
rect 3430 1940 3438 1942
rect 3430 1936 3432 1940
rect 3436 1936 3438 1940
rect 3430 1934 3438 1936
rect 3454 1940 3462 1942
rect 3454 1936 3456 1940
rect 3460 1936 3462 1940
rect 3454 1934 3462 1936
rect 3478 1940 3486 1942
rect 3478 1936 3480 1940
rect 3484 1936 3486 1940
rect 3478 1934 3486 1936
rect 3502 1940 3510 1942
rect 3502 1936 3504 1940
rect 3508 1936 3510 1940
rect 3502 1934 3510 1936
rect 3526 1940 3534 1942
rect 3526 1936 3528 1940
rect 3532 1936 3534 1940
rect 3526 1934 3534 1936
rect 3550 1940 3558 1942
rect 3550 1936 3552 1940
rect 3556 1936 3558 1940
rect 3550 1934 3558 1936
rect 3574 1940 3582 1942
rect 3574 1936 3576 1940
rect 3580 1936 3582 1940
rect 3574 1934 3582 1936
rect 3598 1940 3606 1942
rect 3598 1936 3600 1940
rect 3604 1936 3606 1940
rect 3598 1934 3606 1936
rect 3622 1940 3630 1942
rect 3622 1936 3624 1940
rect 3628 1936 3630 1940
rect 3622 1934 3630 1936
rect 3646 1940 3654 1942
rect 3646 1936 3648 1940
rect 3652 1936 3654 1940
rect 3646 1934 3654 1936
rect 3670 1940 3678 1942
rect 3670 1936 3672 1940
rect 3676 1936 3678 1940
rect 3670 1934 3678 1936
rect 3694 1940 3702 1942
rect 3694 1936 3696 1940
rect 3700 1936 3702 1940
rect 3694 1934 3702 1936
rect 3910 1940 3918 1942
rect 3910 1936 3912 1940
rect 3916 1936 3918 1940
rect 3910 1934 3918 1936
rect 3934 1940 3942 1942
rect 3934 1936 3936 1940
rect 3940 1936 3942 1940
rect 3934 1934 3942 1936
rect 3958 1940 3966 1942
rect 3958 1936 3960 1940
rect 3964 1936 3966 1940
rect 3958 1934 3966 1936
rect 3982 1940 3990 1942
rect 3982 1936 3984 1940
rect 3988 1936 3990 1940
rect 3982 1934 3990 1936
rect 4006 1940 4014 1942
rect 4006 1936 4008 1940
rect 4012 1936 4014 1940
rect 4006 1934 4014 1936
rect 4030 1940 4038 1942
rect 4030 1936 4032 1940
rect 4036 1936 4038 1940
rect 4030 1934 4038 1936
rect 4054 1940 4062 1942
rect 4054 1936 4056 1940
rect 4060 1936 4062 1940
rect 4054 1934 4062 1936
rect 4078 1940 4086 1942
rect 4078 1936 4080 1940
rect 4084 1936 4086 1940
rect 4078 1934 4086 1936
rect 4102 1940 4110 1942
rect 4102 1936 4104 1940
rect 4108 1936 4110 1940
rect 4102 1934 4110 1936
rect 4126 1940 4134 1942
rect 4126 1936 4128 1940
rect 4132 1936 4134 1940
rect 4126 1934 4134 1936
rect 4150 1940 4158 1942
rect 4150 1936 4152 1940
rect 4156 1936 4158 1940
rect 4150 1934 4158 1936
rect 4174 1940 4182 1942
rect 4174 1936 4176 1940
rect 4180 1936 4182 1940
rect 4174 1934 4182 1936
rect 4198 1940 4206 1942
rect 4198 1936 4200 1940
rect 4204 1936 4206 1940
rect 4198 1934 4206 1936
rect 4222 1940 4230 1942
rect 4222 1936 4224 1940
rect 4228 1936 4230 1940
rect 4222 1934 4230 1936
rect 4246 1940 4254 1942
rect 4246 1936 4248 1940
rect 4252 1936 4254 1940
rect 4246 1934 4254 1936
rect 4270 1940 4278 1942
rect 4270 1936 4272 1940
rect 4276 1936 4278 1940
rect 4270 1934 4278 1936
rect 4294 1940 4302 1942
rect 4294 1936 4296 1940
rect 4300 1936 4302 1940
rect 4294 1934 4302 1936
rect 4510 1940 4518 1942
rect 4510 1936 4512 1940
rect 4516 1936 4518 1940
rect 4510 1934 4518 1936
rect 4534 1940 4542 1942
rect 4534 1936 4536 1940
rect 4540 1936 4542 1940
rect 4534 1934 4542 1936
rect 4558 1940 4566 1942
rect 4558 1936 4560 1940
rect 4564 1936 4566 1940
rect 4558 1934 4566 1936
rect 4582 1940 4590 1942
rect 4582 1936 4584 1940
rect 4588 1936 4590 1940
rect 4582 1934 4590 1936
rect 4606 1940 4614 1942
rect 4606 1936 4608 1940
rect 4612 1936 4614 1940
rect 4606 1934 4614 1936
rect 4630 1940 4638 1942
rect 4630 1936 4632 1940
rect 4636 1936 4638 1940
rect 4630 1934 4638 1936
rect 4654 1940 4662 1942
rect 4654 1936 4656 1940
rect 4660 1936 4662 1940
rect 4654 1934 4662 1936
rect 4678 1940 4686 1942
rect 4678 1936 4680 1940
rect 4684 1936 4686 1940
rect 4678 1934 4686 1936
rect 4702 1940 4710 1942
rect 4702 1936 4704 1940
rect 4708 1936 4710 1940
rect 4702 1934 4710 1936
rect 4726 1940 4734 1942
rect 4726 1936 4728 1940
rect 4732 1936 4734 1940
rect 4726 1934 4734 1936
rect 4750 1940 4758 1942
rect 4750 1936 4752 1940
rect 4756 1936 4758 1940
rect 4750 1934 4758 1936
rect 4774 1940 4782 1942
rect 4774 1936 4776 1940
rect 4780 1936 4782 1940
rect 4774 1934 4782 1936
rect 4798 1934 4800 1942
rect 5710 1940 5718 1942
rect 5710 1936 5712 1940
rect 5716 1936 5718 1940
rect 5710 1934 5718 1936
rect 5734 1940 5742 1942
rect 5734 1936 5736 1940
rect 5740 1936 5742 1940
rect 5734 1934 5742 1936
rect 5758 1940 5766 1942
rect 5758 1936 5760 1940
rect 5764 1936 5766 1940
rect 5758 1934 5766 1936
rect 5782 1940 5790 1942
rect 5782 1936 5784 1940
rect 5788 1936 5790 1940
rect 5782 1934 5790 1936
rect 5806 1940 5814 1942
rect 5806 1936 5808 1940
rect 5812 1936 5814 1940
rect 5806 1934 5814 1936
rect 5830 1940 5838 1942
rect 5830 1936 5832 1940
rect 5836 1936 5838 1940
rect 5830 1934 5838 1936
rect 5854 1940 5862 1942
rect 5854 1936 5856 1940
rect 5860 1936 5862 1940
rect 5854 1934 5862 1936
rect 5878 1940 5886 1942
rect 5878 1936 5880 1940
rect 5884 1936 5886 1940
rect 5878 1934 5886 1936
rect 5902 1940 5910 1942
rect 5902 1936 5904 1940
rect 5908 1936 5910 1940
rect 5902 1934 5910 1936
rect 5926 1940 5934 1942
rect 5926 1936 5928 1940
rect 5932 1936 5934 1940
rect 5926 1934 5934 1936
rect 5950 1940 5958 1942
rect 5950 1936 5952 1940
rect 5956 1936 5958 1940
rect 5950 1934 5958 1936
rect 5974 1940 5982 1942
rect 5974 1936 5976 1940
rect 5980 1936 5982 1940
rect 5974 1934 5982 1936
rect 5998 1940 6006 1942
rect 5998 1936 6000 1940
rect 6004 1936 6006 1940
rect 5998 1934 6006 1936
rect 6022 1940 6030 1942
rect 6022 1936 6024 1940
rect 6028 1936 6030 1940
rect 6022 1934 6030 1936
rect 6046 1940 6054 1942
rect 6046 1936 6048 1940
rect 6052 1936 6054 1940
rect 6046 1934 6054 1936
rect 6070 1940 6078 1942
rect 6070 1936 6072 1940
rect 6076 1936 6078 1940
rect 6070 1934 6078 1936
rect 6094 1940 6102 1942
rect 6094 1936 6096 1940
rect 6100 1936 6102 1940
rect 6094 1934 6102 1936
rect 6310 1940 6318 1942
rect 6310 1936 6312 1940
rect 6316 1936 6318 1940
rect 6310 1934 6318 1936
rect 6334 1940 6342 1942
rect 6334 1936 6336 1940
rect 6340 1936 6342 1940
rect 6334 1934 6342 1936
rect 6358 1940 6366 1942
rect 6358 1936 6360 1940
rect 6364 1936 6366 1940
rect 6358 1934 6366 1936
rect 6382 1940 6390 1942
rect 6382 1936 6384 1940
rect 6388 1936 6390 1940
rect 6382 1934 6390 1936
rect 6406 1940 6414 1942
rect 6406 1936 6408 1940
rect 6412 1936 6414 1940
rect 6406 1934 6414 1936
rect 6430 1940 6438 1942
rect 6430 1936 6432 1940
rect 6436 1936 6438 1940
rect 6430 1934 6438 1936
rect 6454 1940 6462 1942
rect 6454 1936 6456 1940
rect 6460 1936 6462 1940
rect 6454 1934 6462 1936
rect 6478 1940 6486 1942
rect 6478 1936 6480 1940
rect 6484 1936 6486 1940
rect 6478 1934 6486 1936
rect 6502 1940 6510 1942
rect 6502 1936 6504 1940
rect 6508 1936 6510 1940
rect 6502 1934 6510 1936
rect 6526 1940 6534 1942
rect 6526 1936 6528 1940
rect 6532 1936 6534 1940
rect 6526 1934 6534 1936
rect 6550 1940 6558 1942
rect 6550 1936 6552 1940
rect 6556 1936 6558 1940
rect 6550 1934 6558 1936
rect 6574 1940 6582 1942
rect 6574 1936 6576 1940
rect 6580 1936 6582 1940
rect 6574 1934 6582 1936
rect 6598 1940 6606 1942
rect 6598 1936 6600 1940
rect 6604 1936 6606 1940
rect 6598 1934 6606 1936
rect 6622 1940 6630 1942
rect 6622 1936 6624 1940
rect 6628 1936 6630 1940
rect 6622 1934 6630 1936
rect 6646 1940 6654 1942
rect 6646 1936 6648 1940
rect 6652 1936 6654 1940
rect 6646 1934 6654 1936
rect 6670 1940 6678 1942
rect 6670 1936 6672 1940
rect 6676 1936 6678 1940
rect 6670 1934 6678 1936
rect 6694 1940 6702 1942
rect 6694 1936 6696 1940
rect 6700 1936 6702 1940
rect 6694 1934 6702 1936
rect 6910 1940 6918 1942
rect 6910 1936 6912 1940
rect 6916 1936 6918 1940
rect 6910 1934 6918 1936
rect 6934 1940 6942 1942
rect 6934 1936 6936 1940
rect 6940 1936 6942 1940
rect 6934 1934 6942 1936
rect 6958 1940 6966 1942
rect 6958 1936 6960 1940
rect 6964 1936 6966 1940
rect 6958 1934 6966 1936
rect 6982 1940 6990 1942
rect 6982 1936 6984 1940
rect 6988 1936 6990 1940
rect 6982 1934 6990 1936
rect 7006 1940 7014 1942
rect 7006 1936 7008 1940
rect 7012 1936 7014 1940
rect 7006 1934 7014 1936
rect 7030 1940 7038 1942
rect 7030 1936 7032 1940
rect 7036 1936 7038 1940
rect 7030 1934 7038 1936
rect 7054 1940 7062 1942
rect 7054 1936 7056 1940
rect 7060 1936 7062 1940
rect 7054 1934 7062 1936
rect 7078 1940 7086 1942
rect 7078 1936 7080 1940
rect 7084 1936 7086 1940
rect 7078 1934 7086 1936
rect 7102 1940 7110 1942
rect 7102 1936 7104 1940
rect 7108 1936 7110 1940
rect 7102 1934 7110 1936
rect 7126 1940 7134 1942
rect 7126 1936 7128 1940
rect 7132 1936 7134 1940
rect 7126 1934 7134 1936
rect 7150 1940 7158 1942
rect 7150 1936 7152 1940
rect 7156 1936 7158 1940
rect 7150 1934 7158 1936
rect 7174 1940 7182 1942
rect 7174 1936 7176 1940
rect 7180 1936 7182 1940
rect 7174 1934 7182 1936
rect 7198 1934 7200 1942
rect 2410 1928 2418 1930
rect 2410 1924 2412 1928
rect 2416 1924 2418 1928
rect 2410 1922 2418 1924
rect 2434 1928 2442 1930
rect 2434 1924 2436 1928
rect 2440 1924 2442 1928
rect 2434 1922 2442 1924
rect 2458 1928 2466 1930
rect 2458 1924 2460 1928
rect 2464 1924 2466 1928
rect 2458 1922 2466 1924
rect 2482 1928 2490 1930
rect 2482 1924 2484 1928
rect 2488 1924 2490 1928
rect 2482 1922 2490 1924
rect 2698 1928 2706 1930
rect 2698 1924 2700 1928
rect 2704 1924 2706 1928
rect 2698 1922 2706 1924
rect 2722 1928 2730 1930
rect 2722 1924 2724 1928
rect 2728 1924 2730 1928
rect 2722 1922 2730 1924
rect 2746 1928 2754 1930
rect 2746 1924 2748 1928
rect 2752 1924 2754 1928
rect 2746 1922 2754 1924
rect 2770 1928 2778 1930
rect 2770 1924 2772 1928
rect 2776 1924 2778 1928
rect 2770 1922 2778 1924
rect 2794 1928 2802 1930
rect 2794 1924 2796 1928
rect 2800 1924 2802 1928
rect 2794 1922 2802 1924
rect 2818 1928 2826 1930
rect 2818 1924 2820 1928
rect 2824 1924 2826 1928
rect 2818 1922 2826 1924
rect 2842 1928 2850 1930
rect 2842 1924 2844 1928
rect 2848 1924 2850 1928
rect 2842 1922 2850 1924
rect 2866 1928 2874 1930
rect 2866 1924 2868 1928
rect 2872 1924 2874 1928
rect 2866 1922 2874 1924
rect 2890 1928 2898 1930
rect 2890 1924 2892 1928
rect 2896 1924 2898 1928
rect 2890 1922 2898 1924
rect 2914 1928 2922 1930
rect 2914 1924 2916 1928
rect 2920 1924 2922 1928
rect 2914 1922 2922 1924
rect 2938 1928 2946 1930
rect 2938 1924 2940 1928
rect 2944 1924 2946 1928
rect 2938 1922 2946 1924
rect 2962 1928 2970 1930
rect 2962 1924 2964 1928
rect 2968 1924 2970 1928
rect 2962 1922 2970 1924
rect 2986 1928 2994 1930
rect 2986 1924 2988 1928
rect 2992 1924 2994 1928
rect 2986 1922 2994 1924
rect 3010 1928 3018 1930
rect 3010 1924 3012 1928
rect 3016 1924 3018 1928
rect 3010 1922 3018 1924
rect 3034 1928 3042 1930
rect 3034 1924 3036 1928
rect 3040 1924 3042 1928
rect 3034 1922 3042 1924
rect 3058 1928 3066 1930
rect 3058 1924 3060 1928
rect 3064 1924 3066 1928
rect 3058 1922 3066 1924
rect 3082 1928 3090 1930
rect 3082 1924 3084 1928
rect 3088 1924 3090 1928
rect 3082 1922 3090 1924
rect 3298 1928 3306 1930
rect 3298 1924 3300 1928
rect 3304 1924 3306 1928
rect 3298 1922 3306 1924
rect 3322 1928 3330 1930
rect 3322 1924 3324 1928
rect 3328 1924 3330 1928
rect 3322 1922 3330 1924
rect 3346 1928 3354 1930
rect 3346 1924 3348 1928
rect 3352 1924 3354 1928
rect 3346 1922 3354 1924
rect 3370 1928 3378 1930
rect 3370 1924 3372 1928
rect 3376 1924 3378 1928
rect 3370 1922 3378 1924
rect 3394 1928 3402 1930
rect 3394 1924 3396 1928
rect 3400 1924 3402 1928
rect 3394 1922 3402 1924
rect 3418 1928 3426 1930
rect 3418 1924 3420 1928
rect 3424 1924 3426 1928
rect 3418 1922 3426 1924
rect 3442 1928 3450 1930
rect 3442 1924 3444 1928
rect 3448 1924 3450 1928
rect 3442 1922 3450 1924
rect 3466 1928 3474 1930
rect 3466 1924 3468 1928
rect 3472 1924 3474 1928
rect 3466 1922 3474 1924
rect 3490 1928 3498 1930
rect 3490 1924 3492 1928
rect 3496 1924 3498 1928
rect 3490 1922 3498 1924
rect 3514 1928 3522 1930
rect 3514 1924 3516 1928
rect 3520 1924 3522 1928
rect 3514 1922 3522 1924
rect 3538 1928 3546 1930
rect 3538 1924 3540 1928
rect 3544 1924 3546 1928
rect 3538 1922 3546 1924
rect 3562 1928 3570 1930
rect 3562 1924 3564 1928
rect 3568 1924 3570 1928
rect 3562 1922 3570 1924
rect 3586 1928 3594 1930
rect 3586 1924 3588 1928
rect 3592 1924 3594 1928
rect 3586 1922 3594 1924
rect 3610 1928 3618 1930
rect 3610 1924 3612 1928
rect 3616 1924 3618 1928
rect 3610 1922 3618 1924
rect 3634 1928 3642 1930
rect 3634 1924 3636 1928
rect 3640 1924 3642 1928
rect 3634 1922 3642 1924
rect 3658 1928 3666 1930
rect 3658 1924 3660 1928
rect 3664 1924 3666 1928
rect 3658 1922 3666 1924
rect 3682 1928 3690 1930
rect 3682 1924 3684 1928
rect 3688 1924 3690 1928
rect 3682 1922 3690 1924
rect 3898 1928 3906 1930
rect 3898 1924 3900 1928
rect 3904 1924 3906 1928
rect 3898 1922 3906 1924
rect 3922 1928 3930 1930
rect 3922 1924 3924 1928
rect 3928 1924 3930 1928
rect 3922 1922 3930 1924
rect 3946 1928 3954 1930
rect 3946 1924 3948 1928
rect 3952 1924 3954 1928
rect 3946 1922 3954 1924
rect 3970 1928 3978 1930
rect 3970 1924 3972 1928
rect 3976 1924 3978 1928
rect 3970 1922 3978 1924
rect 3994 1928 4002 1930
rect 3994 1924 3996 1928
rect 4000 1924 4002 1928
rect 3994 1922 4002 1924
rect 4018 1928 4026 1930
rect 4018 1924 4020 1928
rect 4024 1924 4026 1928
rect 4018 1922 4026 1924
rect 4042 1928 4050 1930
rect 4042 1924 4044 1928
rect 4048 1924 4050 1928
rect 4042 1922 4050 1924
rect 4066 1928 4074 1930
rect 4066 1924 4068 1928
rect 4072 1924 4074 1928
rect 4066 1922 4074 1924
rect 4090 1928 4098 1930
rect 4090 1924 4092 1928
rect 4096 1924 4098 1928
rect 4090 1922 4098 1924
rect 4114 1928 4122 1930
rect 4114 1924 4116 1928
rect 4120 1924 4122 1928
rect 4114 1922 4122 1924
rect 4138 1928 4146 1930
rect 4138 1924 4140 1928
rect 4144 1924 4146 1928
rect 4138 1922 4146 1924
rect 4162 1928 4170 1930
rect 4162 1924 4164 1928
rect 4168 1924 4170 1928
rect 4162 1922 4170 1924
rect 4186 1928 4194 1930
rect 4186 1924 4188 1928
rect 4192 1924 4194 1928
rect 4186 1922 4194 1924
rect 4210 1928 4218 1930
rect 4210 1924 4212 1928
rect 4216 1924 4218 1928
rect 4210 1922 4218 1924
rect 4234 1928 4242 1930
rect 4234 1924 4236 1928
rect 4240 1924 4242 1928
rect 4234 1922 4242 1924
rect 4258 1928 4266 1930
rect 4258 1924 4260 1928
rect 4264 1924 4266 1928
rect 4258 1922 4266 1924
rect 4282 1928 4290 1930
rect 4282 1924 4284 1928
rect 4288 1924 4290 1928
rect 4282 1922 4290 1924
rect 4498 1928 4506 1930
rect 4498 1924 4500 1928
rect 4504 1924 4506 1928
rect 4498 1922 4506 1924
rect 4522 1928 4530 1930
rect 4522 1924 4524 1928
rect 4528 1924 4530 1928
rect 4522 1922 4530 1924
rect 4546 1928 4554 1930
rect 4546 1924 4548 1928
rect 4552 1924 4554 1928
rect 4546 1922 4554 1924
rect 4570 1928 4578 1930
rect 4570 1924 4572 1928
rect 4576 1924 4578 1928
rect 4570 1922 4578 1924
rect 4594 1928 4602 1930
rect 4594 1924 4596 1928
rect 4600 1924 4602 1928
rect 4594 1922 4602 1924
rect 4618 1928 4626 1930
rect 4618 1924 4620 1928
rect 4624 1924 4626 1928
rect 4618 1922 4626 1924
rect 4642 1928 4650 1930
rect 4642 1924 4644 1928
rect 4648 1924 4650 1928
rect 4642 1922 4650 1924
rect 4666 1928 4674 1930
rect 4666 1924 4668 1928
rect 4672 1924 4674 1928
rect 4666 1922 4674 1924
rect 4690 1928 4698 1930
rect 4690 1924 4692 1928
rect 4696 1924 4698 1928
rect 4690 1922 4698 1924
rect 4714 1928 4722 1930
rect 4714 1924 4716 1928
rect 4720 1924 4722 1928
rect 4714 1922 4722 1924
rect 4738 1928 4746 1930
rect 4738 1924 4740 1928
rect 4744 1924 4746 1928
rect 4738 1922 4746 1924
rect 4762 1928 4770 1930
rect 4762 1924 4764 1928
rect 4768 1924 4770 1928
rect 4762 1922 4770 1924
rect 4786 1928 4794 1930
rect 4786 1924 4788 1928
rect 4792 1924 4794 1928
rect 4786 1922 4794 1924
rect 5698 1928 5706 1930
rect 5698 1924 5700 1928
rect 5704 1924 5706 1928
rect 5698 1922 5706 1924
rect 5722 1928 5730 1930
rect 5722 1924 5724 1928
rect 5728 1924 5730 1928
rect 5722 1922 5730 1924
rect 5746 1928 5754 1930
rect 5746 1924 5748 1928
rect 5752 1924 5754 1928
rect 5746 1922 5754 1924
rect 5770 1928 5778 1930
rect 5770 1924 5772 1928
rect 5776 1924 5778 1928
rect 5770 1922 5778 1924
rect 5794 1928 5802 1930
rect 5794 1924 5796 1928
rect 5800 1924 5802 1928
rect 5794 1922 5802 1924
rect 5818 1928 5826 1930
rect 5818 1924 5820 1928
rect 5824 1924 5826 1928
rect 5818 1922 5826 1924
rect 5842 1928 5850 1930
rect 5842 1924 5844 1928
rect 5848 1924 5850 1928
rect 5842 1922 5850 1924
rect 5866 1928 5874 1930
rect 5866 1924 5868 1928
rect 5872 1924 5874 1928
rect 5866 1922 5874 1924
rect 5890 1928 5898 1930
rect 5890 1924 5892 1928
rect 5896 1924 5898 1928
rect 5890 1922 5898 1924
rect 5914 1928 5922 1930
rect 5914 1924 5916 1928
rect 5920 1924 5922 1928
rect 5914 1922 5922 1924
rect 5938 1928 5946 1930
rect 5938 1924 5940 1928
rect 5944 1924 5946 1928
rect 5938 1922 5946 1924
rect 5962 1928 5970 1930
rect 5962 1924 5964 1928
rect 5968 1924 5970 1928
rect 5962 1922 5970 1924
rect 5986 1928 5994 1930
rect 5986 1924 5988 1928
rect 5992 1924 5994 1928
rect 5986 1922 5994 1924
rect 6010 1928 6018 1930
rect 6010 1924 6012 1928
rect 6016 1924 6018 1928
rect 6010 1922 6018 1924
rect 6034 1928 6042 1930
rect 6034 1924 6036 1928
rect 6040 1924 6042 1928
rect 6034 1922 6042 1924
rect 6058 1928 6066 1930
rect 6058 1924 6060 1928
rect 6064 1924 6066 1928
rect 6058 1922 6066 1924
rect 6082 1928 6090 1930
rect 6082 1924 6084 1928
rect 6088 1924 6090 1928
rect 6082 1922 6090 1924
rect 6298 1928 6306 1930
rect 6298 1924 6300 1928
rect 6304 1924 6306 1928
rect 6298 1922 6306 1924
rect 6322 1928 6330 1930
rect 6322 1924 6324 1928
rect 6328 1924 6330 1928
rect 6322 1922 6330 1924
rect 6346 1928 6354 1930
rect 6346 1924 6348 1928
rect 6352 1924 6354 1928
rect 6346 1922 6354 1924
rect 6370 1928 6378 1930
rect 6370 1924 6372 1928
rect 6376 1924 6378 1928
rect 6370 1922 6378 1924
rect 6394 1928 6402 1930
rect 6394 1924 6396 1928
rect 6400 1924 6402 1928
rect 6394 1922 6402 1924
rect 6418 1928 6426 1930
rect 6418 1924 6420 1928
rect 6424 1924 6426 1928
rect 6418 1922 6426 1924
rect 6442 1928 6450 1930
rect 6442 1924 6444 1928
rect 6448 1924 6450 1928
rect 6442 1922 6450 1924
rect 6466 1928 6474 1930
rect 6466 1924 6468 1928
rect 6472 1924 6474 1928
rect 6466 1922 6474 1924
rect 6490 1928 6498 1930
rect 6490 1924 6492 1928
rect 6496 1924 6498 1928
rect 6490 1922 6498 1924
rect 6514 1928 6522 1930
rect 6514 1924 6516 1928
rect 6520 1924 6522 1928
rect 6514 1922 6522 1924
rect 6538 1928 6546 1930
rect 6538 1924 6540 1928
rect 6544 1924 6546 1928
rect 6538 1922 6546 1924
rect 6562 1928 6570 1930
rect 6562 1924 6564 1928
rect 6568 1924 6570 1928
rect 6562 1922 6570 1924
rect 6586 1928 6594 1930
rect 6586 1924 6588 1928
rect 6592 1924 6594 1928
rect 6586 1922 6594 1924
rect 6610 1928 6618 1930
rect 6610 1924 6612 1928
rect 6616 1924 6618 1928
rect 6610 1922 6618 1924
rect 6634 1928 6642 1930
rect 6634 1924 6636 1928
rect 6640 1924 6642 1928
rect 6634 1922 6642 1924
rect 6658 1928 6666 1930
rect 6658 1924 6660 1928
rect 6664 1924 6666 1928
rect 6658 1922 6666 1924
rect 6682 1928 6690 1930
rect 6682 1924 6684 1928
rect 6688 1924 6690 1928
rect 6682 1922 6690 1924
rect 6898 1928 6906 1930
rect 6898 1924 6900 1928
rect 6904 1924 6906 1928
rect 6898 1922 6906 1924
rect 6922 1928 6930 1930
rect 6922 1924 6924 1928
rect 6928 1924 6930 1928
rect 6922 1922 6930 1924
rect 6946 1928 6954 1930
rect 6946 1924 6948 1928
rect 6952 1924 6954 1928
rect 6946 1922 6954 1924
rect 6970 1928 6978 1930
rect 6970 1924 6972 1928
rect 6976 1924 6978 1928
rect 6970 1922 6978 1924
rect 6994 1928 7002 1930
rect 6994 1924 6996 1928
rect 7000 1924 7002 1928
rect 6994 1922 7002 1924
rect 7018 1928 7026 1930
rect 7018 1924 7020 1928
rect 7024 1924 7026 1928
rect 7018 1922 7026 1924
rect 7042 1928 7050 1930
rect 7042 1924 7044 1928
rect 7048 1924 7050 1928
rect 7042 1922 7050 1924
rect 7066 1928 7074 1930
rect 7066 1924 7068 1928
rect 7072 1924 7074 1928
rect 7066 1922 7074 1924
rect 7090 1928 7098 1930
rect 7090 1924 7092 1928
rect 7096 1924 7098 1928
rect 7090 1922 7098 1924
rect 7114 1928 7122 1930
rect 7114 1924 7116 1928
rect 7120 1924 7122 1928
rect 7114 1922 7122 1924
rect 7138 1928 7146 1930
rect 7138 1924 7140 1928
rect 7144 1924 7146 1928
rect 7138 1922 7146 1924
rect 7162 1928 7170 1930
rect 7162 1924 7164 1928
rect 7168 1924 7170 1928
rect 7162 1922 7170 1924
rect 7186 1928 7194 1930
rect 7186 1924 7188 1928
rect 7192 1924 7194 1928
rect 7186 1922 7194 1924
rect 2400 1916 2406 1918
rect 2404 1912 2406 1916
rect 2400 1910 2406 1912
rect 2422 1916 2430 1918
rect 2422 1912 2424 1916
rect 2428 1912 2430 1916
rect 2422 1910 2430 1912
rect 2446 1916 2454 1918
rect 2446 1912 2448 1916
rect 2452 1912 2454 1916
rect 2446 1910 2454 1912
rect 2470 1916 2478 1918
rect 2470 1912 2472 1916
rect 2476 1912 2478 1916
rect 2470 1910 2478 1912
rect 2494 1916 2502 1918
rect 2494 1912 2496 1916
rect 2500 1912 2502 1916
rect 2494 1910 2502 1912
rect 2710 1916 2718 1918
rect 2710 1912 2712 1916
rect 2716 1912 2718 1916
rect 2710 1910 2718 1912
rect 2734 1916 2742 1918
rect 2734 1912 2736 1916
rect 2740 1912 2742 1916
rect 2734 1910 2742 1912
rect 2758 1916 2766 1918
rect 2758 1912 2760 1916
rect 2764 1912 2766 1916
rect 2758 1910 2766 1912
rect 2782 1916 2790 1918
rect 2782 1912 2784 1916
rect 2788 1912 2790 1916
rect 2782 1910 2790 1912
rect 2806 1916 2814 1918
rect 2806 1912 2808 1916
rect 2812 1912 2814 1916
rect 2806 1910 2814 1912
rect 2830 1916 2838 1918
rect 2830 1912 2832 1916
rect 2836 1912 2838 1916
rect 2830 1910 2838 1912
rect 2854 1916 2862 1918
rect 2854 1912 2856 1916
rect 2860 1912 2862 1916
rect 2854 1910 2862 1912
rect 2878 1916 2886 1918
rect 2878 1912 2880 1916
rect 2884 1912 2886 1916
rect 2878 1910 2886 1912
rect 2902 1916 2910 1918
rect 2902 1912 2904 1916
rect 2908 1912 2910 1916
rect 2902 1910 2910 1912
rect 2926 1916 2934 1918
rect 2926 1912 2928 1916
rect 2932 1912 2934 1916
rect 2926 1910 2934 1912
rect 2950 1916 2958 1918
rect 2950 1912 2952 1916
rect 2956 1912 2958 1916
rect 2950 1910 2958 1912
rect 2974 1916 2982 1918
rect 2974 1912 2976 1916
rect 2980 1912 2982 1916
rect 2974 1910 2982 1912
rect 2998 1916 3006 1918
rect 2998 1912 3000 1916
rect 3004 1912 3006 1916
rect 2998 1910 3006 1912
rect 3022 1916 3030 1918
rect 3022 1912 3024 1916
rect 3028 1912 3030 1916
rect 3022 1910 3030 1912
rect 3046 1916 3054 1918
rect 3046 1912 3048 1916
rect 3052 1912 3054 1916
rect 3046 1910 3054 1912
rect 3070 1916 3078 1918
rect 3070 1912 3072 1916
rect 3076 1912 3078 1916
rect 3070 1910 3078 1912
rect 3094 1916 3102 1918
rect 3094 1912 3096 1916
rect 3100 1912 3102 1916
rect 3094 1910 3102 1912
rect 3310 1916 3318 1918
rect 3310 1912 3312 1916
rect 3316 1912 3318 1916
rect 3310 1910 3318 1912
rect 3334 1916 3342 1918
rect 3334 1912 3336 1916
rect 3340 1912 3342 1916
rect 3334 1910 3342 1912
rect 3358 1916 3366 1918
rect 3358 1912 3360 1916
rect 3364 1912 3366 1916
rect 3358 1910 3366 1912
rect 3382 1916 3390 1918
rect 3382 1912 3384 1916
rect 3388 1912 3390 1916
rect 3382 1910 3390 1912
rect 3406 1916 3414 1918
rect 3406 1912 3408 1916
rect 3412 1912 3414 1916
rect 3406 1910 3414 1912
rect 3430 1916 3438 1918
rect 3430 1912 3432 1916
rect 3436 1912 3438 1916
rect 3430 1910 3438 1912
rect 3454 1916 3462 1918
rect 3454 1912 3456 1916
rect 3460 1912 3462 1916
rect 3454 1910 3462 1912
rect 3478 1916 3486 1918
rect 3478 1912 3480 1916
rect 3484 1912 3486 1916
rect 3478 1910 3486 1912
rect 3502 1916 3510 1918
rect 3502 1912 3504 1916
rect 3508 1912 3510 1916
rect 3502 1910 3510 1912
rect 3526 1916 3534 1918
rect 3526 1912 3528 1916
rect 3532 1912 3534 1916
rect 3526 1910 3534 1912
rect 3550 1916 3558 1918
rect 3550 1912 3552 1916
rect 3556 1912 3558 1916
rect 3550 1910 3558 1912
rect 3574 1916 3582 1918
rect 3574 1912 3576 1916
rect 3580 1912 3582 1916
rect 3574 1910 3582 1912
rect 3598 1916 3606 1918
rect 3598 1912 3600 1916
rect 3604 1912 3606 1916
rect 3598 1910 3606 1912
rect 3622 1916 3630 1918
rect 3622 1912 3624 1916
rect 3628 1912 3630 1916
rect 3622 1910 3630 1912
rect 3646 1916 3654 1918
rect 3646 1912 3648 1916
rect 3652 1912 3654 1916
rect 3646 1910 3654 1912
rect 3670 1916 3678 1918
rect 3670 1912 3672 1916
rect 3676 1912 3678 1916
rect 3670 1910 3678 1912
rect 3694 1916 3702 1918
rect 3694 1912 3696 1916
rect 3700 1912 3702 1916
rect 3694 1910 3702 1912
rect 3910 1916 3918 1918
rect 3910 1912 3912 1916
rect 3916 1912 3918 1916
rect 3910 1910 3918 1912
rect 3934 1916 3942 1918
rect 3934 1912 3936 1916
rect 3940 1912 3942 1916
rect 3934 1910 3942 1912
rect 3958 1916 3966 1918
rect 3958 1912 3960 1916
rect 3964 1912 3966 1916
rect 3958 1910 3966 1912
rect 3982 1916 3990 1918
rect 3982 1912 3984 1916
rect 3988 1912 3990 1916
rect 3982 1910 3990 1912
rect 4006 1916 4014 1918
rect 4006 1912 4008 1916
rect 4012 1912 4014 1916
rect 4006 1910 4014 1912
rect 4030 1916 4038 1918
rect 4030 1912 4032 1916
rect 4036 1912 4038 1916
rect 4030 1910 4038 1912
rect 4054 1916 4062 1918
rect 4054 1912 4056 1916
rect 4060 1912 4062 1916
rect 4054 1910 4062 1912
rect 4078 1916 4086 1918
rect 4078 1912 4080 1916
rect 4084 1912 4086 1916
rect 4078 1910 4086 1912
rect 4102 1916 4110 1918
rect 4102 1912 4104 1916
rect 4108 1912 4110 1916
rect 4102 1910 4110 1912
rect 4126 1916 4134 1918
rect 4126 1912 4128 1916
rect 4132 1912 4134 1916
rect 4126 1910 4134 1912
rect 4150 1916 4158 1918
rect 4150 1912 4152 1916
rect 4156 1912 4158 1916
rect 4150 1910 4158 1912
rect 4174 1916 4182 1918
rect 4174 1912 4176 1916
rect 4180 1912 4182 1916
rect 4174 1910 4182 1912
rect 4198 1916 4206 1918
rect 4198 1912 4200 1916
rect 4204 1912 4206 1916
rect 4198 1910 4206 1912
rect 4222 1916 4230 1918
rect 4222 1912 4224 1916
rect 4228 1912 4230 1916
rect 4222 1910 4230 1912
rect 4246 1916 4254 1918
rect 4246 1912 4248 1916
rect 4252 1912 4254 1916
rect 4246 1910 4254 1912
rect 4270 1916 4278 1918
rect 4270 1912 4272 1916
rect 4276 1912 4278 1916
rect 4270 1910 4278 1912
rect 4294 1916 4302 1918
rect 4294 1912 4296 1916
rect 4300 1912 4302 1916
rect 4294 1910 4302 1912
rect 4510 1916 4518 1918
rect 4510 1912 4512 1916
rect 4516 1912 4518 1916
rect 4510 1910 4518 1912
rect 4534 1916 4542 1918
rect 4534 1912 4536 1916
rect 4540 1912 4542 1916
rect 4534 1910 4542 1912
rect 4558 1916 4566 1918
rect 4558 1912 4560 1916
rect 4564 1912 4566 1916
rect 4558 1910 4566 1912
rect 4582 1916 4590 1918
rect 4582 1912 4584 1916
rect 4588 1912 4590 1916
rect 4582 1910 4590 1912
rect 4606 1916 4614 1918
rect 4606 1912 4608 1916
rect 4612 1912 4614 1916
rect 4606 1910 4614 1912
rect 4630 1916 4638 1918
rect 4630 1912 4632 1916
rect 4636 1912 4638 1916
rect 4630 1910 4638 1912
rect 4654 1916 4662 1918
rect 4654 1912 4656 1916
rect 4660 1912 4662 1916
rect 4654 1910 4662 1912
rect 4678 1916 4686 1918
rect 4678 1912 4680 1916
rect 4684 1912 4686 1916
rect 4678 1910 4686 1912
rect 4702 1916 4710 1918
rect 4702 1912 4704 1916
rect 4708 1912 4710 1916
rect 4702 1910 4710 1912
rect 4726 1916 4734 1918
rect 4726 1912 4728 1916
rect 4732 1912 4734 1916
rect 4726 1910 4734 1912
rect 4750 1916 4758 1918
rect 4750 1912 4752 1916
rect 4756 1912 4758 1916
rect 4750 1910 4758 1912
rect 4774 1916 4782 1918
rect 4774 1912 4776 1916
rect 4780 1912 4782 1916
rect 4774 1910 4782 1912
rect 4798 1910 4800 1918
rect 5710 1916 5718 1918
rect 5710 1912 5712 1916
rect 5716 1912 5718 1916
rect 5710 1910 5718 1912
rect 5734 1916 5742 1918
rect 5734 1912 5736 1916
rect 5740 1912 5742 1916
rect 5734 1910 5742 1912
rect 5758 1916 5766 1918
rect 5758 1912 5760 1916
rect 5764 1912 5766 1916
rect 5758 1910 5766 1912
rect 5782 1916 5790 1918
rect 5782 1912 5784 1916
rect 5788 1912 5790 1916
rect 5782 1910 5790 1912
rect 5806 1916 5814 1918
rect 5806 1912 5808 1916
rect 5812 1912 5814 1916
rect 5806 1910 5814 1912
rect 5830 1916 5838 1918
rect 5830 1912 5832 1916
rect 5836 1912 5838 1916
rect 5830 1910 5838 1912
rect 5854 1916 5862 1918
rect 5854 1912 5856 1916
rect 5860 1912 5862 1916
rect 5854 1910 5862 1912
rect 5878 1916 5886 1918
rect 5878 1912 5880 1916
rect 5884 1912 5886 1916
rect 5878 1910 5886 1912
rect 5902 1916 5910 1918
rect 5902 1912 5904 1916
rect 5908 1912 5910 1916
rect 5902 1910 5910 1912
rect 5926 1916 5934 1918
rect 5926 1912 5928 1916
rect 5932 1912 5934 1916
rect 5926 1910 5934 1912
rect 5950 1916 5958 1918
rect 5950 1912 5952 1916
rect 5956 1912 5958 1916
rect 5950 1910 5958 1912
rect 5974 1916 5982 1918
rect 5974 1912 5976 1916
rect 5980 1912 5982 1916
rect 5974 1910 5982 1912
rect 5998 1916 6006 1918
rect 5998 1912 6000 1916
rect 6004 1912 6006 1916
rect 5998 1910 6006 1912
rect 6022 1916 6030 1918
rect 6022 1912 6024 1916
rect 6028 1912 6030 1916
rect 6022 1910 6030 1912
rect 6046 1916 6054 1918
rect 6046 1912 6048 1916
rect 6052 1912 6054 1916
rect 6046 1910 6054 1912
rect 6070 1916 6078 1918
rect 6070 1912 6072 1916
rect 6076 1912 6078 1916
rect 6070 1910 6078 1912
rect 6094 1916 6102 1918
rect 6094 1912 6096 1916
rect 6100 1912 6102 1916
rect 6094 1910 6102 1912
rect 6310 1916 6318 1918
rect 6310 1912 6312 1916
rect 6316 1912 6318 1916
rect 6310 1910 6318 1912
rect 6334 1916 6342 1918
rect 6334 1912 6336 1916
rect 6340 1912 6342 1916
rect 6334 1910 6342 1912
rect 6358 1916 6366 1918
rect 6358 1912 6360 1916
rect 6364 1912 6366 1916
rect 6358 1910 6366 1912
rect 6382 1916 6390 1918
rect 6382 1912 6384 1916
rect 6388 1912 6390 1916
rect 6382 1910 6390 1912
rect 6406 1916 6414 1918
rect 6406 1912 6408 1916
rect 6412 1912 6414 1916
rect 6406 1910 6414 1912
rect 6430 1916 6438 1918
rect 6430 1912 6432 1916
rect 6436 1912 6438 1916
rect 6430 1910 6438 1912
rect 6454 1916 6462 1918
rect 6454 1912 6456 1916
rect 6460 1912 6462 1916
rect 6454 1910 6462 1912
rect 6478 1916 6486 1918
rect 6478 1912 6480 1916
rect 6484 1912 6486 1916
rect 6478 1910 6486 1912
rect 6502 1916 6510 1918
rect 6502 1912 6504 1916
rect 6508 1912 6510 1916
rect 6502 1910 6510 1912
rect 6526 1916 6534 1918
rect 6526 1912 6528 1916
rect 6532 1912 6534 1916
rect 6526 1910 6534 1912
rect 6550 1916 6558 1918
rect 6550 1912 6552 1916
rect 6556 1912 6558 1916
rect 6550 1910 6558 1912
rect 6574 1916 6582 1918
rect 6574 1912 6576 1916
rect 6580 1912 6582 1916
rect 6574 1910 6582 1912
rect 6598 1916 6606 1918
rect 6598 1912 6600 1916
rect 6604 1912 6606 1916
rect 6598 1910 6606 1912
rect 6622 1916 6630 1918
rect 6622 1912 6624 1916
rect 6628 1912 6630 1916
rect 6622 1910 6630 1912
rect 6646 1916 6654 1918
rect 6646 1912 6648 1916
rect 6652 1912 6654 1916
rect 6646 1910 6654 1912
rect 6670 1916 6678 1918
rect 6670 1912 6672 1916
rect 6676 1912 6678 1916
rect 6670 1910 6678 1912
rect 6694 1916 6702 1918
rect 6694 1912 6696 1916
rect 6700 1912 6702 1916
rect 6694 1910 6702 1912
rect 6910 1916 6918 1918
rect 6910 1912 6912 1916
rect 6916 1912 6918 1916
rect 6910 1910 6918 1912
rect 6934 1916 6942 1918
rect 6934 1912 6936 1916
rect 6940 1912 6942 1916
rect 6934 1910 6942 1912
rect 6958 1916 6966 1918
rect 6958 1912 6960 1916
rect 6964 1912 6966 1916
rect 6958 1910 6966 1912
rect 6982 1916 6990 1918
rect 6982 1912 6984 1916
rect 6988 1912 6990 1916
rect 6982 1910 6990 1912
rect 7006 1916 7014 1918
rect 7006 1912 7008 1916
rect 7012 1912 7014 1916
rect 7006 1910 7014 1912
rect 7030 1916 7038 1918
rect 7030 1912 7032 1916
rect 7036 1912 7038 1916
rect 7030 1910 7038 1912
rect 7054 1916 7062 1918
rect 7054 1912 7056 1916
rect 7060 1912 7062 1916
rect 7054 1910 7062 1912
rect 7078 1916 7086 1918
rect 7078 1912 7080 1916
rect 7084 1912 7086 1916
rect 7078 1910 7086 1912
rect 7102 1916 7110 1918
rect 7102 1912 7104 1916
rect 7108 1912 7110 1916
rect 7102 1910 7110 1912
rect 7126 1916 7134 1918
rect 7126 1912 7128 1916
rect 7132 1912 7134 1916
rect 7126 1910 7134 1912
rect 7150 1916 7158 1918
rect 7150 1912 7152 1916
rect 7156 1912 7158 1916
rect 7150 1910 7158 1912
rect 7174 1916 7182 1918
rect 7174 1912 7176 1916
rect 7180 1912 7182 1916
rect 7174 1910 7182 1912
rect 7198 1910 7200 1918
rect 2410 1904 2418 1906
rect 2410 1900 2412 1904
rect 2416 1900 2418 1904
rect 2410 1898 2418 1900
rect 2434 1904 2442 1906
rect 2434 1900 2436 1904
rect 2440 1900 2442 1904
rect 2434 1898 2442 1900
rect 2458 1904 2466 1906
rect 2458 1900 2460 1904
rect 2464 1900 2466 1904
rect 2458 1898 2466 1900
rect 2482 1904 2490 1906
rect 2482 1900 2484 1904
rect 2488 1900 2490 1904
rect 2482 1898 2490 1900
rect 2698 1904 2706 1906
rect 2698 1900 2700 1904
rect 2704 1900 2706 1904
rect 2698 1898 2706 1900
rect 2722 1904 2730 1906
rect 2722 1900 2724 1904
rect 2728 1900 2730 1904
rect 2722 1898 2730 1900
rect 2746 1904 2754 1906
rect 2746 1900 2748 1904
rect 2752 1900 2754 1904
rect 2746 1898 2754 1900
rect 2770 1904 2778 1906
rect 2770 1900 2772 1904
rect 2776 1900 2778 1904
rect 2770 1898 2778 1900
rect 2794 1904 2802 1906
rect 2794 1900 2796 1904
rect 2800 1900 2802 1904
rect 2794 1898 2802 1900
rect 2818 1904 2826 1906
rect 2818 1900 2820 1904
rect 2824 1900 2826 1904
rect 2818 1898 2826 1900
rect 2842 1904 2850 1906
rect 2842 1900 2844 1904
rect 2848 1900 2850 1904
rect 2842 1898 2850 1900
rect 2866 1904 2874 1906
rect 2866 1900 2868 1904
rect 2872 1900 2874 1904
rect 2866 1898 2874 1900
rect 2890 1904 2898 1906
rect 2890 1900 2892 1904
rect 2896 1900 2898 1904
rect 2890 1898 2898 1900
rect 2914 1904 2922 1906
rect 2914 1900 2916 1904
rect 2920 1900 2922 1904
rect 2914 1898 2922 1900
rect 2938 1904 2946 1906
rect 2938 1900 2940 1904
rect 2944 1900 2946 1904
rect 2938 1898 2946 1900
rect 2962 1904 2970 1906
rect 2962 1900 2964 1904
rect 2968 1900 2970 1904
rect 2962 1898 2970 1900
rect 2986 1904 2994 1906
rect 2986 1900 2988 1904
rect 2992 1900 2994 1904
rect 2986 1898 2994 1900
rect 3010 1904 3018 1906
rect 3010 1900 3012 1904
rect 3016 1900 3018 1904
rect 3010 1898 3018 1900
rect 3034 1904 3042 1906
rect 3034 1900 3036 1904
rect 3040 1900 3042 1904
rect 3034 1898 3042 1900
rect 3058 1904 3066 1906
rect 3058 1900 3060 1904
rect 3064 1900 3066 1904
rect 3058 1898 3066 1900
rect 3082 1904 3090 1906
rect 3082 1900 3084 1904
rect 3088 1900 3090 1904
rect 3082 1898 3090 1900
rect 3298 1904 3306 1906
rect 3298 1900 3300 1904
rect 3304 1900 3306 1904
rect 3298 1898 3306 1900
rect 3322 1904 3330 1906
rect 3322 1900 3324 1904
rect 3328 1900 3330 1904
rect 3322 1898 3330 1900
rect 3346 1904 3354 1906
rect 3346 1900 3348 1904
rect 3352 1900 3354 1904
rect 3346 1898 3354 1900
rect 3370 1904 3378 1906
rect 3370 1900 3372 1904
rect 3376 1900 3378 1904
rect 3370 1898 3378 1900
rect 3394 1904 3402 1906
rect 3394 1900 3396 1904
rect 3400 1900 3402 1904
rect 3394 1898 3402 1900
rect 3418 1904 3426 1906
rect 3418 1900 3420 1904
rect 3424 1900 3426 1904
rect 3418 1898 3426 1900
rect 3442 1904 3450 1906
rect 3442 1900 3444 1904
rect 3448 1900 3450 1904
rect 3442 1898 3450 1900
rect 3466 1904 3474 1906
rect 3466 1900 3468 1904
rect 3472 1900 3474 1904
rect 3466 1898 3474 1900
rect 3490 1904 3498 1906
rect 3490 1900 3492 1904
rect 3496 1900 3498 1904
rect 3490 1898 3498 1900
rect 3514 1904 3522 1906
rect 3514 1900 3516 1904
rect 3520 1900 3522 1904
rect 3514 1898 3522 1900
rect 3538 1904 3546 1906
rect 3538 1900 3540 1904
rect 3544 1900 3546 1904
rect 3538 1898 3546 1900
rect 3562 1904 3570 1906
rect 3562 1900 3564 1904
rect 3568 1900 3570 1904
rect 3562 1898 3570 1900
rect 3586 1904 3594 1906
rect 3586 1900 3588 1904
rect 3592 1900 3594 1904
rect 3586 1898 3594 1900
rect 3610 1904 3618 1906
rect 3610 1900 3612 1904
rect 3616 1900 3618 1904
rect 3610 1898 3618 1900
rect 3634 1904 3642 1906
rect 3634 1900 3636 1904
rect 3640 1900 3642 1904
rect 3634 1898 3642 1900
rect 3658 1904 3666 1906
rect 3658 1900 3660 1904
rect 3664 1900 3666 1904
rect 3658 1898 3666 1900
rect 3682 1904 3690 1906
rect 3682 1900 3684 1904
rect 3688 1900 3690 1904
rect 3682 1898 3690 1900
rect 3898 1904 3906 1906
rect 3898 1900 3900 1904
rect 3904 1900 3906 1904
rect 3898 1898 3906 1900
rect 3922 1904 3930 1906
rect 3922 1900 3924 1904
rect 3928 1900 3930 1904
rect 3922 1898 3930 1900
rect 3946 1904 3954 1906
rect 3946 1900 3948 1904
rect 3952 1900 3954 1904
rect 3946 1898 3954 1900
rect 3970 1904 3978 1906
rect 3970 1900 3972 1904
rect 3976 1900 3978 1904
rect 3970 1898 3978 1900
rect 3994 1904 4002 1906
rect 3994 1900 3996 1904
rect 4000 1900 4002 1904
rect 3994 1898 4002 1900
rect 4018 1904 4026 1906
rect 4018 1900 4020 1904
rect 4024 1900 4026 1904
rect 4018 1898 4026 1900
rect 4042 1904 4050 1906
rect 4042 1900 4044 1904
rect 4048 1900 4050 1904
rect 4042 1898 4050 1900
rect 4066 1904 4074 1906
rect 4066 1900 4068 1904
rect 4072 1900 4074 1904
rect 4066 1898 4074 1900
rect 4090 1904 4098 1906
rect 4090 1900 4092 1904
rect 4096 1900 4098 1904
rect 4090 1898 4098 1900
rect 4114 1904 4122 1906
rect 4114 1900 4116 1904
rect 4120 1900 4122 1904
rect 4114 1898 4122 1900
rect 4138 1904 4146 1906
rect 4138 1900 4140 1904
rect 4144 1900 4146 1904
rect 4138 1898 4146 1900
rect 4162 1904 4170 1906
rect 4162 1900 4164 1904
rect 4168 1900 4170 1904
rect 4162 1898 4170 1900
rect 4186 1904 4194 1906
rect 4186 1900 4188 1904
rect 4192 1900 4194 1904
rect 4186 1898 4194 1900
rect 4210 1904 4218 1906
rect 4210 1900 4212 1904
rect 4216 1900 4218 1904
rect 4210 1898 4218 1900
rect 4234 1904 4242 1906
rect 4234 1900 4236 1904
rect 4240 1900 4242 1904
rect 4234 1898 4242 1900
rect 4258 1904 4266 1906
rect 4258 1900 4260 1904
rect 4264 1900 4266 1904
rect 4258 1898 4266 1900
rect 4282 1904 4290 1906
rect 4282 1900 4284 1904
rect 4288 1900 4290 1904
rect 4282 1898 4290 1900
rect 4498 1904 4506 1906
rect 4498 1900 4500 1904
rect 4504 1900 4506 1904
rect 4498 1898 4506 1900
rect 4522 1904 4530 1906
rect 4522 1900 4524 1904
rect 4528 1900 4530 1904
rect 4522 1898 4530 1900
rect 4546 1904 4554 1906
rect 4546 1900 4548 1904
rect 4552 1900 4554 1904
rect 4546 1898 4554 1900
rect 4570 1904 4578 1906
rect 4570 1900 4572 1904
rect 4576 1900 4578 1904
rect 4570 1898 4578 1900
rect 4594 1904 4602 1906
rect 4594 1900 4596 1904
rect 4600 1900 4602 1904
rect 4594 1898 4602 1900
rect 4618 1904 4626 1906
rect 4618 1900 4620 1904
rect 4624 1900 4626 1904
rect 4618 1898 4626 1900
rect 4642 1904 4650 1906
rect 4642 1900 4644 1904
rect 4648 1900 4650 1904
rect 4642 1898 4650 1900
rect 4666 1904 4674 1906
rect 4666 1900 4668 1904
rect 4672 1900 4674 1904
rect 4666 1898 4674 1900
rect 4690 1904 4698 1906
rect 4690 1900 4692 1904
rect 4696 1900 4698 1904
rect 4690 1898 4698 1900
rect 4714 1904 4722 1906
rect 4714 1900 4716 1904
rect 4720 1900 4722 1904
rect 4714 1898 4722 1900
rect 4738 1904 4746 1906
rect 4738 1900 4740 1904
rect 4744 1900 4746 1904
rect 4738 1898 4746 1900
rect 4762 1904 4770 1906
rect 4762 1900 4764 1904
rect 4768 1900 4770 1904
rect 4762 1898 4770 1900
rect 4786 1904 4794 1906
rect 4786 1900 4788 1904
rect 4792 1900 4794 1904
rect 4786 1898 4794 1900
rect 5698 1904 5706 1906
rect 5698 1900 5700 1904
rect 5704 1900 5706 1904
rect 5698 1898 5706 1900
rect 5722 1904 5730 1906
rect 5722 1900 5724 1904
rect 5728 1900 5730 1904
rect 5722 1898 5730 1900
rect 5746 1904 5754 1906
rect 5746 1900 5748 1904
rect 5752 1900 5754 1904
rect 5746 1898 5754 1900
rect 5770 1904 5778 1906
rect 5770 1900 5772 1904
rect 5776 1900 5778 1904
rect 5770 1898 5778 1900
rect 5794 1904 5802 1906
rect 5794 1900 5796 1904
rect 5800 1900 5802 1904
rect 5794 1898 5802 1900
rect 5818 1904 5826 1906
rect 5818 1900 5820 1904
rect 5824 1900 5826 1904
rect 5818 1898 5826 1900
rect 5842 1904 5850 1906
rect 5842 1900 5844 1904
rect 5848 1900 5850 1904
rect 5842 1898 5850 1900
rect 5866 1904 5874 1906
rect 5866 1900 5868 1904
rect 5872 1900 5874 1904
rect 5866 1898 5874 1900
rect 5890 1904 5898 1906
rect 5890 1900 5892 1904
rect 5896 1900 5898 1904
rect 5890 1898 5898 1900
rect 5914 1904 5922 1906
rect 5914 1900 5916 1904
rect 5920 1900 5922 1904
rect 5914 1898 5922 1900
rect 5938 1904 5946 1906
rect 5938 1900 5940 1904
rect 5944 1900 5946 1904
rect 5938 1898 5946 1900
rect 5962 1904 5970 1906
rect 5962 1900 5964 1904
rect 5968 1900 5970 1904
rect 5962 1898 5970 1900
rect 5986 1904 5994 1906
rect 5986 1900 5988 1904
rect 5992 1900 5994 1904
rect 5986 1898 5994 1900
rect 6010 1904 6018 1906
rect 6010 1900 6012 1904
rect 6016 1900 6018 1904
rect 6010 1898 6018 1900
rect 6034 1904 6042 1906
rect 6034 1900 6036 1904
rect 6040 1900 6042 1904
rect 6034 1898 6042 1900
rect 6058 1904 6066 1906
rect 6058 1900 6060 1904
rect 6064 1900 6066 1904
rect 6058 1898 6066 1900
rect 6082 1904 6090 1906
rect 6082 1900 6084 1904
rect 6088 1900 6090 1904
rect 6082 1898 6090 1900
rect 6298 1904 6306 1906
rect 6298 1900 6300 1904
rect 6304 1900 6306 1904
rect 6298 1898 6306 1900
rect 6322 1904 6330 1906
rect 6322 1900 6324 1904
rect 6328 1900 6330 1904
rect 6322 1898 6330 1900
rect 6346 1904 6354 1906
rect 6346 1900 6348 1904
rect 6352 1900 6354 1904
rect 6346 1898 6354 1900
rect 6370 1904 6378 1906
rect 6370 1900 6372 1904
rect 6376 1900 6378 1904
rect 6370 1898 6378 1900
rect 6394 1904 6402 1906
rect 6394 1900 6396 1904
rect 6400 1900 6402 1904
rect 6394 1898 6402 1900
rect 6418 1904 6426 1906
rect 6418 1900 6420 1904
rect 6424 1900 6426 1904
rect 6418 1898 6426 1900
rect 6442 1904 6450 1906
rect 6442 1900 6444 1904
rect 6448 1900 6450 1904
rect 6442 1898 6450 1900
rect 6466 1904 6474 1906
rect 6466 1900 6468 1904
rect 6472 1900 6474 1904
rect 6466 1898 6474 1900
rect 6490 1904 6498 1906
rect 6490 1900 6492 1904
rect 6496 1900 6498 1904
rect 6490 1898 6498 1900
rect 6514 1904 6522 1906
rect 6514 1900 6516 1904
rect 6520 1900 6522 1904
rect 6514 1898 6522 1900
rect 6538 1904 6546 1906
rect 6538 1900 6540 1904
rect 6544 1900 6546 1904
rect 6538 1898 6546 1900
rect 6562 1904 6570 1906
rect 6562 1900 6564 1904
rect 6568 1900 6570 1904
rect 6562 1898 6570 1900
rect 6586 1904 6594 1906
rect 6586 1900 6588 1904
rect 6592 1900 6594 1904
rect 6586 1898 6594 1900
rect 6610 1904 6618 1906
rect 6610 1900 6612 1904
rect 6616 1900 6618 1904
rect 6610 1898 6618 1900
rect 6634 1904 6642 1906
rect 6634 1900 6636 1904
rect 6640 1900 6642 1904
rect 6634 1898 6642 1900
rect 6658 1904 6666 1906
rect 6658 1900 6660 1904
rect 6664 1900 6666 1904
rect 6658 1898 6666 1900
rect 6682 1904 6690 1906
rect 6682 1900 6684 1904
rect 6688 1900 6690 1904
rect 6682 1898 6690 1900
rect 6898 1904 6906 1906
rect 6898 1900 6900 1904
rect 6904 1900 6906 1904
rect 6898 1898 6906 1900
rect 6922 1904 6930 1906
rect 6922 1900 6924 1904
rect 6928 1900 6930 1904
rect 6922 1898 6930 1900
rect 6946 1904 6954 1906
rect 6946 1900 6948 1904
rect 6952 1900 6954 1904
rect 6946 1898 6954 1900
rect 6970 1904 6978 1906
rect 6970 1900 6972 1904
rect 6976 1900 6978 1904
rect 6970 1898 6978 1900
rect 6994 1904 7002 1906
rect 6994 1900 6996 1904
rect 7000 1900 7002 1904
rect 6994 1898 7002 1900
rect 7018 1904 7026 1906
rect 7018 1900 7020 1904
rect 7024 1900 7026 1904
rect 7018 1898 7026 1900
rect 7042 1904 7050 1906
rect 7042 1900 7044 1904
rect 7048 1900 7050 1904
rect 7042 1898 7050 1900
rect 7066 1904 7074 1906
rect 7066 1900 7068 1904
rect 7072 1900 7074 1904
rect 7066 1898 7074 1900
rect 7090 1904 7098 1906
rect 7090 1900 7092 1904
rect 7096 1900 7098 1904
rect 7090 1898 7098 1900
rect 7114 1904 7122 1906
rect 7114 1900 7116 1904
rect 7120 1900 7122 1904
rect 7114 1898 7122 1900
rect 7138 1904 7146 1906
rect 7138 1900 7140 1904
rect 7144 1900 7146 1904
rect 7138 1898 7146 1900
rect 7162 1904 7170 1906
rect 7162 1900 7164 1904
rect 7168 1900 7170 1904
rect 7162 1898 7170 1900
rect 7186 1904 7194 1906
rect 7186 1900 7188 1904
rect 7192 1900 7194 1904
rect 7186 1898 7194 1900
rect 2400 1892 2406 1894
rect 2404 1888 2406 1892
rect 2400 1886 2406 1888
rect 2422 1892 2430 1894
rect 2422 1888 2424 1892
rect 2428 1888 2430 1892
rect 2422 1886 2430 1888
rect 2446 1892 2454 1894
rect 2446 1888 2448 1892
rect 2452 1888 2454 1892
rect 2446 1886 2454 1888
rect 2470 1892 2478 1894
rect 2470 1888 2472 1892
rect 2476 1888 2478 1892
rect 2470 1886 2478 1888
rect 2494 1892 2502 1894
rect 2494 1888 2496 1892
rect 2500 1888 2502 1892
rect 2494 1886 2502 1888
rect 2710 1892 2718 1894
rect 2710 1888 2712 1892
rect 2716 1888 2718 1892
rect 2710 1886 2718 1888
rect 2734 1892 2742 1894
rect 2734 1888 2736 1892
rect 2740 1888 2742 1892
rect 2734 1886 2742 1888
rect 2758 1892 2766 1894
rect 2758 1888 2760 1892
rect 2764 1888 2766 1892
rect 2758 1886 2766 1888
rect 2782 1892 2790 1894
rect 2782 1888 2784 1892
rect 2788 1888 2790 1892
rect 2782 1886 2790 1888
rect 2806 1892 2814 1894
rect 2806 1888 2808 1892
rect 2812 1888 2814 1892
rect 2806 1886 2814 1888
rect 2830 1892 2838 1894
rect 2830 1888 2832 1892
rect 2836 1888 2838 1892
rect 2830 1886 2838 1888
rect 2854 1892 2862 1894
rect 2854 1888 2856 1892
rect 2860 1888 2862 1892
rect 2854 1886 2862 1888
rect 2878 1892 2886 1894
rect 2878 1888 2880 1892
rect 2884 1888 2886 1892
rect 2878 1886 2886 1888
rect 2902 1892 2910 1894
rect 2902 1888 2904 1892
rect 2908 1888 2910 1892
rect 2902 1886 2910 1888
rect 2926 1892 2934 1894
rect 2926 1888 2928 1892
rect 2932 1888 2934 1892
rect 2926 1886 2934 1888
rect 2950 1892 2958 1894
rect 2950 1888 2952 1892
rect 2956 1888 2958 1892
rect 2950 1886 2958 1888
rect 2974 1892 2982 1894
rect 2974 1888 2976 1892
rect 2980 1888 2982 1892
rect 2974 1886 2982 1888
rect 2998 1892 3006 1894
rect 2998 1888 3000 1892
rect 3004 1888 3006 1892
rect 2998 1886 3006 1888
rect 3022 1892 3030 1894
rect 3022 1888 3024 1892
rect 3028 1888 3030 1892
rect 3022 1886 3030 1888
rect 3046 1892 3054 1894
rect 3046 1888 3048 1892
rect 3052 1888 3054 1892
rect 3046 1886 3054 1888
rect 3070 1892 3078 1894
rect 3070 1888 3072 1892
rect 3076 1888 3078 1892
rect 3070 1886 3078 1888
rect 3094 1892 3102 1894
rect 3094 1888 3096 1892
rect 3100 1888 3102 1892
rect 3094 1886 3102 1888
rect 3310 1892 3318 1894
rect 3310 1888 3312 1892
rect 3316 1888 3318 1892
rect 3310 1886 3318 1888
rect 3334 1892 3342 1894
rect 3334 1888 3336 1892
rect 3340 1888 3342 1892
rect 3334 1886 3342 1888
rect 3358 1892 3366 1894
rect 3358 1888 3360 1892
rect 3364 1888 3366 1892
rect 3358 1886 3366 1888
rect 3382 1892 3390 1894
rect 3382 1888 3384 1892
rect 3388 1888 3390 1892
rect 3382 1886 3390 1888
rect 3406 1892 3414 1894
rect 3406 1888 3408 1892
rect 3412 1888 3414 1892
rect 3406 1886 3414 1888
rect 3430 1892 3438 1894
rect 3430 1888 3432 1892
rect 3436 1888 3438 1892
rect 3430 1886 3438 1888
rect 3454 1892 3462 1894
rect 3454 1888 3456 1892
rect 3460 1888 3462 1892
rect 3454 1886 3462 1888
rect 3478 1892 3486 1894
rect 3478 1888 3480 1892
rect 3484 1888 3486 1892
rect 3478 1886 3486 1888
rect 3502 1892 3510 1894
rect 3502 1888 3504 1892
rect 3508 1888 3510 1892
rect 3502 1886 3510 1888
rect 3526 1892 3534 1894
rect 3526 1888 3528 1892
rect 3532 1888 3534 1892
rect 3526 1886 3534 1888
rect 3550 1892 3558 1894
rect 3550 1888 3552 1892
rect 3556 1888 3558 1892
rect 3550 1886 3558 1888
rect 3574 1892 3582 1894
rect 3574 1888 3576 1892
rect 3580 1888 3582 1892
rect 3574 1886 3582 1888
rect 3598 1892 3606 1894
rect 3598 1888 3600 1892
rect 3604 1888 3606 1892
rect 3598 1886 3606 1888
rect 3622 1892 3630 1894
rect 3622 1888 3624 1892
rect 3628 1888 3630 1892
rect 3622 1886 3630 1888
rect 3646 1892 3654 1894
rect 3646 1888 3648 1892
rect 3652 1888 3654 1892
rect 3646 1886 3654 1888
rect 3670 1892 3678 1894
rect 3670 1888 3672 1892
rect 3676 1888 3678 1892
rect 3670 1886 3678 1888
rect 3694 1892 3702 1894
rect 3694 1888 3696 1892
rect 3700 1888 3702 1892
rect 3694 1886 3702 1888
rect 3910 1892 3918 1894
rect 3910 1888 3912 1892
rect 3916 1888 3918 1892
rect 3910 1886 3918 1888
rect 3934 1892 3942 1894
rect 3934 1888 3936 1892
rect 3940 1888 3942 1892
rect 3934 1886 3942 1888
rect 3958 1892 3966 1894
rect 3958 1888 3960 1892
rect 3964 1888 3966 1892
rect 3958 1886 3966 1888
rect 3982 1892 3990 1894
rect 3982 1888 3984 1892
rect 3988 1888 3990 1892
rect 3982 1886 3990 1888
rect 4006 1892 4014 1894
rect 4006 1888 4008 1892
rect 4012 1888 4014 1892
rect 4006 1886 4014 1888
rect 4030 1892 4038 1894
rect 4030 1888 4032 1892
rect 4036 1888 4038 1892
rect 4030 1886 4038 1888
rect 4054 1892 4062 1894
rect 4054 1888 4056 1892
rect 4060 1888 4062 1892
rect 4054 1886 4062 1888
rect 4078 1892 4086 1894
rect 4078 1888 4080 1892
rect 4084 1888 4086 1892
rect 4078 1886 4086 1888
rect 4102 1892 4110 1894
rect 4102 1888 4104 1892
rect 4108 1888 4110 1892
rect 4102 1886 4110 1888
rect 4126 1892 4134 1894
rect 4126 1888 4128 1892
rect 4132 1888 4134 1892
rect 4126 1886 4134 1888
rect 4150 1892 4158 1894
rect 4150 1888 4152 1892
rect 4156 1888 4158 1892
rect 4150 1886 4158 1888
rect 4174 1892 4182 1894
rect 4174 1888 4176 1892
rect 4180 1888 4182 1892
rect 4174 1886 4182 1888
rect 4198 1892 4206 1894
rect 4198 1888 4200 1892
rect 4204 1888 4206 1892
rect 4198 1886 4206 1888
rect 4222 1892 4230 1894
rect 4222 1888 4224 1892
rect 4228 1888 4230 1892
rect 4222 1886 4230 1888
rect 4246 1892 4254 1894
rect 4246 1888 4248 1892
rect 4252 1888 4254 1892
rect 4246 1886 4254 1888
rect 4270 1892 4278 1894
rect 4270 1888 4272 1892
rect 4276 1888 4278 1892
rect 4270 1886 4278 1888
rect 4294 1892 4302 1894
rect 4294 1888 4296 1892
rect 4300 1888 4302 1892
rect 4294 1886 4302 1888
rect 4510 1892 4518 1894
rect 4510 1888 4512 1892
rect 4516 1888 4518 1892
rect 4510 1886 4518 1888
rect 4534 1892 4542 1894
rect 4534 1888 4536 1892
rect 4540 1888 4542 1892
rect 4534 1886 4542 1888
rect 4558 1892 4566 1894
rect 4558 1888 4560 1892
rect 4564 1888 4566 1892
rect 4558 1886 4566 1888
rect 4582 1892 4590 1894
rect 4582 1888 4584 1892
rect 4588 1888 4590 1892
rect 4582 1886 4590 1888
rect 4606 1892 4614 1894
rect 4606 1888 4608 1892
rect 4612 1888 4614 1892
rect 4606 1886 4614 1888
rect 4630 1892 4638 1894
rect 4630 1888 4632 1892
rect 4636 1888 4638 1892
rect 4630 1886 4638 1888
rect 4654 1892 4662 1894
rect 4654 1888 4656 1892
rect 4660 1888 4662 1892
rect 4654 1886 4662 1888
rect 4678 1892 4686 1894
rect 4678 1888 4680 1892
rect 4684 1888 4686 1892
rect 4678 1886 4686 1888
rect 4702 1892 4710 1894
rect 4702 1888 4704 1892
rect 4708 1888 4710 1892
rect 4702 1886 4710 1888
rect 4726 1892 4734 1894
rect 4726 1888 4728 1892
rect 4732 1888 4734 1892
rect 4726 1886 4734 1888
rect 4750 1892 4758 1894
rect 4750 1888 4752 1892
rect 4756 1888 4758 1892
rect 4750 1886 4758 1888
rect 4774 1892 4782 1894
rect 4774 1888 4776 1892
rect 4780 1888 4782 1892
rect 4774 1886 4782 1888
rect 4798 1886 4800 1894
rect 5710 1892 5718 1894
rect 5710 1888 5712 1892
rect 5716 1888 5718 1892
rect 5710 1886 5718 1888
rect 5734 1892 5742 1894
rect 5734 1888 5736 1892
rect 5740 1888 5742 1892
rect 5734 1886 5742 1888
rect 5758 1892 5766 1894
rect 5758 1888 5760 1892
rect 5764 1888 5766 1892
rect 5758 1886 5766 1888
rect 5782 1892 5790 1894
rect 5782 1888 5784 1892
rect 5788 1888 5790 1892
rect 5782 1886 5790 1888
rect 5806 1892 5814 1894
rect 5806 1888 5808 1892
rect 5812 1888 5814 1892
rect 5806 1886 5814 1888
rect 5830 1892 5838 1894
rect 5830 1888 5832 1892
rect 5836 1888 5838 1892
rect 5830 1886 5838 1888
rect 5854 1892 5862 1894
rect 5854 1888 5856 1892
rect 5860 1888 5862 1892
rect 5854 1886 5862 1888
rect 5878 1892 5886 1894
rect 5878 1888 5880 1892
rect 5884 1888 5886 1892
rect 5878 1886 5886 1888
rect 5902 1892 5910 1894
rect 5902 1888 5904 1892
rect 5908 1888 5910 1892
rect 5902 1886 5910 1888
rect 5926 1892 5934 1894
rect 5926 1888 5928 1892
rect 5932 1888 5934 1892
rect 5926 1886 5934 1888
rect 5950 1892 5958 1894
rect 5950 1888 5952 1892
rect 5956 1888 5958 1892
rect 5950 1886 5958 1888
rect 5974 1892 5982 1894
rect 5974 1888 5976 1892
rect 5980 1888 5982 1892
rect 5974 1886 5982 1888
rect 5998 1892 6006 1894
rect 5998 1888 6000 1892
rect 6004 1888 6006 1892
rect 5998 1886 6006 1888
rect 6022 1892 6030 1894
rect 6022 1888 6024 1892
rect 6028 1888 6030 1892
rect 6022 1886 6030 1888
rect 6046 1892 6054 1894
rect 6046 1888 6048 1892
rect 6052 1888 6054 1892
rect 6046 1886 6054 1888
rect 6070 1892 6078 1894
rect 6070 1888 6072 1892
rect 6076 1888 6078 1892
rect 6070 1886 6078 1888
rect 6094 1892 6102 1894
rect 6094 1888 6096 1892
rect 6100 1888 6102 1892
rect 6094 1886 6102 1888
rect 6310 1892 6318 1894
rect 6310 1888 6312 1892
rect 6316 1888 6318 1892
rect 6310 1886 6318 1888
rect 6334 1892 6342 1894
rect 6334 1888 6336 1892
rect 6340 1888 6342 1892
rect 6334 1886 6342 1888
rect 6358 1892 6366 1894
rect 6358 1888 6360 1892
rect 6364 1888 6366 1892
rect 6358 1886 6366 1888
rect 6382 1892 6390 1894
rect 6382 1888 6384 1892
rect 6388 1888 6390 1892
rect 6382 1886 6390 1888
rect 6406 1892 6414 1894
rect 6406 1888 6408 1892
rect 6412 1888 6414 1892
rect 6406 1886 6414 1888
rect 6430 1892 6438 1894
rect 6430 1888 6432 1892
rect 6436 1888 6438 1892
rect 6430 1886 6438 1888
rect 6454 1892 6462 1894
rect 6454 1888 6456 1892
rect 6460 1888 6462 1892
rect 6454 1886 6462 1888
rect 6478 1892 6486 1894
rect 6478 1888 6480 1892
rect 6484 1888 6486 1892
rect 6478 1886 6486 1888
rect 6502 1892 6510 1894
rect 6502 1888 6504 1892
rect 6508 1888 6510 1892
rect 6502 1886 6510 1888
rect 6526 1892 6534 1894
rect 6526 1888 6528 1892
rect 6532 1888 6534 1892
rect 6526 1886 6534 1888
rect 6550 1892 6558 1894
rect 6550 1888 6552 1892
rect 6556 1888 6558 1892
rect 6550 1886 6558 1888
rect 6574 1892 6582 1894
rect 6574 1888 6576 1892
rect 6580 1888 6582 1892
rect 6574 1886 6582 1888
rect 6598 1892 6606 1894
rect 6598 1888 6600 1892
rect 6604 1888 6606 1892
rect 6598 1886 6606 1888
rect 6622 1892 6630 1894
rect 6622 1888 6624 1892
rect 6628 1888 6630 1892
rect 6622 1886 6630 1888
rect 6646 1892 6654 1894
rect 6646 1888 6648 1892
rect 6652 1888 6654 1892
rect 6646 1886 6654 1888
rect 6670 1892 6678 1894
rect 6670 1888 6672 1892
rect 6676 1888 6678 1892
rect 6670 1886 6678 1888
rect 6694 1892 6702 1894
rect 6694 1888 6696 1892
rect 6700 1888 6702 1892
rect 6694 1886 6702 1888
rect 6910 1892 6918 1894
rect 6910 1888 6912 1892
rect 6916 1888 6918 1892
rect 6910 1886 6918 1888
rect 6934 1892 6942 1894
rect 6934 1888 6936 1892
rect 6940 1888 6942 1892
rect 6934 1886 6942 1888
rect 6958 1892 6966 1894
rect 6958 1888 6960 1892
rect 6964 1888 6966 1892
rect 6958 1886 6966 1888
rect 6982 1892 6990 1894
rect 6982 1888 6984 1892
rect 6988 1888 6990 1892
rect 6982 1886 6990 1888
rect 7006 1892 7014 1894
rect 7006 1888 7008 1892
rect 7012 1888 7014 1892
rect 7006 1886 7014 1888
rect 7030 1892 7038 1894
rect 7030 1888 7032 1892
rect 7036 1888 7038 1892
rect 7030 1886 7038 1888
rect 7054 1892 7062 1894
rect 7054 1888 7056 1892
rect 7060 1888 7062 1892
rect 7054 1886 7062 1888
rect 7078 1892 7086 1894
rect 7078 1888 7080 1892
rect 7084 1888 7086 1892
rect 7078 1886 7086 1888
rect 7102 1892 7110 1894
rect 7102 1888 7104 1892
rect 7108 1888 7110 1892
rect 7102 1886 7110 1888
rect 7126 1892 7134 1894
rect 7126 1888 7128 1892
rect 7132 1888 7134 1892
rect 7126 1886 7134 1888
rect 7150 1892 7158 1894
rect 7150 1888 7152 1892
rect 7156 1888 7158 1892
rect 7150 1886 7158 1888
rect 7174 1892 7182 1894
rect 7174 1888 7176 1892
rect 7180 1888 7182 1892
rect 7174 1886 7182 1888
rect 7198 1886 7200 1894
rect 2410 1880 2418 1882
rect 2410 1876 2412 1880
rect 2416 1876 2418 1880
rect 2410 1874 2418 1876
rect 2434 1880 2442 1882
rect 2434 1876 2436 1880
rect 2440 1876 2442 1880
rect 2434 1874 2442 1876
rect 2458 1880 2466 1882
rect 2458 1876 2460 1880
rect 2464 1876 2466 1880
rect 2458 1874 2466 1876
rect 2482 1880 2490 1882
rect 2482 1876 2484 1880
rect 2488 1876 2490 1880
rect 2482 1874 2490 1876
rect 2698 1880 2706 1882
rect 2698 1876 2700 1880
rect 2704 1876 2706 1880
rect 2698 1874 2706 1876
rect 2722 1880 2730 1882
rect 2722 1876 2724 1880
rect 2728 1876 2730 1880
rect 2722 1874 2730 1876
rect 2746 1880 2754 1882
rect 2746 1876 2748 1880
rect 2752 1876 2754 1880
rect 2746 1874 2754 1876
rect 2770 1880 2778 1882
rect 2770 1876 2772 1880
rect 2776 1876 2778 1880
rect 2770 1874 2778 1876
rect 2794 1880 2802 1882
rect 2794 1876 2796 1880
rect 2800 1876 2802 1880
rect 2794 1874 2802 1876
rect 2818 1880 2826 1882
rect 2818 1876 2820 1880
rect 2824 1876 2826 1880
rect 2818 1874 2826 1876
rect 2842 1880 2850 1882
rect 2842 1876 2844 1880
rect 2848 1876 2850 1880
rect 2842 1874 2850 1876
rect 2866 1880 2874 1882
rect 2866 1876 2868 1880
rect 2872 1876 2874 1880
rect 2866 1874 2874 1876
rect 2890 1880 2898 1882
rect 2890 1876 2892 1880
rect 2896 1876 2898 1880
rect 2890 1874 2898 1876
rect 2914 1880 2922 1882
rect 2914 1876 2916 1880
rect 2920 1876 2922 1880
rect 2914 1874 2922 1876
rect 2938 1880 2946 1882
rect 2938 1876 2940 1880
rect 2944 1876 2946 1880
rect 2938 1874 2946 1876
rect 2962 1880 2970 1882
rect 2962 1876 2964 1880
rect 2968 1876 2970 1880
rect 2962 1874 2970 1876
rect 2986 1880 2994 1882
rect 2986 1876 2988 1880
rect 2992 1876 2994 1880
rect 2986 1874 2994 1876
rect 3010 1880 3018 1882
rect 3010 1876 3012 1880
rect 3016 1876 3018 1880
rect 3010 1874 3018 1876
rect 3034 1880 3042 1882
rect 3034 1876 3036 1880
rect 3040 1876 3042 1880
rect 3034 1874 3042 1876
rect 3058 1880 3066 1882
rect 3058 1876 3060 1880
rect 3064 1876 3066 1880
rect 3058 1874 3066 1876
rect 3082 1880 3090 1882
rect 3082 1876 3084 1880
rect 3088 1876 3090 1880
rect 3082 1874 3090 1876
rect 3298 1880 3306 1882
rect 3298 1876 3300 1880
rect 3304 1876 3306 1880
rect 3298 1874 3306 1876
rect 3322 1880 3330 1882
rect 3322 1876 3324 1880
rect 3328 1876 3330 1880
rect 3322 1874 3330 1876
rect 3346 1880 3354 1882
rect 3346 1876 3348 1880
rect 3352 1876 3354 1880
rect 3346 1874 3354 1876
rect 3370 1880 3378 1882
rect 3370 1876 3372 1880
rect 3376 1876 3378 1880
rect 3370 1874 3378 1876
rect 3394 1880 3402 1882
rect 3394 1876 3396 1880
rect 3400 1876 3402 1880
rect 3394 1874 3402 1876
rect 3418 1880 3426 1882
rect 3418 1876 3420 1880
rect 3424 1876 3426 1880
rect 3418 1874 3426 1876
rect 3442 1880 3450 1882
rect 3442 1876 3444 1880
rect 3448 1876 3450 1880
rect 3442 1874 3450 1876
rect 3466 1880 3474 1882
rect 3466 1876 3468 1880
rect 3472 1876 3474 1880
rect 3466 1874 3474 1876
rect 3490 1880 3498 1882
rect 3490 1876 3492 1880
rect 3496 1876 3498 1880
rect 3490 1874 3498 1876
rect 3514 1880 3522 1882
rect 3514 1876 3516 1880
rect 3520 1876 3522 1880
rect 3514 1874 3522 1876
rect 3538 1880 3546 1882
rect 3538 1876 3540 1880
rect 3544 1876 3546 1880
rect 3538 1874 3546 1876
rect 3562 1880 3570 1882
rect 3562 1876 3564 1880
rect 3568 1876 3570 1880
rect 3562 1874 3570 1876
rect 3586 1880 3594 1882
rect 3586 1876 3588 1880
rect 3592 1876 3594 1880
rect 3586 1874 3594 1876
rect 3610 1880 3618 1882
rect 3610 1876 3612 1880
rect 3616 1876 3618 1880
rect 3610 1874 3618 1876
rect 3634 1880 3642 1882
rect 3634 1876 3636 1880
rect 3640 1876 3642 1880
rect 3634 1874 3642 1876
rect 3658 1880 3666 1882
rect 3658 1876 3660 1880
rect 3664 1876 3666 1880
rect 3658 1874 3666 1876
rect 3682 1880 3690 1882
rect 3682 1876 3684 1880
rect 3688 1876 3690 1880
rect 3682 1874 3690 1876
rect 3898 1880 3906 1882
rect 3898 1876 3900 1880
rect 3904 1876 3906 1880
rect 3898 1874 3906 1876
rect 3922 1880 3930 1882
rect 3922 1876 3924 1880
rect 3928 1876 3930 1880
rect 3922 1874 3930 1876
rect 3946 1880 3954 1882
rect 3946 1876 3948 1880
rect 3952 1876 3954 1880
rect 3946 1874 3954 1876
rect 3970 1880 3978 1882
rect 3970 1876 3972 1880
rect 3976 1876 3978 1880
rect 3970 1874 3978 1876
rect 3994 1880 4002 1882
rect 3994 1876 3996 1880
rect 4000 1876 4002 1880
rect 3994 1874 4002 1876
rect 4018 1880 4026 1882
rect 4018 1876 4020 1880
rect 4024 1876 4026 1880
rect 4018 1874 4026 1876
rect 4042 1880 4050 1882
rect 4042 1876 4044 1880
rect 4048 1876 4050 1880
rect 4042 1874 4050 1876
rect 4066 1880 4074 1882
rect 4066 1876 4068 1880
rect 4072 1876 4074 1880
rect 4066 1874 4074 1876
rect 4090 1880 4098 1882
rect 4090 1876 4092 1880
rect 4096 1876 4098 1880
rect 4090 1874 4098 1876
rect 4114 1880 4122 1882
rect 4114 1876 4116 1880
rect 4120 1876 4122 1880
rect 4114 1874 4122 1876
rect 4138 1880 4146 1882
rect 4138 1876 4140 1880
rect 4144 1876 4146 1880
rect 4138 1874 4146 1876
rect 4162 1880 4170 1882
rect 4162 1876 4164 1880
rect 4168 1876 4170 1880
rect 4162 1874 4170 1876
rect 4186 1880 4194 1882
rect 4186 1876 4188 1880
rect 4192 1876 4194 1880
rect 4186 1874 4194 1876
rect 4210 1880 4218 1882
rect 4210 1876 4212 1880
rect 4216 1876 4218 1880
rect 4210 1874 4218 1876
rect 4234 1880 4242 1882
rect 4234 1876 4236 1880
rect 4240 1876 4242 1880
rect 4234 1874 4242 1876
rect 4258 1880 4266 1882
rect 4258 1876 4260 1880
rect 4264 1876 4266 1880
rect 4258 1874 4266 1876
rect 4282 1880 4290 1882
rect 4282 1876 4284 1880
rect 4288 1876 4290 1880
rect 4282 1874 4290 1876
rect 4498 1880 4506 1882
rect 4498 1876 4500 1880
rect 4504 1876 4506 1880
rect 4498 1874 4506 1876
rect 4522 1880 4530 1882
rect 4522 1876 4524 1880
rect 4528 1876 4530 1880
rect 4522 1874 4530 1876
rect 4546 1880 4554 1882
rect 4546 1876 4548 1880
rect 4552 1876 4554 1880
rect 4546 1874 4554 1876
rect 4570 1880 4578 1882
rect 4570 1876 4572 1880
rect 4576 1876 4578 1880
rect 4570 1874 4578 1876
rect 4594 1880 4602 1882
rect 4594 1876 4596 1880
rect 4600 1876 4602 1880
rect 4594 1874 4602 1876
rect 4618 1880 4626 1882
rect 4618 1876 4620 1880
rect 4624 1876 4626 1880
rect 4618 1874 4626 1876
rect 4642 1880 4650 1882
rect 4642 1876 4644 1880
rect 4648 1876 4650 1880
rect 4642 1874 4650 1876
rect 4666 1880 4674 1882
rect 4666 1876 4668 1880
rect 4672 1876 4674 1880
rect 4666 1874 4674 1876
rect 4690 1880 4698 1882
rect 4690 1876 4692 1880
rect 4696 1876 4698 1880
rect 4690 1874 4698 1876
rect 4714 1880 4722 1882
rect 4714 1876 4716 1880
rect 4720 1876 4722 1880
rect 4714 1874 4722 1876
rect 4738 1880 4746 1882
rect 4738 1876 4740 1880
rect 4744 1876 4746 1880
rect 4738 1874 4746 1876
rect 4762 1880 4770 1882
rect 4762 1876 4764 1880
rect 4768 1876 4770 1880
rect 4762 1874 4770 1876
rect 4786 1880 4794 1882
rect 4786 1876 4788 1880
rect 4792 1876 4794 1880
rect 4786 1874 4794 1876
rect 5698 1880 5706 1882
rect 5698 1876 5700 1880
rect 5704 1876 5706 1880
rect 5698 1874 5706 1876
rect 5722 1880 5730 1882
rect 5722 1876 5724 1880
rect 5728 1876 5730 1880
rect 5722 1874 5730 1876
rect 5746 1880 5754 1882
rect 5746 1876 5748 1880
rect 5752 1876 5754 1880
rect 5746 1874 5754 1876
rect 5770 1880 5778 1882
rect 5770 1876 5772 1880
rect 5776 1876 5778 1880
rect 5770 1874 5778 1876
rect 5794 1880 5802 1882
rect 5794 1876 5796 1880
rect 5800 1876 5802 1880
rect 5794 1874 5802 1876
rect 5818 1880 5826 1882
rect 5818 1876 5820 1880
rect 5824 1876 5826 1880
rect 5818 1874 5826 1876
rect 5842 1880 5850 1882
rect 5842 1876 5844 1880
rect 5848 1876 5850 1880
rect 5842 1874 5850 1876
rect 5866 1880 5874 1882
rect 5866 1876 5868 1880
rect 5872 1876 5874 1880
rect 5866 1874 5874 1876
rect 5890 1880 5898 1882
rect 5890 1876 5892 1880
rect 5896 1876 5898 1880
rect 5890 1874 5898 1876
rect 5914 1880 5922 1882
rect 5914 1876 5916 1880
rect 5920 1876 5922 1880
rect 5914 1874 5922 1876
rect 5938 1880 5946 1882
rect 5938 1876 5940 1880
rect 5944 1876 5946 1880
rect 5938 1874 5946 1876
rect 5962 1880 5970 1882
rect 5962 1876 5964 1880
rect 5968 1876 5970 1880
rect 5962 1874 5970 1876
rect 5986 1880 5994 1882
rect 5986 1876 5988 1880
rect 5992 1876 5994 1880
rect 5986 1874 5994 1876
rect 6010 1880 6018 1882
rect 6010 1876 6012 1880
rect 6016 1876 6018 1880
rect 6010 1874 6018 1876
rect 6034 1880 6042 1882
rect 6034 1876 6036 1880
rect 6040 1876 6042 1880
rect 6034 1874 6042 1876
rect 6058 1880 6066 1882
rect 6058 1876 6060 1880
rect 6064 1876 6066 1880
rect 6058 1874 6066 1876
rect 6082 1880 6090 1882
rect 6082 1876 6084 1880
rect 6088 1876 6090 1880
rect 6082 1874 6090 1876
rect 6298 1880 6306 1882
rect 6298 1876 6300 1880
rect 6304 1876 6306 1880
rect 6298 1874 6306 1876
rect 6322 1880 6330 1882
rect 6322 1876 6324 1880
rect 6328 1876 6330 1880
rect 6322 1874 6330 1876
rect 6346 1880 6354 1882
rect 6346 1876 6348 1880
rect 6352 1876 6354 1880
rect 6346 1874 6354 1876
rect 6370 1880 6378 1882
rect 6370 1876 6372 1880
rect 6376 1876 6378 1880
rect 6370 1874 6378 1876
rect 6394 1880 6402 1882
rect 6394 1876 6396 1880
rect 6400 1876 6402 1880
rect 6394 1874 6402 1876
rect 6418 1880 6426 1882
rect 6418 1876 6420 1880
rect 6424 1876 6426 1880
rect 6418 1874 6426 1876
rect 6442 1880 6450 1882
rect 6442 1876 6444 1880
rect 6448 1876 6450 1880
rect 6442 1874 6450 1876
rect 6466 1880 6474 1882
rect 6466 1876 6468 1880
rect 6472 1876 6474 1880
rect 6466 1874 6474 1876
rect 6490 1880 6498 1882
rect 6490 1876 6492 1880
rect 6496 1876 6498 1880
rect 6490 1874 6498 1876
rect 6514 1880 6522 1882
rect 6514 1876 6516 1880
rect 6520 1876 6522 1880
rect 6514 1874 6522 1876
rect 6538 1880 6546 1882
rect 6538 1876 6540 1880
rect 6544 1876 6546 1880
rect 6538 1874 6546 1876
rect 6562 1880 6570 1882
rect 6562 1876 6564 1880
rect 6568 1876 6570 1880
rect 6562 1874 6570 1876
rect 6586 1880 6594 1882
rect 6586 1876 6588 1880
rect 6592 1876 6594 1880
rect 6586 1874 6594 1876
rect 6610 1880 6618 1882
rect 6610 1876 6612 1880
rect 6616 1876 6618 1880
rect 6610 1874 6618 1876
rect 6634 1880 6642 1882
rect 6634 1876 6636 1880
rect 6640 1876 6642 1880
rect 6634 1874 6642 1876
rect 6658 1880 6666 1882
rect 6658 1876 6660 1880
rect 6664 1876 6666 1880
rect 6658 1874 6666 1876
rect 6682 1880 6690 1882
rect 6682 1876 6684 1880
rect 6688 1876 6690 1880
rect 6682 1874 6690 1876
rect 6898 1880 6906 1882
rect 6898 1876 6900 1880
rect 6904 1876 6906 1880
rect 6898 1874 6906 1876
rect 6922 1880 6930 1882
rect 6922 1876 6924 1880
rect 6928 1876 6930 1880
rect 6922 1874 6930 1876
rect 6946 1880 6954 1882
rect 6946 1876 6948 1880
rect 6952 1876 6954 1880
rect 6946 1874 6954 1876
rect 6970 1880 6978 1882
rect 6970 1876 6972 1880
rect 6976 1876 6978 1880
rect 6970 1874 6978 1876
rect 6994 1880 7002 1882
rect 6994 1876 6996 1880
rect 7000 1876 7002 1880
rect 6994 1874 7002 1876
rect 7018 1880 7026 1882
rect 7018 1876 7020 1880
rect 7024 1876 7026 1880
rect 7018 1874 7026 1876
rect 7042 1880 7050 1882
rect 7042 1876 7044 1880
rect 7048 1876 7050 1880
rect 7042 1874 7050 1876
rect 7066 1880 7074 1882
rect 7066 1876 7068 1880
rect 7072 1876 7074 1880
rect 7066 1874 7074 1876
rect 7090 1880 7098 1882
rect 7090 1876 7092 1880
rect 7096 1876 7098 1880
rect 7090 1874 7098 1876
rect 7114 1880 7122 1882
rect 7114 1876 7116 1880
rect 7120 1876 7122 1880
rect 7114 1874 7122 1876
rect 7138 1880 7146 1882
rect 7138 1876 7140 1880
rect 7144 1876 7146 1880
rect 7138 1874 7146 1876
rect 7162 1880 7170 1882
rect 7162 1876 7164 1880
rect 7168 1876 7170 1880
rect 7162 1874 7170 1876
rect 7186 1880 7194 1882
rect 7186 1876 7188 1880
rect 7192 1876 7194 1880
rect 7186 1874 7194 1876
rect 2400 1868 2406 1870
rect 2404 1864 2406 1868
rect 2400 1862 2406 1864
rect 2422 1868 2430 1870
rect 2422 1864 2424 1868
rect 2428 1864 2430 1868
rect 2422 1862 2430 1864
rect 2446 1868 2454 1870
rect 2446 1864 2448 1868
rect 2452 1864 2454 1868
rect 2446 1862 2454 1864
rect 2470 1868 2478 1870
rect 2470 1864 2472 1868
rect 2476 1864 2478 1868
rect 2470 1862 2478 1864
rect 2494 1868 2502 1870
rect 2494 1864 2496 1868
rect 2500 1864 2502 1868
rect 2494 1862 2502 1864
rect 2710 1868 2718 1870
rect 2710 1864 2712 1868
rect 2716 1864 2718 1868
rect 2710 1862 2718 1864
rect 2734 1868 2742 1870
rect 2734 1864 2736 1868
rect 2740 1864 2742 1868
rect 2734 1862 2742 1864
rect 2758 1868 2766 1870
rect 2758 1864 2760 1868
rect 2764 1864 2766 1868
rect 2758 1862 2766 1864
rect 2782 1868 2790 1870
rect 2782 1864 2784 1868
rect 2788 1864 2790 1868
rect 2782 1862 2790 1864
rect 2806 1868 2814 1870
rect 2806 1864 2808 1868
rect 2812 1864 2814 1868
rect 2806 1862 2814 1864
rect 2830 1868 2838 1870
rect 2830 1864 2832 1868
rect 2836 1864 2838 1868
rect 2830 1862 2838 1864
rect 2854 1868 2862 1870
rect 2854 1864 2856 1868
rect 2860 1864 2862 1868
rect 2854 1862 2862 1864
rect 2878 1868 2886 1870
rect 2878 1864 2880 1868
rect 2884 1864 2886 1868
rect 2878 1862 2886 1864
rect 2902 1868 2910 1870
rect 2902 1864 2904 1868
rect 2908 1864 2910 1868
rect 2902 1862 2910 1864
rect 2926 1868 2934 1870
rect 2926 1864 2928 1868
rect 2932 1864 2934 1868
rect 2926 1862 2934 1864
rect 2950 1868 2958 1870
rect 2950 1864 2952 1868
rect 2956 1864 2958 1868
rect 2950 1862 2958 1864
rect 2974 1868 2982 1870
rect 2974 1864 2976 1868
rect 2980 1864 2982 1868
rect 2974 1862 2982 1864
rect 2998 1868 3006 1870
rect 2998 1864 3000 1868
rect 3004 1864 3006 1868
rect 2998 1862 3006 1864
rect 3022 1868 3030 1870
rect 3022 1864 3024 1868
rect 3028 1864 3030 1868
rect 3022 1862 3030 1864
rect 3046 1868 3054 1870
rect 3046 1864 3048 1868
rect 3052 1864 3054 1868
rect 3046 1862 3054 1864
rect 3070 1868 3078 1870
rect 3070 1864 3072 1868
rect 3076 1864 3078 1868
rect 3070 1862 3078 1864
rect 3094 1868 3102 1870
rect 3094 1864 3096 1868
rect 3100 1864 3102 1868
rect 3094 1862 3102 1864
rect 3310 1868 3318 1870
rect 3310 1864 3312 1868
rect 3316 1864 3318 1868
rect 3310 1862 3318 1864
rect 3334 1868 3342 1870
rect 3334 1864 3336 1868
rect 3340 1864 3342 1868
rect 3334 1862 3342 1864
rect 3358 1868 3366 1870
rect 3358 1864 3360 1868
rect 3364 1864 3366 1868
rect 3358 1862 3366 1864
rect 3382 1868 3390 1870
rect 3382 1864 3384 1868
rect 3388 1864 3390 1868
rect 3382 1862 3390 1864
rect 3406 1868 3414 1870
rect 3406 1864 3408 1868
rect 3412 1864 3414 1868
rect 3406 1862 3414 1864
rect 3430 1868 3438 1870
rect 3430 1864 3432 1868
rect 3436 1864 3438 1868
rect 3430 1862 3438 1864
rect 3454 1868 3462 1870
rect 3454 1864 3456 1868
rect 3460 1864 3462 1868
rect 3454 1862 3462 1864
rect 3478 1868 3486 1870
rect 3478 1864 3480 1868
rect 3484 1864 3486 1868
rect 3478 1862 3486 1864
rect 3502 1868 3510 1870
rect 3502 1864 3504 1868
rect 3508 1864 3510 1868
rect 3502 1862 3510 1864
rect 3526 1868 3534 1870
rect 3526 1864 3528 1868
rect 3532 1864 3534 1868
rect 3526 1862 3534 1864
rect 3550 1868 3558 1870
rect 3550 1864 3552 1868
rect 3556 1864 3558 1868
rect 3550 1862 3558 1864
rect 3574 1868 3582 1870
rect 3574 1864 3576 1868
rect 3580 1864 3582 1868
rect 3574 1862 3582 1864
rect 3598 1868 3606 1870
rect 3598 1864 3600 1868
rect 3604 1864 3606 1868
rect 3598 1862 3606 1864
rect 3622 1868 3630 1870
rect 3622 1864 3624 1868
rect 3628 1864 3630 1868
rect 3622 1862 3630 1864
rect 3646 1868 3654 1870
rect 3646 1864 3648 1868
rect 3652 1864 3654 1868
rect 3646 1862 3654 1864
rect 3670 1868 3678 1870
rect 3670 1864 3672 1868
rect 3676 1864 3678 1868
rect 3670 1862 3678 1864
rect 3694 1868 3702 1870
rect 3694 1864 3696 1868
rect 3700 1864 3702 1868
rect 3694 1862 3702 1864
rect 3910 1868 3918 1870
rect 3910 1864 3912 1868
rect 3916 1864 3918 1868
rect 3910 1862 3918 1864
rect 3934 1868 3942 1870
rect 3934 1864 3936 1868
rect 3940 1864 3942 1868
rect 3934 1862 3942 1864
rect 3958 1868 3966 1870
rect 3958 1864 3960 1868
rect 3964 1864 3966 1868
rect 3958 1862 3966 1864
rect 3982 1868 3990 1870
rect 3982 1864 3984 1868
rect 3988 1864 3990 1868
rect 3982 1862 3990 1864
rect 4006 1868 4014 1870
rect 4006 1864 4008 1868
rect 4012 1864 4014 1868
rect 4006 1862 4014 1864
rect 4030 1868 4038 1870
rect 4030 1864 4032 1868
rect 4036 1864 4038 1868
rect 4030 1862 4038 1864
rect 4054 1868 4062 1870
rect 4054 1864 4056 1868
rect 4060 1864 4062 1868
rect 4054 1862 4062 1864
rect 4078 1868 4086 1870
rect 4078 1864 4080 1868
rect 4084 1864 4086 1868
rect 4078 1862 4086 1864
rect 4102 1868 4110 1870
rect 4102 1864 4104 1868
rect 4108 1864 4110 1868
rect 4102 1862 4110 1864
rect 4126 1868 4134 1870
rect 4126 1864 4128 1868
rect 4132 1864 4134 1868
rect 4126 1862 4134 1864
rect 4150 1868 4158 1870
rect 4150 1864 4152 1868
rect 4156 1864 4158 1868
rect 4150 1862 4158 1864
rect 4174 1868 4182 1870
rect 4174 1864 4176 1868
rect 4180 1864 4182 1868
rect 4174 1862 4182 1864
rect 4198 1868 4206 1870
rect 4198 1864 4200 1868
rect 4204 1864 4206 1868
rect 4198 1862 4206 1864
rect 4222 1868 4230 1870
rect 4222 1864 4224 1868
rect 4228 1864 4230 1868
rect 4222 1862 4230 1864
rect 4246 1868 4254 1870
rect 4246 1864 4248 1868
rect 4252 1864 4254 1868
rect 4246 1862 4254 1864
rect 4270 1868 4278 1870
rect 4270 1864 4272 1868
rect 4276 1864 4278 1868
rect 4270 1862 4278 1864
rect 4294 1868 4302 1870
rect 4294 1864 4296 1868
rect 4300 1864 4302 1868
rect 4294 1862 4302 1864
rect 4510 1868 4518 1870
rect 4510 1864 4512 1868
rect 4516 1864 4518 1868
rect 4510 1862 4518 1864
rect 4534 1868 4542 1870
rect 4534 1864 4536 1868
rect 4540 1864 4542 1868
rect 4534 1862 4542 1864
rect 4558 1868 4566 1870
rect 4558 1864 4560 1868
rect 4564 1864 4566 1868
rect 4558 1862 4566 1864
rect 4582 1868 4590 1870
rect 4582 1864 4584 1868
rect 4588 1864 4590 1868
rect 4582 1862 4590 1864
rect 4606 1868 4614 1870
rect 4606 1864 4608 1868
rect 4612 1864 4614 1868
rect 4606 1862 4614 1864
rect 4630 1868 4638 1870
rect 4630 1864 4632 1868
rect 4636 1864 4638 1868
rect 4630 1862 4638 1864
rect 4654 1868 4662 1870
rect 4654 1864 4656 1868
rect 4660 1864 4662 1868
rect 4654 1862 4662 1864
rect 4678 1868 4686 1870
rect 4678 1864 4680 1868
rect 4684 1864 4686 1868
rect 4678 1862 4686 1864
rect 4702 1868 4710 1870
rect 4702 1864 4704 1868
rect 4708 1864 4710 1868
rect 4702 1862 4710 1864
rect 4726 1868 4734 1870
rect 4726 1864 4728 1868
rect 4732 1864 4734 1868
rect 4726 1862 4734 1864
rect 4750 1868 4758 1870
rect 4750 1864 4752 1868
rect 4756 1864 4758 1868
rect 4750 1862 4758 1864
rect 4774 1868 4782 1870
rect 4774 1864 4776 1868
rect 4780 1864 4782 1868
rect 4774 1862 4782 1864
rect 4798 1862 4800 1870
rect 5710 1868 5718 1870
rect 5710 1864 5712 1868
rect 5716 1864 5718 1868
rect 5710 1862 5718 1864
rect 5734 1868 5742 1870
rect 5734 1864 5736 1868
rect 5740 1864 5742 1868
rect 5734 1862 5742 1864
rect 5758 1868 5766 1870
rect 5758 1864 5760 1868
rect 5764 1864 5766 1868
rect 5758 1862 5766 1864
rect 5782 1868 5790 1870
rect 5782 1864 5784 1868
rect 5788 1864 5790 1868
rect 5782 1862 5790 1864
rect 5806 1868 5814 1870
rect 5806 1864 5808 1868
rect 5812 1864 5814 1868
rect 5806 1862 5814 1864
rect 5830 1868 5838 1870
rect 5830 1864 5832 1868
rect 5836 1864 5838 1868
rect 5830 1862 5838 1864
rect 5854 1868 5862 1870
rect 5854 1864 5856 1868
rect 5860 1864 5862 1868
rect 5854 1862 5862 1864
rect 5878 1868 5886 1870
rect 5878 1864 5880 1868
rect 5884 1864 5886 1868
rect 5878 1862 5886 1864
rect 5902 1868 5910 1870
rect 5902 1864 5904 1868
rect 5908 1864 5910 1868
rect 5902 1862 5910 1864
rect 5926 1868 5934 1870
rect 5926 1864 5928 1868
rect 5932 1864 5934 1868
rect 5926 1862 5934 1864
rect 5950 1868 5958 1870
rect 5950 1864 5952 1868
rect 5956 1864 5958 1868
rect 5950 1862 5958 1864
rect 5974 1868 5982 1870
rect 5974 1864 5976 1868
rect 5980 1864 5982 1868
rect 5974 1862 5982 1864
rect 5998 1868 6006 1870
rect 5998 1864 6000 1868
rect 6004 1864 6006 1868
rect 5998 1862 6006 1864
rect 6022 1868 6030 1870
rect 6022 1864 6024 1868
rect 6028 1864 6030 1868
rect 6022 1862 6030 1864
rect 6046 1868 6054 1870
rect 6046 1864 6048 1868
rect 6052 1864 6054 1868
rect 6046 1862 6054 1864
rect 6070 1868 6078 1870
rect 6070 1864 6072 1868
rect 6076 1864 6078 1868
rect 6070 1862 6078 1864
rect 6094 1868 6102 1870
rect 6094 1864 6096 1868
rect 6100 1864 6102 1868
rect 6094 1862 6102 1864
rect 6310 1868 6318 1870
rect 6310 1864 6312 1868
rect 6316 1864 6318 1868
rect 6310 1862 6318 1864
rect 6334 1868 6342 1870
rect 6334 1864 6336 1868
rect 6340 1864 6342 1868
rect 6334 1862 6342 1864
rect 6358 1868 6366 1870
rect 6358 1864 6360 1868
rect 6364 1864 6366 1868
rect 6358 1862 6366 1864
rect 6382 1868 6390 1870
rect 6382 1864 6384 1868
rect 6388 1864 6390 1868
rect 6382 1862 6390 1864
rect 6406 1868 6414 1870
rect 6406 1864 6408 1868
rect 6412 1864 6414 1868
rect 6406 1862 6414 1864
rect 6430 1868 6438 1870
rect 6430 1864 6432 1868
rect 6436 1864 6438 1868
rect 6430 1862 6438 1864
rect 6454 1868 6462 1870
rect 6454 1864 6456 1868
rect 6460 1864 6462 1868
rect 6454 1862 6462 1864
rect 6478 1868 6486 1870
rect 6478 1864 6480 1868
rect 6484 1864 6486 1868
rect 6478 1862 6486 1864
rect 6502 1868 6510 1870
rect 6502 1864 6504 1868
rect 6508 1864 6510 1868
rect 6502 1862 6510 1864
rect 6526 1868 6534 1870
rect 6526 1864 6528 1868
rect 6532 1864 6534 1868
rect 6526 1862 6534 1864
rect 6550 1868 6558 1870
rect 6550 1864 6552 1868
rect 6556 1864 6558 1868
rect 6550 1862 6558 1864
rect 6574 1868 6582 1870
rect 6574 1864 6576 1868
rect 6580 1864 6582 1868
rect 6574 1862 6582 1864
rect 6598 1868 6606 1870
rect 6598 1864 6600 1868
rect 6604 1864 6606 1868
rect 6598 1862 6606 1864
rect 6622 1868 6630 1870
rect 6622 1864 6624 1868
rect 6628 1864 6630 1868
rect 6622 1862 6630 1864
rect 6646 1868 6654 1870
rect 6646 1864 6648 1868
rect 6652 1864 6654 1868
rect 6646 1862 6654 1864
rect 6670 1868 6678 1870
rect 6670 1864 6672 1868
rect 6676 1864 6678 1868
rect 6670 1862 6678 1864
rect 6694 1868 6702 1870
rect 6694 1864 6696 1868
rect 6700 1864 6702 1868
rect 6694 1862 6702 1864
rect 6910 1868 6918 1870
rect 6910 1864 6912 1868
rect 6916 1864 6918 1868
rect 6910 1862 6918 1864
rect 6934 1868 6942 1870
rect 6934 1864 6936 1868
rect 6940 1864 6942 1868
rect 6934 1862 6942 1864
rect 6958 1868 6966 1870
rect 6958 1864 6960 1868
rect 6964 1864 6966 1868
rect 6958 1862 6966 1864
rect 6982 1868 6990 1870
rect 6982 1864 6984 1868
rect 6988 1864 6990 1868
rect 6982 1862 6990 1864
rect 7006 1868 7014 1870
rect 7006 1864 7008 1868
rect 7012 1864 7014 1868
rect 7006 1862 7014 1864
rect 7030 1868 7038 1870
rect 7030 1864 7032 1868
rect 7036 1864 7038 1868
rect 7030 1862 7038 1864
rect 7054 1868 7062 1870
rect 7054 1864 7056 1868
rect 7060 1864 7062 1868
rect 7054 1862 7062 1864
rect 7078 1868 7086 1870
rect 7078 1864 7080 1868
rect 7084 1864 7086 1868
rect 7078 1862 7086 1864
rect 7102 1868 7110 1870
rect 7102 1864 7104 1868
rect 7108 1864 7110 1868
rect 7102 1862 7110 1864
rect 7126 1868 7134 1870
rect 7126 1864 7128 1868
rect 7132 1864 7134 1868
rect 7126 1862 7134 1864
rect 7150 1868 7158 1870
rect 7150 1864 7152 1868
rect 7156 1864 7158 1868
rect 7150 1862 7158 1864
rect 7174 1868 7182 1870
rect 7174 1864 7176 1868
rect 7180 1864 7182 1868
rect 7174 1862 7182 1864
rect 7198 1862 7200 1870
rect 2410 1856 2418 1858
rect 2410 1852 2412 1856
rect 2416 1852 2418 1856
rect 2410 1850 2418 1852
rect 2434 1856 2442 1858
rect 2434 1852 2436 1856
rect 2440 1852 2442 1856
rect 2434 1850 2442 1852
rect 2458 1856 2466 1858
rect 2458 1852 2460 1856
rect 2464 1852 2466 1856
rect 2458 1850 2466 1852
rect 2482 1856 2490 1858
rect 2482 1852 2484 1856
rect 2488 1852 2490 1856
rect 2482 1850 2490 1852
rect 2698 1856 2706 1858
rect 2698 1852 2700 1856
rect 2704 1852 2706 1856
rect 2698 1850 2706 1852
rect 2722 1856 2730 1858
rect 2722 1852 2724 1856
rect 2728 1852 2730 1856
rect 2722 1850 2730 1852
rect 2746 1856 2754 1858
rect 2746 1852 2748 1856
rect 2752 1852 2754 1856
rect 2746 1850 2754 1852
rect 2770 1856 2778 1858
rect 2770 1852 2772 1856
rect 2776 1852 2778 1856
rect 2770 1850 2778 1852
rect 2794 1856 2802 1858
rect 2794 1852 2796 1856
rect 2800 1852 2802 1856
rect 2794 1850 2802 1852
rect 2818 1856 2826 1858
rect 2818 1852 2820 1856
rect 2824 1852 2826 1856
rect 2818 1850 2826 1852
rect 2842 1856 2850 1858
rect 2842 1852 2844 1856
rect 2848 1852 2850 1856
rect 2842 1850 2850 1852
rect 2866 1856 2874 1858
rect 2866 1852 2868 1856
rect 2872 1852 2874 1856
rect 2866 1850 2874 1852
rect 2890 1856 2898 1858
rect 2890 1852 2892 1856
rect 2896 1852 2898 1856
rect 2890 1850 2898 1852
rect 2914 1856 2922 1858
rect 2914 1852 2916 1856
rect 2920 1852 2922 1856
rect 2914 1850 2922 1852
rect 2938 1856 2946 1858
rect 2938 1852 2940 1856
rect 2944 1852 2946 1856
rect 2938 1850 2946 1852
rect 2962 1856 2970 1858
rect 2962 1852 2964 1856
rect 2968 1852 2970 1856
rect 2962 1850 2970 1852
rect 2986 1856 2994 1858
rect 2986 1852 2988 1856
rect 2992 1852 2994 1856
rect 2986 1850 2994 1852
rect 3010 1856 3018 1858
rect 3010 1852 3012 1856
rect 3016 1852 3018 1856
rect 3010 1850 3018 1852
rect 3034 1856 3042 1858
rect 3034 1852 3036 1856
rect 3040 1852 3042 1856
rect 3034 1850 3042 1852
rect 3058 1856 3066 1858
rect 3058 1852 3060 1856
rect 3064 1852 3066 1856
rect 3058 1850 3066 1852
rect 3082 1856 3090 1858
rect 3082 1852 3084 1856
rect 3088 1852 3090 1856
rect 3082 1850 3090 1852
rect 3298 1856 3306 1858
rect 3298 1852 3300 1856
rect 3304 1852 3306 1856
rect 3298 1850 3306 1852
rect 3322 1856 3330 1858
rect 3322 1852 3324 1856
rect 3328 1852 3330 1856
rect 3322 1850 3330 1852
rect 3346 1856 3354 1858
rect 3346 1852 3348 1856
rect 3352 1852 3354 1856
rect 3346 1850 3354 1852
rect 3370 1856 3378 1858
rect 3370 1852 3372 1856
rect 3376 1852 3378 1856
rect 3370 1850 3378 1852
rect 3394 1856 3402 1858
rect 3394 1852 3396 1856
rect 3400 1852 3402 1856
rect 3394 1850 3402 1852
rect 3418 1856 3426 1858
rect 3418 1852 3420 1856
rect 3424 1852 3426 1856
rect 3418 1850 3426 1852
rect 3442 1856 3450 1858
rect 3442 1852 3444 1856
rect 3448 1852 3450 1856
rect 3442 1850 3450 1852
rect 3466 1856 3474 1858
rect 3466 1852 3468 1856
rect 3472 1852 3474 1856
rect 3466 1850 3474 1852
rect 3490 1856 3498 1858
rect 3490 1852 3492 1856
rect 3496 1852 3498 1856
rect 3490 1850 3498 1852
rect 3514 1856 3522 1858
rect 3514 1852 3516 1856
rect 3520 1852 3522 1856
rect 3514 1850 3522 1852
rect 3538 1856 3546 1858
rect 3538 1852 3540 1856
rect 3544 1852 3546 1856
rect 3538 1850 3546 1852
rect 3562 1856 3570 1858
rect 3562 1852 3564 1856
rect 3568 1852 3570 1856
rect 3562 1850 3570 1852
rect 3586 1856 3594 1858
rect 3586 1852 3588 1856
rect 3592 1852 3594 1856
rect 3586 1850 3594 1852
rect 3610 1856 3618 1858
rect 3610 1852 3612 1856
rect 3616 1852 3618 1856
rect 3610 1850 3618 1852
rect 3634 1856 3642 1858
rect 3634 1852 3636 1856
rect 3640 1852 3642 1856
rect 3634 1850 3642 1852
rect 3658 1856 3666 1858
rect 3658 1852 3660 1856
rect 3664 1852 3666 1856
rect 3658 1850 3666 1852
rect 3682 1856 3690 1858
rect 3682 1852 3684 1856
rect 3688 1852 3690 1856
rect 3682 1850 3690 1852
rect 3898 1856 3906 1858
rect 3898 1852 3900 1856
rect 3904 1852 3906 1856
rect 3898 1850 3906 1852
rect 3922 1856 3930 1858
rect 3922 1852 3924 1856
rect 3928 1852 3930 1856
rect 3922 1850 3930 1852
rect 3946 1856 3954 1858
rect 3946 1852 3948 1856
rect 3952 1852 3954 1856
rect 3946 1850 3954 1852
rect 3970 1856 3978 1858
rect 3970 1852 3972 1856
rect 3976 1852 3978 1856
rect 3970 1850 3978 1852
rect 3994 1856 4002 1858
rect 3994 1852 3996 1856
rect 4000 1852 4002 1856
rect 3994 1850 4002 1852
rect 4018 1856 4026 1858
rect 4018 1852 4020 1856
rect 4024 1852 4026 1856
rect 4018 1850 4026 1852
rect 4042 1856 4050 1858
rect 4042 1852 4044 1856
rect 4048 1852 4050 1856
rect 4042 1850 4050 1852
rect 4066 1856 4074 1858
rect 4066 1852 4068 1856
rect 4072 1852 4074 1856
rect 4066 1850 4074 1852
rect 4090 1856 4098 1858
rect 4090 1852 4092 1856
rect 4096 1852 4098 1856
rect 4090 1850 4098 1852
rect 4114 1856 4122 1858
rect 4114 1852 4116 1856
rect 4120 1852 4122 1856
rect 4114 1850 4122 1852
rect 4138 1856 4146 1858
rect 4138 1852 4140 1856
rect 4144 1852 4146 1856
rect 4138 1850 4146 1852
rect 4162 1856 4170 1858
rect 4162 1852 4164 1856
rect 4168 1852 4170 1856
rect 4162 1850 4170 1852
rect 4186 1856 4194 1858
rect 4186 1852 4188 1856
rect 4192 1852 4194 1856
rect 4186 1850 4194 1852
rect 4210 1856 4218 1858
rect 4210 1852 4212 1856
rect 4216 1852 4218 1856
rect 4210 1850 4218 1852
rect 4234 1856 4242 1858
rect 4234 1852 4236 1856
rect 4240 1852 4242 1856
rect 4234 1850 4242 1852
rect 4258 1856 4266 1858
rect 4258 1852 4260 1856
rect 4264 1852 4266 1856
rect 4258 1850 4266 1852
rect 4282 1856 4290 1858
rect 4282 1852 4284 1856
rect 4288 1852 4290 1856
rect 4282 1850 4290 1852
rect 4498 1856 4506 1858
rect 4498 1852 4500 1856
rect 4504 1852 4506 1856
rect 4498 1850 4506 1852
rect 4522 1856 4530 1858
rect 4522 1852 4524 1856
rect 4528 1852 4530 1856
rect 4522 1850 4530 1852
rect 4546 1856 4554 1858
rect 4546 1852 4548 1856
rect 4552 1852 4554 1856
rect 4546 1850 4554 1852
rect 4570 1856 4578 1858
rect 4570 1852 4572 1856
rect 4576 1852 4578 1856
rect 4570 1850 4578 1852
rect 4594 1856 4602 1858
rect 4594 1852 4596 1856
rect 4600 1852 4602 1856
rect 4594 1850 4602 1852
rect 4618 1856 4626 1858
rect 4618 1852 4620 1856
rect 4624 1852 4626 1856
rect 4618 1850 4626 1852
rect 4642 1856 4650 1858
rect 4642 1852 4644 1856
rect 4648 1852 4650 1856
rect 4642 1850 4650 1852
rect 4666 1856 4674 1858
rect 4666 1852 4668 1856
rect 4672 1852 4674 1856
rect 4666 1850 4674 1852
rect 4690 1856 4698 1858
rect 4690 1852 4692 1856
rect 4696 1852 4698 1856
rect 4690 1850 4698 1852
rect 4714 1856 4722 1858
rect 4714 1852 4716 1856
rect 4720 1852 4722 1856
rect 4714 1850 4722 1852
rect 4738 1856 4746 1858
rect 4738 1852 4740 1856
rect 4744 1852 4746 1856
rect 4738 1850 4746 1852
rect 4762 1856 4770 1858
rect 4762 1852 4764 1856
rect 4768 1852 4770 1856
rect 4762 1850 4770 1852
rect 4786 1856 4794 1858
rect 4786 1852 4788 1856
rect 4792 1852 4794 1856
rect 4786 1850 4794 1852
rect 5698 1856 5706 1858
rect 5698 1852 5700 1856
rect 5704 1852 5706 1856
rect 5698 1850 5706 1852
rect 5722 1856 5730 1858
rect 5722 1852 5724 1856
rect 5728 1852 5730 1856
rect 5722 1850 5730 1852
rect 5746 1856 5754 1858
rect 5746 1852 5748 1856
rect 5752 1852 5754 1856
rect 5746 1850 5754 1852
rect 5770 1856 5778 1858
rect 5770 1852 5772 1856
rect 5776 1852 5778 1856
rect 5770 1850 5778 1852
rect 5794 1856 5802 1858
rect 5794 1852 5796 1856
rect 5800 1852 5802 1856
rect 5794 1850 5802 1852
rect 5818 1856 5826 1858
rect 5818 1852 5820 1856
rect 5824 1852 5826 1856
rect 5818 1850 5826 1852
rect 5842 1856 5850 1858
rect 5842 1852 5844 1856
rect 5848 1852 5850 1856
rect 5842 1850 5850 1852
rect 5866 1856 5874 1858
rect 5866 1852 5868 1856
rect 5872 1852 5874 1856
rect 5866 1850 5874 1852
rect 5890 1856 5898 1858
rect 5890 1852 5892 1856
rect 5896 1852 5898 1856
rect 5890 1850 5898 1852
rect 5914 1856 5922 1858
rect 5914 1852 5916 1856
rect 5920 1852 5922 1856
rect 5914 1850 5922 1852
rect 5938 1856 5946 1858
rect 5938 1852 5940 1856
rect 5944 1852 5946 1856
rect 5938 1850 5946 1852
rect 5962 1856 5970 1858
rect 5962 1852 5964 1856
rect 5968 1852 5970 1856
rect 5962 1850 5970 1852
rect 5986 1856 5994 1858
rect 5986 1852 5988 1856
rect 5992 1852 5994 1856
rect 5986 1850 5994 1852
rect 6010 1856 6018 1858
rect 6010 1852 6012 1856
rect 6016 1852 6018 1856
rect 6010 1850 6018 1852
rect 6034 1856 6042 1858
rect 6034 1852 6036 1856
rect 6040 1852 6042 1856
rect 6034 1850 6042 1852
rect 6058 1856 6066 1858
rect 6058 1852 6060 1856
rect 6064 1852 6066 1856
rect 6058 1850 6066 1852
rect 6082 1856 6090 1858
rect 6082 1852 6084 1856
rect 6088 1852 6090 1856
rect 6082 1850 6090 1852
rect 6298 1856 6306 1858
rect 6298 1852 6300 1856
rect 6304 1852 6306 1856
rect 6298 1850 6306 1852
rect 6322 1856 6330 1858
rect 6322 1852 6324 1856
rect 6328 1852 6330 1856
rect 6322 1850 6330 1852
rect 6346 1856 6354 1858
rect 6346 1852 6348 1856
rect 6352 1852 6354 1856
rect 6346 1850 6354 1852
rect 6370 1856 6378 1858
rect 6370 1852 6372 1856
rect 6376 1852 6378 1856
rect 6370 1850 6378 1852
rect 6394 1856 6402 1858
rect 6394 1852 6396 1856
rect 6400 1852 6402 1856
rect 6394 1850 6402 1852
rect 6418 1856 6426 1858
rect 6418 1852 6420 1856
rect 6424 1852 6426 1856
rect 6418 1850 6426 1852
rect 6442 1856 6450 1858
rect 6442 1852 6444 1856
rect 6448 1852 6450 1856
rect 6442 1850 6450 1852
rect 6466 1856 6474 1858
rect 6466 1852 6468 1856
rect 6472 1852 6474 1856
rect 6466 1850 6474 1852
rect 6490 1856 6498 1858
rect 6490 1852 6492 1856
rect 6496 1852 6498 1856
rect 6490 1850 6498 1852
rect 6514 1856 6522 1858
rect 6514 1852 6516 1856
rect 6520 1852 6522 1856
rect 6514 1850 6522 1852
rect 6538 1856 6546 1858
rect 6538 1852 6540 1856
rect 6544 1852 6546 1856
rect 6538 1850 6546 1852
rect 6562 1856 6570 1858
rect 6562 1852 6564 1856
rect 6568 1852 6570 1856
rect 6562 1850 6570 1852
rect 6586 1856 6594 1858
rect 6586 1852 6588 1856
rect 6592 1852 6594 1856
rect 6586 1850 6594 1852
rect 6610 1856 6618 1858
rect 6610 1852 6612 1856
rect 6616 1852 6618 1856
rect 6610 1850 6618 1852
rect 6634 1856 6642 1858
rect 6634 1852 6636 1856
rect 6640 1852 6642 1856
rect 6634 1850 6642 1852
rect 6658 1856 6666 1858
rect 6658 1852 6660 1856
rect 6664 1852 6666 1856
rect 6658 1850 6666 1852
rect 6682 1856 6690 1858
rect 6682 1852 6684 1856
rect 6688 1852 6690 1856
rect 6682 1850 6690 1852
rect 6898 1856 6906 1858
rect 6898 1852 6900 1856
rect 6904 1852 6906 1856
rect 6898 1850 6906 1852
rect 6922 1856 6930 1858
rect 6922 1852 6924 1856
rect 6928 1852 6930 1856
rect 6922 1850 6930 1852
rect 6946 1856 6954 1858
rect 6946 1852 6948 1856
rect 6952 1852 6954 1856
rect 6946 1850 6954 1852
rect 6970 1856 6978 1858
rect 6970 1852 6972 1856
rect 6976 1852 6978 1856
rect 6970 1850 6978 1852
rect 6994 1856 7002 1858
rect 6994 1852 6996 1856
rect 7000 1852 7002 1856
rect 6994 1850 7002 1852
rect 7018 1856 7026 1858
rect 7018 1852 7020 1856
rect 7024 1852 7026 1856
rect 7018 1850 7026 1852
rect 7042 1856 7050 1858
rect 7042 1852 7044 1856
rect 7048 1852 7050 1856
rect 7042 1850 7050 1852
rect 7066 1856 7074 1858
rect 7066 1852 7068 1856
rect 7072 1852 7074 1856
rect 7066 1850 7074 1852
rect 7090 1856 7098 1858
rect 7090 1852 7092 1856
rect 7096 1852 7098 1856
rect 7090 1850 7098 1852
rect 7114 1856 7122 1858
rect 7114 1852 7116 1856
rect 7120 1852 7122 1856
rect 7114 1850 7122 1852
rect 7138 1856 7146 1858
rect 7138 1852 7140 1856
rect 7144 1852 7146 1856
rect 7138 1850 7146 1852
rect 7162 1856 7170 1858
rect 7162 1852 7164 1856
rect 7168 1852 7170 1856
rect 7162 1850 7170 1852
rect 7186 1856 7194 1858
rect 7186 1852 7188 1856
rect 7192 1852 7194 1856
rect 7186 1850 7194 1852
rect 2400 1844 2406 1846
rect 2404 1840 2406 1844
rect 2400 1838 2406 1840
rect 2422 1844 2430 1846
rect 2422 1840 2424 1844
rect 2428 1840 2430 1844
rect 2422 1838 2430 1840
rect 2446 1844 2454 1846
rect 2446 1840 2448 1844
rect 2452 1840 2454 1844
rect 2446 1838 2454 1840
rect 2470 1844 2478 1846
rect 2470 1840 2472 1844
rect 2476 1840 2478 1844
rect 2470 1838 2478 1840
rect 2494 1844 2502 1846
rect 2494 1840 2496 1844
rect 2500 1840 2502 1844
rect 2494 1838 2502 1840
rect 2710 1844 2718 1846
rect 2710 1840 2712 1844
rect 2716 1840 2718 1844
rect 2710 1838 2718 1840
rect 2734 1844 2742 1846
rect 2734 1840 2736 1844
rect 2740 1840 2742 1844
rect 2734 1838 2742 1840
rect 2758 1844 2766 1846
rect 2758 1840 2760 1844
rect 2764 1840 2766 1844
rect 2758 1838 2766 1840
rect 2782 1844 2790 1846
rect 2782 1840 2784 1844
rect 2788 1840 2790 1844
rect 2782 1838 2790 1840
rect 2806 1844 2814 1846
rect 2806 1840 2808 1844
rect 2812 1840 2814 1844
rect 2806 1838 2814 1840
rect 2830 1844 2838 1846
rect 2830 1840 2832 1844
rect 2836 1840 2838 1844
rect 2830 1838 2838 1840
rect 2854 1844 2862 1846
rect 2854 1840 2856 1844
rect 2860 1840 2862 1844
rect 2854 1838 2862 1840
rect 2878 1844 2886 1846
rect 2878 1840 2880 1844
rect 2884 1840 2886 1844
rect 2878 1838 2886 1840
rect 2902 1844 2910 1846
rect 2902 1840 2904 1844
rect 2908 1840 2910 1844
rect 2902 1838 2910 1840
rect 2926 1844 2934 1846
rect 2926 1840 2928 1844
rect 2932 1840 2934 1844
rect 2926 1838 2934 1840
rect 2950 1844 2958 1846
rect 2950 1840 2952 1844
rect 2956 1840 2958 1844
rect 2950 1838 2958 1840
rect 2974 1844 2982 1846
rect 2974 1840 2976 1844
rect 2980 1840 2982 1844
rect 2974 1838 2982 1840
rect 2998 1844 3006 1846
rect 2998 1840 3000 1844
rect 3004 1840 3006 1844
rect 2998 1838 3006 1840
rect 3022 1844 3030 1846
rect 3022 1840 3024 1844
rect 3028 1840 3030 1844
rect 3022 1838 3030 1840
rect 3046 1844 3054 1846
rect 3046 1840 3048 1844
rect 3052 1840 3054 1844
rect 3046 1838 3054 1840
rect 3070 1844 3078 1846
rect 3070 1840 3072 1844
rect 3076 1840 3078 1844
rect 3070 1838 3078 1840
rect 3094 1844 3102 1846
rect 3094 1840 3096 1844
rect 3100 1840 3102 1844
rect 3094 1838 3102 1840
rect 3310 1844 3318 1846
rect 3310 1840 3312 1844
rect 3316 1840 3318 1844
rect 3310 1838 3318 1840
rect 3334 1844 3342 1846
rect 3334 1840 3336 1844
rect 3340 1840 3342 1844
rect 3334 1838 3342 1840
rect 3358 1844 3366 1846
rect 3358 1840 3360 1844
rect 3364 1840 3366 1844
rect 3358 1838 3366 1840
rect 3382 1844 3390 1846
rect 3382 1840 3384 1844
rect 3388 1840 3390 1844
rect 3382 1838 3390 1840
rect 3406 1844 3414 1846
rect 3406 1840 3408 1844
rect 3412 1840 3414 1844
rect 3406 1838 3414 1840
rect 3430 1844 3438 1846
rect 3430 1840 3432 1844
rect 3436 1840 3438 1844
rect 3430 1838 3438 1840
rect 3454 1844 3462 1846
rect 3454 1840 3456 1844
rect 3460 1840 3462 1844
rect 3454 1838 3462 1840
rect 3478 1844 3486 1846
rect 3478 1840 3480 1844
rect 3484 1840 3486 1844
rect 3478 1838 3486 1840
rect 3502 1844 3510 1846
rect 3502 1840 3504 1844
rect 3508 1840 3510 1844
rect 3502 1838 3510 1840
rect 3526 1844 3534 1846
rect 3526 1840 3528 1844
rect 3532 1840 3534 1844
rect 3526 1838 3534 1840
rect 3550 1844 3558 1846
rect 3550 1840 3552 1844
rect 3556 1840 3558 1844
rect 3550 1838 3558 1840
rect 3574 1844 3582 1846
rect 3574 1840 3576 1844
rect 3580 1840 3582 1844
rect 3574 1838 3582 1840
rect 3598 1844 3606 1846
rect 3598 1840 3600 1844
rect 3604 1840 3606 1844
rect 3598 1838 3606 1840
rect 3622 1844 3630 1846
rect 3622 1840 3624 1844
rect 3628 1840 3630 1844
rect 3622 1838 3630 1840
rect 3646 1844 3654 1846
rect 3646 1840 3648 1844
rect 3652 1840 3654 1844
rect 3646 1838 3654 1840
rect 3670 1844 3678 1846
rect 3670 1840 3672 1844
rect 3676 1840 3678 1844
rect 3670 1838 3678 1840
rect 3694 1844 3702 1846
rect 3694 1840 3696 1844
rect 3700 1840 3702 1844
rect 3694 1838 3702 1840
rect 3910 1844 3918 1846
rect 3910 1840 3912 1844
rect 3916 1840 3918 1844
rect 3910 1838 3918 1840
rect 3934 1844 3942 1846
rect 3934 1840 3936 1844
rect 3940 1840 3942 1844
rect 3934 1838 3942 1840
rect 3958 1844 3966 1846
rect 3958 1840 3960 1844
rect 3964 1840 3966 1844
rect 3958 1838 3966 1840
rect 3982 1844 3990 1846
rect 3982 1840 3984 1844
rect 3988 1840 3990 1844
rect 3982 1838 3990 1840
rect 4006 1844 4014 1846
rect 4006 1840 4008 1844
rect 4012 1840 4014 1844
rect 4006 1838 4014 1840
rect 4030 1844 4038 1846
rect 4030 1840 4032 1844
rect 4036 1840 4038 1844
rect 4030 1838 4038 1840
rect 4054 1844 4062 1846
rect 4054 1840 4056 1844
rect 4060 1840 4062 1844
rect 4054 1838 4062 1840
rect 4078 1844 4086 1846
rect 4078 1840 4080 1844
rect 4084 1840 4086 1844
rect 4078 1838 4086 1840
rect 4102 1844 4110 1846
rect 4102 1840 4104 1844
rect 4108 1840 4110 1844
rect 4102 1838 4110 1840
rect 4126 1844 4134 1846
rect 4126 1840 4128 1844
rect 4132 1840 4134 1844
rect 4126 1838 4134 1840
rect 4150 1844 4158 1846
rect 4150 1840 4152 1844
rect 4156 1840 4158 1844
rect 4150 1838 4158 1840
rect 4174 1844 4182 1846
rect 4174 1840 4176 1844
rect 4180 1840 4182 1844
rect 4174 1838 4182 1840
rect 4198 1844 4206 1846
rect 4198 1840 4200 1844
rect 4204 1840 4206 1844
rect 4198 1838 4206 1840
rect 4222 1844 4230 1846
rect 4222 1840 4224 1844
rect 4228 1840 4230 1844
rect 4222 1838 4230 1840
rect 4246 1844 4254 1846
rect 4246 1840 4248 1844
rect 4252 1840 4254 1844
rect 4246 1838 4254 1840
rect 4270 1844 4278 1846
rect 4270 1840 4272 1844
rect 4276 1840 4278 1844
rect 4270 1838 4278 1840
rect 4294 1844 4302 1846
rect 4294 1840 4296 1844
rect 4300 1840 4302 1844
rect 4294 1838 4302 1840
rect 4510 1844 4518 1846
rect 4510 1840 4512 1844
rect 4516 1840 4518 1844
rect 4510 1838 4518 1840
rect 4534 1844 4542 1846
rect 4534 1840 4536 1844
rect 4540 1840 4542 1844
rect 4534 1838 4542 1840
rect 4558 1844 4566 1846
rect 4558 1840 4560 1844
rect 4564 1840 4566 1844
rect 4558 1838 4566 1840
rect 4582 1844 4590 1846
rect 4582 1840 4584 1844
rect 4588 1840 4590 1844
rect 4582 1838 4590 1840
rect 4606 1844 4614 1846
rect 4606 1840 4608 1844
rect 4612 1840 4614 1844
rect 4606 1838 4614 1840
rect 4630 1844 4638 1846
rect 4630 1840 4632 1844
rect 4636 1840 4638 1844
rect 4630 1838 4638 1840
rect 4654 1844 4662 1846
rect 4654 1840 4656 1844
rect 4660 1840 4662 1844
rect 4654 1838 4662 1840
rect 4678 1844 4686 1846
rect 4678 1840 4680 1844
rect 4684 1840 4686 1844
rect 4678 1838 4686 1840
rect 4702 1844 4710 1846
rect 4702 1840 4704 1844
rect 4708 1840 4710 1844
rect 4702 1838 4710 1840
rect 4726 1844 4734 1846
rect 4726 1840 4728 1844
rect 4732 1840 4734 1844
rect 4726 1838 4734 1840
rect 4750 1844 4758 1846
rect 4750 1840 4752 1844
rect 4756 1840 4758 1844
rect 4750 1838 4758 1840
rect 4774 1844 4782 1846
rect 4774 1840 4776 1844
rect 4780 1840 4782 1844
rect 4774 1838 4782 1840
rect 4798 1838 4800 1846
rect 5710 1844 5718 1846
rect 5710 1840 5712 1844
rect 5716 1840 5718 1844
rect 5710 1838 5718 1840
rect 5734 1844 5742 1846
rect 5734 1840 5736 1844
rect 5740 1840 5742 1844
rect 5734 1838 5742 1840
rect 5758 1844 5766 1846
rect 5758 1840 5760 1844
rect 5764 1840 5766 1844
rect 5758 1838 5766 1840
rect 5782 1844 5790 1846
rect 5782 1840 5784 1844
rect 5788 1840 5790 1844
rect 5782 1838 5790 1840
rect 5806 1844 5814 1846
rect 5806 1840 5808 1844
rect 5812 1840 5814 1844
rect 5806 1838 5814 1840
rect 5830 1844 5838 1846
rect 5830 1840 5832 1844
rect 5836 1840 5838 1844
rect 5830 1838 5838 1840
rect 5854 1844 5862 1846
rect 5854 1840 5856 1844
rect 5860 1840 5862 1844
rect 5854 1838 5862 1840
rect 5878 1844 5886 1846
rect 5878 1840 5880 1844
rect 5884 1840 5886 1844
rect 5878 1838 5886 1840
rect 5902 1844 5910 1846
rect 5902 1840 5904 1844
rect 5908 1840 5910 1844
rect 5902 1838 5910 1840
rect 5926 1844 5934 1846
rect 5926 1840 5928 1844
rect 5932 1840 5934 1844
rect 5926 1838 5934 1840
rect 5950 1844 5958 1846
rect 5950 1840 5952 1844
rect 5956 1840 5958 1844
rect 5950 1838 5958 1840
rect 5974 1844 5982 1846
rect 5974 1840 5976 1844
rect 5980 1840 5982 1844
rect 5974 1838 5982 1840
rect 5998 1844 6006 1846
rect 5998 1840 6000 1844
rect 6004 1840 6006 1844
rect 5998 1838 6006 1840
rect 6022 1844 6030 1846
rect 6022 1840 6024 1844
rect 6028 1840 6030 1844
rect 6022 1838 6030 1840
rect 6046 1844 6054 1846
rect 6046 1840 6048 1844
rect 6052 1840 6054 1844
rect 6046 1838 6054 1840
rect 6070 1844 6078 1846
rect 6070 1840 6072 1844
rect 6076 1840 6078 1844
rect 6070 1838 6078 1840
rect 6094 1844 6102 1846
rect 6094 1840 6096 1844
rect 6100 1840 6102 1844
rect 6094 1838 6102 1840
rect 6310 1844 6318 1846
rect 6310 1840 6312 1844
rect 6316 1840 6318 1844
rect 6310 1838 6318 1840
rect 6334 1844 6342 1846
rect 6334 1840 6336 1844
rect 6340 1840 6342 1844
rect 6334 1838 6342 1840
rect 6358 1844 6366 1846
rect 6358 1840 6360 1844
rect 6364 1840 6366 1844
rect 6358 1838 6366 1840
rect 6382 1844 6390 1846
rect 6382 1840 6384 1844
rect 6388 1840 6390 1844
rect 6382 1838 6390 1840
rect 6406 1844 6414 1846
rect 6406 1840 6408 1844
rect 6412 1840 6414 1844
rect 6406 1838 6414 1840
rect 6430 1844 6438 1846
rect 6430 1840 6432 1844
rect 6436 1840 6438 1844
rect 6430 1838 6438 1840
rect 6454 1844 6462 1846
rect 6454 1840 6456 1844
rect 6460 1840 6462 1844
rect 6454 1838 6462 1840
rect 6478 1844 6486 1846
rect 6478 1840 6480 1844
rect 6484 1840 6486 1844
rect 6478 1838 6486 1840
rect 6502 1844 6510 1846
rect 6502 1840 6504 1844
rect 6508 1840 6510 1844
rect 6502 1838 6510 1840
rect 6526 1844 6534 1846
rect 6526 1840 6528 1844
rect 6532 1840 6534 1844
rect 6526 1838 6534 1840
rect 6550 1844 6558 1846
rect 6550 1840 6552 1844
rect 6556 1840 6558 1844
rect 6550 1838 6558 1840
rect 6574 1844 6582 1846
rect 6574 1840 6576 1844
rect 6580 1840 6582 1844
rect 6574 1838 6582 1840
rect 6598 1844 6606 1846
rect 6598 1840 6600 1844
rect 6604 1840 6606 1844
rect 6598 1838 6606 1840
rect 6622 1844 6630 1846
rect 6622 1840 6624 1844
rect 6628 1840 6630 1844
rect 6622 1838 6630 1840
rect 6646 1844 6654 1846
rect 6646 1840 6648 1844
rect 6652 1840 6654 1844
rect 6646 1838 6654 1840
rect 6670 1844 6678 1846
rect 6670 1840 6672 1844
rect 6676 1840 6678 1844
rect 6670 1838 6678 1840
rect 6694 1844 6702 1846
rect 6694 1840 6696 1844
rect 6700 1840 6702 1844
rect 6694 1838 6702 1840
rect 6910 1844 6918 1846
rect 6910 1840 6912 1844
rect 6916 1840 6918 1844
rect 6910 1838 6918 1840
rect 6934 1844 6942 1846
rect 6934 1840 6936 1844
rect 6940 1840 6942 1844
rect 6934 1838 6942 1840
rect 6958 1844 6966 1846
rect 6958 1840 6960 1844
rect 6964 1840 6966 1844
rect 6958 1838 6966 1840
rect 6982 1844 6990 1846
rect 6982 1840 6984 1844
rect 6988 1840 6990 1844
rect 6982 1838 6990 1840
rect 7006 1844 7014 1846
rect 7006 1840 7008 1844
rect 7012 1840 7014 1844
rect 7006 1838 7014 1840
rect 7030 1844 7038 1846
rect 7030 1840 7032 1844
rect 7036 1840 7038 1844
rect 7030 1838 7038 1840
rect 7054 1844 7062 1846
rect 7054 1840 7056 1844
rect 7060 1840 7062 1844
rect 7054 1838 7062 1840
rect 7078 1844 7086 1846
rect 7078 1840 7080 1844
rect 7084 1840 7086 1844
rect 7078 1838 7086 1840
rect 7102 1844 7110 1846
rect 7102 1840 7104 1844
rect 7108 1840 7110 1844
rect 7102 1838 7110 1840
rect 7126 1844 7134 1846
rect 7126 1840 7128 1844
rect 7132 1840 7134 1844
rect 7126 1838 7134 1840
rect 7150 1844 7158 1846
rect 7150 1840 7152 1844
rect 7156 1840 7158 1844
rect 7150 1838 7158 1840
rect 7174 1844 7182 1846
rect 7174 1840 7176 1844
rect 7180 1840 7182 1844
rect 7174 1838 7182 1840
rect 7198 1838 7200 1846
rect 2410 1832 2418 1834
rect 2410 1828 2412 1832
rect 2416 1828 2418 1832
rect 2410 1826 2418 1828
rect 2434 1832 2442 1834
rect 2434 1828 2436 1832
rect 2440 1828 2442 1832
rect 2434 1826 2442 1828
rect 2458 1832 2466 1834
rect 2458 1828 2460 1832
rect 2464 1828 2466 1832
rect 2458 1826 2466 1828
rect 2482 1832 2490 1834
rect 2482 1828 2484 1832
rect 2488 1828 2490 1832
rect 2482 1826 2490 1828
rect 2698 1832 2706 1834
rect 2698 1828 2700 1832
rect 2704 1828 2706 1832
rect 2698 1826 2706 1828
rect 2722 1832 2730 1834
rect 2722 1828 2724 1832
rect 2728 1828 2730 1832
rect 2722 1826 2730 1828
rect 2746 1832 2754 1834
rect 2746 1828 2748 1832
rect 2752 1828 2754 1832
rect 2746 1826 2754 1828
rect 2770 1832 2778 1834
rect 2770 1828 2772 1832
rect 2776 1828 2778 1832
rect 2770 1826 2778 1828
rect 2794 1832 2802 1834
rect 2794 1828 2796 1832
rect 2800 1828 2802 1832
rect 2794 1826 2802 1828
rect 2818 1832 2826 1834
rect 2818 1828 2820 1832
rect 2824 1828 2826 1832
rect 2818 1826 2826 1828
rect 2842 1832 2850 1834
rect 2842 1828 2844 1832
rect 2848 1828 2850 1832
rect 2842 1826 2850 1828
rect 2866 1832 2874 1834
rect 2866 1828 2868 1832
rect 2872 1828 2874 1832
rect 2866 1826 2874 1828
rect 2890 1832 2898 1834
rect 2890 1828 2892 1832
rect 2896 1828 2898 1832
rect 2890 1826 2898 1828
rect 2914 1832 2922 1834
rect 2914 1828 2916 1832
rect 2920 1828 2922 1832
rect 2914 1826 2922 1828
rect 2938 1832 2946 1834
rect 2938 1828 2940 1832
rect 2944 1828 2946 1832
rect 2938 1826 2946 1828
rect 2962 1832 2970 1834
rect 2962 1828 2964 1832
rect 2968 1828 2970 1832
rect 2962 1826 2970 1828
rect 2986 1832 2994 1834
rect 2986 1828 2988 1832
rect 2992 1828 2994 1832
rect 2986 1826 2994 1828
rect 3010 1832 3018 1834
rect 3010 1828 3012 1832
rect 3016 1828 3018 1832
rect 3010 1826 3018 1828
rect 3034 1832 3042 1834
rect 3034 1828 3036 1832
rect 3040 1828 3042 1832
rect 3034 1826 3042 1828
rect 3058 1832 3066 1834
rect 3058 1828 3060 1832
rect 3064 1828 3066 1832
rect 3058 1826 3066 1828
rect 3082 1832 3090 1834
rect 3082 1828 3084 1832
rect 3088 1828 3090 1832
rect 3082 1826 3090 1828
rect 3298 1832 3306 1834
rect 3298 1828 3300 1832
rect 3304 1828 3306 1832
rect 3298 1826 3306 1828
rect 3322 1832 3330 1834
rect 3322 1828 3324 1832
rect 3328 1828 3330 1832
rect 3322 1826 3330 1828
rect 3346 1832 3354 1834
rect 3346 1828 3348 1832
rect 3352 1828 3354 1832
rect 3346 1826 3354 1828
rect 3370 1832 3378 1834
rect 3370 1828 3372 1832
rect 3376 1828 3378 1832
rect 3370 1826 3378 1828
rect 3394 1832 3402 1834
rect 3394 1828 3396 1832
rect 3400 1828 3402 1832
rect 3394 1826 3402 1828
rect 3418 1832 3426 1834
rect 3418 1828 3420 1832
rect 3424 1828 3426 1832
rect 3418 1826 3426 1828
rect 3442 1832 3450 1834
rect 3442 1828 3444 1832
rect 3448 1828 3450 1832
rect 3442 1826 3450 1828
rect 3466 1832 3474 1834
rect 3466 1828 3468 1832
rect 3472 1828 3474 1832
rect 3466 1826 3474 1828
rect 3490 1832 3498 1834
rect 3490 1828 3492 1832
rect 3496 1828 3498 1832
rect 3490 1826 3498 1828
rect 3514 1832 3522 1834
rect 3514 1828 3516 1832
rect 3520 1828 3522 1832
rect 3514 1826 3522 1828
rect 3538 1832 3546 1834
rect 3538 1828 3540 1832
rect 3544 1828 3546 1832
rect 3538 1826 3546 1828
rect 3562 1832 3570 1834
rect 3562 1828 3564 1832
rect 3568 1828 3570 1832
rect 3562 1826 3570 1828
rect 3586 1832 3594 1834
rect 3586 1828 3588 1832
rect 3592 1828 3594 1832
rect 3586 1826 3594 1828
rect 3610 1832 3618 1834
rect 3610 1828 3612 1832
rect 3616 1828 3618 1832
rect 3610 1826 3618 1828
rect 3634 1832 3642 1834
rect 3634 1828 3636 1832
rect 3640 1828 3642 1832
rect 3634 1826 3642 1828
rect 3658 1832 3666 1834
rect 3658 1828 3660 1832
rect 3664 1828 3666 1832
rect 3658 1826 3666 1828
rect 3682 1832 3690 1834
rect 3682 1828 3684 1832
rect 3688 1828 3690 1832
rect 3682 1826 3690 1828
rect 3898 1832 3906 1834
rect 3898 1828 3900 1832
rect 3904 1828 3906 1832
rect 3898 1826 3906 1828
rect 3922 1832 3930 1834
rect 3922 1828 3924 1832
rect 3928 1828 3930 1832
rect 3922 1826 3930 1828
rect 3946 1832 3954 1834
rect 3946 1828 3948 1832
rect 3952 1828 3954 1832
rect 3946 1826 3954 1828
rect 3970 1832 3978 1834
rect 3970 1828 3972 1832
rect 3976 1828 3978 1832
rect 3970 1826 3978 1828
rect 3994 1832 4002 1834
rect 3994 1828 3996 1832
rect 4000 1828 4002 1832
rect 3994 1826 4002 1828
rect 4018 1832 4026 1834
rect 4018 1828 4020 1832
rect 4024 1828 4026 1832
rect 4018 1826 4026 1828
rect 4042 1832 4050 1834
rect 4042 1828 4044 1832
rect 4048 1828 4050 1832
rect 4042 1826 4050 1828
rect 4066 1832 4074 1834
rect 4066 1828 4068 1832
rect 4072 1828 4074 1832
rect 4066 1826 4074 1828
rect 4090 1832 4098 1834
rect 4090 1828 4092 1832
rect 4096 1828 4098 1832
rect 4090 1826 4098 1828
rect 4114 1832 4122 1834
rect 4114 1828 4116 1832
rect 4120 1828 4122 1832
rect 4114 1826 4122 1828
rect 4138 1832 4146 1834
rect 4138 1828 4140 1832
rect 4144 1828 4146 1832
rect 4138 1826 4146 1828
rect 4162 1832 4170 1834
rect 4162 1828 4164 1832
rect 4168 1828 4170 1832
rect 4162 1826 4170 1828
rect 4186 1832 4194 1834
rect 4186 1828 4188 1832
rect 4192 1828 4194 1832
rect 4186 1826 4194 1828
rect 4210 1832 4218 1834
rect 4210 1828 4212 1832
rect 4216 1828 4218 1832
rect 4210 1826 4218 1828
rect 4234 1832 4242 1834
rect 4234 1828 4236 1832
rect 4240 1828 4242 1832
rect 4234 1826 4242 1828
rect 4258 1832 4266 1834
rect 4258 1828 4260 1832
rect 4264 1828 4266 1832
rect 4258 1826 4266 1828
rect 4282 1832 4290 1834
rect 4282 1828 4284 1832
rect 4288 1828 4290 1832
rect 4282 1826 4290 1828
rect 4498 1832 4506 1834
rect 4498 1828 4500 1832
rect 4504 1828 4506 1832
rect 4498 1826 4506 1828
rect 4522 1832 4530 1834
rect 4522 1828 4524 1832
rect 4528 1828 4530 1832
rect 4522 1826 4530 1828
rect 4546 1832 4554 1834
rect 4546 1828 4548 1832
rect 4552 1828 4554 1832
rect 4546 1826 4554 1828
rect 4570 1832 4578 1834
rect 4570 1828 4572 1832
rect 4576 1828 4578 1832
rect 4570 1826 4578 1828
rect 4594 1832 4602 1834
rect 4594 1828 4596 1832
rect 4600 1828 4602 1832
rect 4594 1826 4602 1828
rect 4618 1832 4626 1834
rect 4618 1828 4620 1832
rect 4624 1828 4626 1832
rect 4618 1826 4626 1828
rect 4642 1832 4650 1834
rect 4642 1828 4644 1832
rect 4648 1828 4650 1832
rect 4642 1826 4650 1828
rect 4666 1832 4674 1834
rect 4666 1828 4668 1832
rect 4672 1828 4674 1832
rect 4666 1826 4674 1828
rect 4690 1832 4698 1834
rect 4690 1828 4692 1832
rect 4696 1828 4698 1832
rect 4690 1826 4698 1828
rect 4714 1832 4722 1834
rect 4714 1828 4716 1832
rect 4720 1828 4722 1832
rect 4714 1826 4722 1828
rect 4738 1832 4746 1834
rect 4738 1828 4740 1832
rect 4744 1828 4746 1832
rect 4738 1826 4746 1828
rect 4762 1832 4770 1834
rect 4762 1828 4764 1832
rect 4768 1828 4770 1832
rect 4762 1826 4770 1828
rect 4786 1832 4794 1834
rect 4786 1828 4788 1832
rect 4792 1828 4794 1832
rect 4786 1826 4794 1828
rect 5698 1832 5706 1834
rect 5698 1828 5700 1832
rect 5704 1828 5706 1832
rect 5698 1826 5706 1828
rect 5722 1832 5730 1834
rect 5722 1828 5724 1832
rect 5728 1828 5730 1832
rect 5722 1826 5730 1828
rect 5746 1832 5754 1834
rect 5746 1828 5748 1832
rect 5752 1828 5754 1832
rect 5746 1826 5754 1828
rect 5770 1832 5778 1834
rect 5770 1828 5772 1832
rect 5776 1828 5778 1832
rect 5770 1826 5778 1828
rect 5794 1832 5802 1834
rect 5794 1828 5796 1832
rect 5800 1828 5802 1832
rect 5794 1826 5802 1828
rect 5818 1832 5826 1834
rect 5818 1828 5820 1832
rect 5824 1828 5826 1832
rect 5818 1826 5826 1828
rect 5842 1832 5850 1834
rect 5842 1828 5844 1832
rect 5848 1828 5850 1832
rect 5842 1826 5850 1828
rect 5866 1832 5874 1834
rect 5866 1828 5868 1832
rect 5872 1828 5874 1832
rect 5866 1826 5874 1828
rect 5890 1832 5898 1834
rect 5890 1828 5892 1832
rect 5896 1828 5898 1832
rect 5890 1826 5898 1828
rect 5914 1832 5922 1834
rect 5914 1828 5916 1832
rect 5920 1828 5922 1832
rect 5914 1826 5922 1828
rect 5938 1832 5946 1834
rect 5938 1828 5940 1832
rect 5944 1828 5946 1832
rect 5938 1826 5946 1828
rect 5962 1832 5970 1834
rect 5962 1828 5964 1832
rect 5968 1828 5970 1832
rect 5962 1826 5970 1828
rect 5986 1832 5994 1834
rect 5986 1828 5988 1832
rect 5992 1828 5994 1832
rect 5986 1826 5994 1828
rect 6010 1832 6018 1834
rect 6010 1828 6012 1832
rect 6016 1828 6018 1832
rect 6010 1826 6018 1828
rect 6034 1832 6042 1834
rect 6034 1828 6036 1832
rect 6040 1828 6042 1832
rect 6034 1826 6042 1828
rect 6058 1832 6066 1834
rect 6058 1828 6060 1832
rect 6064 1828 6066 1832
rect 6058 1826 6066 1828
rect 6082 1832 6090 1834
rect 6082 1828 6084 1832
rect 6088 1828 6090 1832
rect 6082 1826 6090 1828
rect 6298 1832 6306 1834
rect 6298 1828 6300 1832
rect 6304 1828 6306 1832
rect 6298 1826 6306 1828
rect 6322 1832 6330 1834
rect 6322 1828 6324 1832
rect 6328 1828 6330 1832
rect 6322 1826 6330 1828
rect 6346 1832 6354 1834
rect 6346 1828 6348 1832
rect 6352 1828 6354 1832
rect 6346 1826 6354 1828
rect 6370 1832 6378 1834
rect 6370 1828 6372 1832
rect 6376 1828 6378 1832
rect 6370 1826 6378 1828
rect 6394 1832 6402 1834
rect 6394 1828 6396 1832
rect 6400 1828 6402 1832
rect 6394 1826 6402 1828
rect 6418 1832 6426 1834
rect 6418 1828 6420 1832
rect 6424 1828 6426 1832
rect 6418 1826 6426 1828
rect 6442 1832 6450 1834
rect 6442 1828 6444 1832
rect 6448 1828 6450 1832
rect 6442 1826 6450 1828
rect 6466 1832 6474 1834
rect 6466 1828 6468 1832
rect 6472 1828 6474 1832
rect 6466 1826 6474 1828
rect 6490 1832 6498 1834
rect 6490 1828 6492 1832
rect 6496 1828 6498 1832
rect 6490 1826 6498 1828
rect 6514 1832 6522 1834
rect 6514 1828 6516 1832
rect 6520 1828 6522 1832
rect 6514 1826 6522 1828
rect 6538 1832 6546 1834
rect 6538 1828 6540 1832
rect 6544 1828 6546 1832
rect 6538 1826 6546 1828
rect 6562 1832 6570 1834
rect 6562 1828 6564 1832
rect 6568 1828 6570 1832
rect 6562 1826 6570 1828
rect 6586 1832 6594 1834
rect 6586 1828 6588 1832
rect 6592 1828 6594 1832
rect 6586 1826 6594 1828
rect 6610 1832 6618 1834
rect 6610 1828 6612 1832
rect 6616 1828 6618 1832
rect 6610 1826 6618 1828
rect 6634 1832 6642 1834
rect 6634 1828 6636 1832
rect 6640 1828 6642 1832
rect 6634 1826 6642 1828
rect 6658 1832 6666 1834
rect 6658 1828 6660 1832
rect 6664 1828 6666 1832
rect 6658 1826 6666 1828
rect 6682 1832 6690 1834
rect 6682 1828 6684 1832
rect 6688 1828 6690 1832
rect 6682 1826 6690 1828
rect 6898 1832 6906 1834
rect 6898 1828 6900 1832
rect 6904 1828 6906 1832
rect 6898 1826 6906 1828
rect 6922 1832 6930 1834
rect 6922 1828 6924 1832
rect 6928 1828 6930 1832
rect 6922 1826 6930 1828
rect 6946 1832 6954 1834
rect 6946 1828 6948 1832
rect 6952 1828 6954 1832
rect 6946 1826 6954 1828
rect 6970 1832 6978 1834
rect 6970 1828 6972 1832
rect 6976 1828 6978 1832
rect 6970 1826 6978 1828
rect 6994 1832 7002 1834
rect 6994 1828 6996 1832
rect 7000 1828 7002 1832
rect 6994 1826 7002 1828
rect 7018 1832 7026 1834
rect 7018 1828 7020 1832
rect 7024 1828 7026 1832
rect 7018 1826 7026 1828
rect 7042 1832 7050 1834
rect 7042 1828 7044 1832
rect 7048 1828 7050 1832
rect 7042 1826 7050 1828
rect 7066 1832 7074 1834
rect 7066 1828 7068 1832
rect 7072 1828 7074 1832
rect 7066 1826 7074 1828
rect 7090 1832 7098 1834
rect 7090 1828 7092 1832
rect 7096 1828 7098 1832
rect 7090 1826 7098 1828
rect 7114 1832 7122 1834
rect 7114 1828 7116 1832
rect 7120 1828 7122 1832
rect 7114 1826 7122 1828
rect 7138 1832 7146 1834
rect 7138 1828 7140 1832
rect 7144 1828 7146 1832
rect 7138 1826 7146 1828
rect 7162 1832 7170 1834
rect 7162 1828 7164 1832
rect 7168 1828 7170 1832
rect 7162 1826 7170 1828
rect 7186 1832 7194 1834
rect 7186 1828 7188 1832
rect 7192 1828 7194 1832
rect 7186 1826 7194 1828
rect 2400 1820 2406 1822
rect 2404 1816 2406 1820
rect 2400 1814 2406 1816
rect 2422 1820 2430 1822
rect 2422 1816 2424 1820
rect 2428 1816 2430 1820
rect 2422 1814 2430 1816
rect 2446 1820 2454 1822
rect 2446 1816 2448 1820
rect 2452 1816 2454 1820
rect 2446 1814 2454 1816
rect 2470 1820 2478 1822
rect 2470 1816 2472 1820
rect 2476 1816 2478 1820
rect 2470 1814 2478 1816
rect 2494 1820 2502 1822
rect 2494 1816 2496 1820
rect 2500 1816 2502 1820
rect 2494 1814 2502 1816
rect 2710 1820 2718 1822
rect 2710 1816 2712 1820
rect 2716 1816 2718 1820
rect 2710 1814 2718 1816
rect 2734 1820 2742 1822
rect 2734 1816 2736 1820
rect 2740 1816 2742 1820
rect 2734 1814 2742 1816
rect 2758 1820 2766 1822
rect 2758 1816 2760 1820
rect 2764 1816 2766 1820
rect 2758 1814 2766 1816
rect 2782 1820 2790 1822
rect 2782 1816 2784 1820
rect 2788 1816 2790 1820
rect 2782 1814 2790 1816
rect 2806 1820 2814 1822
rect 2806 1816 2808 1820
rect 2812 1816 2814 1820
rect 2806 1814 2814 1816
rect 2830 1820 2838 1822
rect 2830 1816 2832 1820
rect 2836 1816 2838 1820
rect 2830 1814 2838 1816
rect 2854 1820 2862 1822
rect 2854 1816 2856 1820
rect 2860 1816 2862 1820
rect 2854 1814 2862 1816
rect 2878 1820 2886 1822
rect 2878 1816 2880 1820
rect 2884 1816 2886 1820
rect 2878 1814 2886 1816
rect 2902 1820 2910 1822
rect 2902 1816 2904 1820
rect 2908 1816 2910 1820
rect 2902 1814 2910 1816
rect 2926 1820 2934 1822
rect 2926 1816 2928 1820
rect 2932 1816 2934 1820
rect 2926 1814 2934 1816
rect 2950 1820 2958 1822
rect 2950 1816 2952 1820
rect 2956 1816 2958 1820
rect 2950 1814 2958 1816
rect 2974 1820 2982 1822
rect 2974 1816 2976 1820
rect 2980 1816 2982 1820
rect 2974 1814 2982 1816
rect 2998 1820 3006 1822
rect 2998 1816 3000 1820
rect 3004 1816 3006 1820
rect 2998 1814 3006 1816
rect 3022 1820 3030 1822
rect 3022 1816 3024 1820
rect 3028 1816 3030 1820
rect 3022 1814 3030 1816
rect 3046 1820 3054 1822
rect 3046 1816 3048 1820
rect 3052 1816 3054 1820
rect 3046 1814 3054 1816
rect 3070 1820 3078 1822
rect 3070 1816 3072 1820
rect 3076 1816 3078 1820
rect 3070 1814 3078 1816
rect 3094 1820 3102 1822
rect 3094 1816 3096 1820
rect 3100 1816 3102 1820
rect 3094 1814 3102 1816
rect 3310 1820 3318 1822
rect 3310 1816 3312 1820
rect 3316 1816 3318 1820
rect 3310 1814 3318 1816
rect 3334 1820 3342 1822
rect 3334 1816 3336 1820
rect 3340 1816 3342 1820
rect 3334 1814 3342 1816
rect 3358 1820 3366 1822
rect 3358 1816 3360 1820
rect 3364 1816 3366 1820
rect 3358 1814 3366 1816
rect 3382 1820 3390 1822
rect 3382 1816 3384 1820
rect 3388 1816 3390 1820
rect 3382 1814 3390 1816
rect 3406 1820 3414 1822
rect 3406 1816 3408 1820
rect 3412 1816 3414 1820
rect 3406 1814 3414 1816
rect 3430 1820 3438 1822
rect 3430 1816 3432 1820
rect 3436 1816 3438 1820
rect 3430 1814 3438 1816
rect 3454 1820 3462 1822
rect 3454 1816 3456 1820
rect 3460 1816 3462 1820
rect 3454 1814 3462 1816
rect 3478 1820 3486 1822
rect 3478 1816 3480 1820
rect 3484 1816 3486 1820
rect 3478 1814 3486 1816
rect 3502 1820 3510 1822
rect 3502 1816 3504 1820
rect 3508 1816 3510 1820
rect 3502 1814 3510 1816
rect 3526 1820 3534 1822
rect 3526 1816 3528 1820
rect 3532 1816 3534 1820
rect 3526 1814 3534 1816
rect 3550 1820 3558 1822
rect 3550 1816 3552 1820
rect 3556 1816 3558 1820
rect 3550 1814 3558 1816
rect 3574 1820 3582 1822
rect 3574 1816 3576 1820
rect 3580 1816 3582 1820
rect 3574 1814 3582 1816
rect 3598 1820 3606 1822
rect 3598 1816 3600 1820
rect 3604 1816 3606 1820
rect 3598 1814 3606 1816
rect 3622 1820 3630 1822
rect 3622 1816 3624 1820
rect 3628 1816 3630 1820
rect 3622 1814 3630 1816
rect 3646 1820 3654 1822
rect 3646 1816 3648 1820
rect 3652 1816 3654 1820
rect 3646 1814 3654 1816
rect 3670 1820 3678 1822
rect 3670 1816 3672 1820
rect 3676 1816 3678 1820
rect 3670 1814 3678 1816
rect 3694 1820 3702 1822
rect 3694 1816 3696 1820
rect 3700 1816 3702 1820
rect 3694 1814 3702 1816
rect 3910 1820 3918 1822
rect 3910 1816 3912 1820
rect 3916 1816 3918 1820
rect 3910 1814 3918 1816
rect 3934 1820 3942 1822
rect 3934 1816 3936 1820
rect 3940 1816 3942 1820
rect 3934 1814 3942 1816
rect 3958 1820 3966 1822
rect 3958 1816 3960 1820
rect 3964 1816 3966 1820
rect 3958 1814 3966 1816
rect 3982 1820 3990 1822
rect 3982 1816 3984 1820
rect 3988 1816 3990 1820
rect 3982 1814 3990 1816
rect 4006 1820 4014 1822
rect 4006 1816 4008 1820
rect 4012 1816 4014 1820
rect 4006 1814 4014 1816
rect 4030 1820 4038 1822
rect 4030 1816 4032 1820
rect 4036 1816 4038 1820
rect 4030 1814 4038 1816
rect 4054 1820 4062 1822
rect 4054 1816 4056 1820
rect 4060 1816 4062 1820
rect 4054 1814 4062 1816
rect 4078 1820 4086 1822
rect 4078 1816 4080 1820
rect 4084 1816 4086 1820
rect 4078 1814 4086 1816
rect 4102 1820 4110 1822
rect 4102 1816 4104 1820
rect 4108 1816 4110 1820
rect 4102 1814 4110 1816
rect 4126 1820 4134 1822
rect 4126 1816 4128 1820
rect 4132 1816 4134 1820
rect 4126 1814 4134 1816
rect 4150 1820 4158 1822
rect 4150 1816 4152 1820
rect 4156 1816 4158 1820
rect 4150 1814 4158 1816
rect 4174 1820 4182 1822
rect 4174 1816 4176 1820
rect 4180 1816 4182 1820
rect 4174 1814 4182 1816
rect 4198 1820 4206 1822
rect 4198 1816 4200 1820
rect 4204 1816 4206 1820
rect 4198 1814 4206 1816
rect 4222 1820 4230 1822
rect 4222 1816 4224 1820
rect 4228 1816 4230 1820
rect 4222 1814 4230 1816
rect 4246 1820 4254 1822
rect 4246 1816 4248 1820
rect 4252 1816 4254 1820
rect 4246 1814 4254 1816
rect 4270 1820 4278 1822
rect 4270 1816 4272 1820
rect 4276 1816 4278 1820
rect 4270 1814 4278 1816
rect 4294 1820 4302 1822
rect 4294 1816 4296 1820
rect 4300 1816 4302 1820
rect 4294 1814 4302 1816
rect 4510 1820 4518 1822
rect 4510 1816 4512 1820
rect 4516 1816 4518 1820
rect 4510 1814 4518 1816
rect 4534 1820 4542 1822
rect 4534 1816 4536 1820
rect 4540 1816 4542 1820
rect 4534 1814 4542 1816
rect 4558 1820 4566 1822
rect 4558 1816 4560 1820
rect 4564 1816 4566 1820
rect 4558 1814 4566 1816
rect 4582 1820 4590 1822
rect 4582 1816 4584 1820
rect 4588 1816 4590 1820
rect 4582 1814 4590 1816
rect 4606 1820 4614 1822
rect 4606 1816 4608 1820
rect 4612 1816 4614 1820
rect 4606 1814 4614 1816
rect 4630 1820 4638 1822
rect 4630 1816 4632 1820
rect 4636 1816 4638 1820
rect 4630 1814 4638 1816
rect 4654 1820 4662 1822
rect 4654 1816 4656 1820
rect 4660 1816 4662 1820
rect 4654 1814 4662 1816
rect 4678 1820 4686 1822
rect 4678 1816 4680 1820
rect 4684 1816 4686 1820
rect 4678 1814 4686 1816
rect 4702 1820 4710 1822
rect 4702 1816 4704 1820
rect 4708 1816 4710 1820
rect 4702 1814 4710 1816
rect 4726 1820 4734 1822
rect 4726 1816 4728 1820
rect 4732 1816 4734 1820
rect 4726 1814 4734 1816
rect 4750 1820 4758 1822
rect 4750 1816 4752 1820
rect 4756 1816 4758 1820
rect 4750 1814 4758 1816
rect 4774 1820 4782 1822
rect 4774 1816 4776 1820
rect 4780 1816 4782 1820
rect 4774 1814 4782 1816
rect 4798 1814 4800 1822
rect 5710 1820 5718 1822
rect 5710 1816 5712 1820
rect 5716 1816 5718 1820
rect 5710 1814 5718 1816
rect 5734 1820 5742 1822
rect 5734 1816 5736 1820
rect 5740 1816 5742 1820
rect 5734 1814 5742 1816
rect 5758 1820 5766 1822
rect 5758 1816 5760 1820
rect 5764 1816 5766 1820
rect 5758 1814 5766 1816
rect 5782 1820 5790 1822
rect 5782 1816 5784 1820
rect 5788 1816 5790 1820
rect 5782 1814 5790 1816
rect 5806 1820 5814 1822
rect 5806 1816 5808 1820
rect 5812 1816 5814 1820
rect 5806 1814 5814 1816
rect 5830 1820 5838 1822
rect 5830 1816 5832 1820
rect 5836 1816 5838 1820
rect 5830 1814 5838 1816
rect 5854 1820 5862 1822
rect 5854 1816 5856 1820
rect 5860 1816 5862 1820
rect 5854 1814 5862 1816
rect 5878 1820 5886 1822
rect 5878 1816 5880 1820
rect 5884 1816 5886 1820
rect 5878 1814 5886 1816
rect 5902 1820 5910 1822
rect 5902 1816 5904 1820
rect 5908 1816 5910 1820
rect 5902 1814 5910 1816
rect 5926 1820 5934 1822
rect 5926 1816 5928 1820
rect 5932 1816 5934 1820
rect 5926 1814 5934 1816
rect 5950 1820 5958 1822
rect 5950 1816 5952 1820
rect 5956 1816 5958 1820
rect 5950 1814 5958 1816
rect 5974 1820 5982 1822
rect 5974 1816 5976 1820
rect 5980 1816 5982 1820
rect 5974 1814 5982 1816
rect 5998 1820 6006 1822
rect 5998 1816 6000 1820
rect 6004 1816 6006 1820
rect 5998 1814 6006 1816
rect 6022 1820 6030 1822
rect 6022 1816 6024 1820
rect 6028 1816 6030 1820
rect 6022 1814 6030 1816
rect 6046 1820 6054 1822
rect 6046 1816 6048 1820
rect 6052 1816 6054 1820
rect 6046 1814 6054 1816
rect 6070 1820 6078 1822
rect 6070 1816 6072 1820
rect 6076 1816 6078 1820
rect 6070 1814 6078 1816
rect 6094 1820 6102 1822
rect 6094 1816 6096 1820
rect 6100 1816 6102 1820
rect 6094 1814 6102 1816
rect 6310 1820 6318 1822
rect 6310 1816 6312 1820
rect 6316 1816 6318 1820
rect 6310 1814 6318 1816
rect 6334 1820 6342 1822
rect 6334 1816 6336 1820
rect 6340 1816 6342 1820
rect 6334 1814 6342 1816
rect 6358 1820 6366 1822
rect 6358 1816 6360 1820
rect 6364 1816 6366 1820
rect 6358 1814 6366 1816
rect 6382 1820 6390 1822
rect 6382 1816 6384 1820
rect 6388 1816 6390 1820
rect 6382 1814 6390 1816
rect 6406 1820 6414 1822
rect 6406 1816 6408 1820
rect 6412 1816 6414 1820
rect 6406 1814 6414 1816
rect 6430 1820 6438 1822
rect 6430 1816 6432 1820
rect 6436 1816 6438 1820
rect 6430 1814 6438 1816
rect 6454 1820 6462 1822
rect 6454 1816 6456 1820
rect 6460 1816 6462 1820
rect 6454 1814 6462 1816
rect 6478 1820 6486 1822
rect 6478 1816 6480 1820
rect 6484 1816 6486 1820
rect 6478 1814 6486 1816
rect 6502 1820 6510 1822
rect 6502 1816 6504 1820
rect 6508 1816 6510 1820
rect 6502 1814 6510 1816
rect 6526 1820 6534 1822
rect 6526 1816 6528 1820
rect 6532 1816 6534 1820
rect 6526 1814 6534 1816
rect 6550 1820 6558 1822
rect 6550 1816 6552 1820
rect 6556 1816 6558 1820
rect 6550 1814 6558 1816
rect 6574 1820 6582 1822
rect 6574 1816 6576 1820
rect 6580 1816 6582 1820
rect 6574 1814 6582 1816
rect 6598 1820 6606 1822
rect 6598 1816 6600 1820
rect 6604 1816 6606 1820
rect 6598 1814 6606 1816
rect 6622 1820 6630 1822
rect 6622 1816 6624 1820
rect 6628 1816 6630 1820
rect 6622 1814 6630 1816
rect 6646 1820 6654 1822
rect 6646 1816 6648 1820
rect 6652 1816 6654 1820
rect 6646 1814 6654 1816
rect 6670 1820 6678 1822
rect 6670 1816 6672 1820
rect 6676 1816 6678 1820
rect 6670 1814 6678 1816
rect 6694 1820 6702 1822
rect 6694 1816 6696 1820
rect 6700 1816 6702 1820
rect 6694 1814 6702 1816
rect 6910 1820 6918 1822
rect 6910 1816 6912 1820
rect 6916 1816 6918 1820
rect 6910 1814 6918 1816
rect 6934 1820 6942 1822
rect 6934 1816 6936 1820
rect 6940 1816 6942 1820
rect 6934 1814 6942 1816
rect 6958 1820 6966 1822
rect 6958 1816 6960 1820
rect 6964 1816 6966 1820
rect 6958 1814 6966 1816
rect 6982 1820 6990 1822
rect 6982 1816 6984 1820
rect 6988 1816 6990 1820
rect 6982 1814 6990 1816
rect 7006 1820 7014 1822
rect 7006 1816 7008 1820
rect 7012 1816 7014 1820
rect 7006 1814 7014 1816
rect 7030 1820 7038 1822
rect 7030 1816 7032 1820
rect 7036 1816 7038 1820
rect 7030 1814 7038 1816
rect 7054 1820 7062 1822
rect 7054 1816 7056 1820
rect 7060 1816 7062 1820
rect 7054 1814 7062 1816
rect 7078 1820 7086 1822
rect 7078 1816 7080 1820
rect 7084 1816 7086 1820
rect 7078 1814 7086 1816
rect 7102 1820 7110 1822
rect 7102 1816 7104 1820
rect 7108 1816 7110 1820
rect 7102 1814 7110 1816
rect 7126 1820 7134 1822
rect 7126 1816 7128 1820
rect 7132 1816 7134 1820
rect 7126 1814 7134 1816
rect 7150 1820 7158 1822
rect 7150 1816 7152 1820
rect 7156 1816 7158 1820
rect 7150 1814 7158 1816
rect 7174 1820 7182 1822
rect 7174 1816 7176 1820
rect 7180 1816 7182 1820
rect 7174 1814 7182 1816
rect 7198 1814 7200 1822
rect 2410 1808 2418 1810
rect 2410 1804 2412 1808
rect 2416 1804 2418 1808
rect 2410 1802 2418 1804
rect 2434 1808 2442 1810
rect 2434 1804 2436 1808
rect 2440 1804 2442 1808
rect 2434 1802 2442 1804
rect 2458 1808 2466 1810
rect 2458 1804 2460 1808
rect 2464 1804 2466 1808
rect 2458 1802 2466 1804
rect 2482 1808 2490 1810
rect 2482 1804 2484 1808
rect 2488 1804 2490 1808
rect 2482 1802 2490 1804
rect 2698 1808 2706 1810
rect 2698 1804 2700 1808
rect 2704 1804 2706 1808
rect 2698 1802 2706 1804
rect 2722 1808 2730 1810
rect 2722 1804 2724 1808
rect 2728 1804 2730 1808
rect 2722 1802 2730 1804
rect 2746 1808 2754 1810
rect 2746 1804 2748 1808
rect 2752 1804 2754 1808
rect 2746 1802 2754 1804
rect 2770 1808 2778 1810
rect 2770 1804 2772 1808
rect 2776 1804 2778 1808
rect 2770 1802 2778 1804
rect 2794 1808 2802 1810
rect 2794 1804 2796 1808
rect 2800 1804 2802 1808
rect 2794 1802 2802 1804
rect 2818 1808 2826 1810
rect 2818 1804 2820 1808
rect 2824 1804 2826 1808
rect 2818 1802 2826 1804
rect 2842 1808 2850 1810
rect 2842 1804 2844 1808
rect 2848 1804 2850 1808
rect 2842 1802 2850 1804
rect 2866 1808 2874 1810
rect 2866 1804 2868 1808
rect 2872 1804 2874 1808
rect 2866 1802 2874 1804
rect 2890 1808 2898 1810
rect 2890 1804 2892 1808
rect 2896 1804 2898 1808
rect 2890 1802 2898 1804
rect 2914 1808 2922 1810
rect 2914 1804 2916 1808
rect 2920 1804 2922 1808
rect 2914 1802 2922 1804
rect 2938 1808 2946 1810
rect 2938 1804 2940 1808
rect 2944 1804 2946 1808
rect 2938 1802 2946 1804
rect 2962 1808 2970 1810
rect 2962 1804 2964 1808
rect 2968 1804 2970 1808
rect 2962 1802 2970 1804
rect 2986 1808 2994 1810
rect 2986 1804 2988 1808
rect 2992 1804 2994 1808
rect 2986 1802 2994 1804
rect 3010 1808 3018 1810
rect 3010 1804 3012 1808
rect 3016 1804 3018 1808
rect 3010 1802 3018 1804
rect 3034 1808 3042 1810
rect 3034 1804 3036 1808
rect 3040 1804 3042 1808
rect 3034 1802 3042 1804
rect 3058 1808 3066 1810
rect 3058 1804 3060 1808
rect 3064 1804 3066 1808
rect 3058 1802 3066 1804
rect 3082 1808 3090 1810
rect 3082 1804 3084 1808
rect 3088 1804 3090 1808
rect 3082 1802 3090 1804
rect 3298 1808 3306 1810
rect 3298 1804 3300 1808
rect 3304 1804 3306 1808
rect 3298 1802 3306 1804
rect 3322 1808 3330 1810
rect 3322 1804 3324 1808
rect 3328 1804 3330 1808
rect 3322 1802 3330 1804
rect 3346 1808 3354 1810
rect 3346 1804 3348 1808
rect 3352 1804 3354 1808
rect 3346 1802 3354 1804
rect 3370 1808 3378 1810
rect 3370 1804 3372 1808
rect 3376 1804 3378 1808
rect 3370 1802 3378 1804
rect 3394 1808 3402 1810
rect 3394 1804 3396 1808
rect 3400 1804 3402 1808
rect 3394 1802 3402 1804
rect 3418 1808 3426 1810
rect 3418 1804 3420 1808
rect 3424 1804 3426 1808
rect 3418 1802 3426 1804
rect 3442 1808 3450 1810
rect 3442 1804 3444 1808
rect 3448 1804 3450 1808
rect 3442 1802 3450 1804
rect 3466 1808 3474 1810
rect 3466 1804 3468 1808
rect 3472 1804 3474 1808
rect 3466 1802 3474 1804
rect 3490 1808 3498 1810
rect 3490 1804 3492 1808
rect 3496 1804 3498 1808
rect 3490 1802 3498 1804
rect 3514 1808 3522 1810
rect 3514 1804 3516 1808
rect 3520 1804 3522 1808
rect 3514 1802 3522 1804
rect 3538 1808 3546 1810
rect 3538 1804 3540 1808
rect 3544 1804 3546 1808
rect 3538 1802 3546 1804
rect 3562 1808 3570 1810
rect 3562 1804 3564 1808
rect 3568 1804 3570 1808
rect 3562 1802 3570 1804
rect 3586 1808 3594 1810
rect 3586 1804 3588 1808
rect 3592 1804 3594 1808
rect 3586 1802 3594 1804
rect 3610 1808 3618 1810
rect 3610 1804 3612 1808
rect 3616 1804 3618 1808
rect 3610 1802 3618 1804
rect 3634 1808 3642 1810
rect 3634 1804 3636 1808
rect 3640 1804 3642 1808
rect 3634 1802 3642 1804
rect 3658 1808 3666 1810
rect 3658 1804 3660 1808
rect 3664 1804 3666 1808
rect 3658 1802 3666 1804
rect 3682 1808 3690 1810
rect 3682 1804 3684 1808
rect 3688 1804 3690 1808
rect 3682 1802 3690 1804
rect 3898 1808 3906 1810
rect 3898 1804 3900 1808
rect 3904 1804 3906 1808
rect 3898 1802 3906 1804
rect 3922 1808 3930 1810
rect 3922 1804 3924 1808
rect 3928 1804 3930 1808
rect 3922 1802 3930 1804
rect 3946 1808 3954 1810
rect 3946 1804 3948 1808
rect 3952 1804 3954 1808
rect 3946 1802 3954 1804
rect 3970 1808 3978 1810
rect 3970 1804 3972 1808
rect 3976 1804 3978 1808
rect 3970 1802 3978 1804
rect 3994 1808 4002 1810
rect 3994 1804 3996 1808
rect 4000 1804 4002 1808
rect 3994 1802 4002 1804
rect 4018 1808 4026 1810
rect 4018 1804 4020 1808
rect 4024 1804 4026 1808
rect 4018 1802 4026 1804
rect 4042 1808 4050 1810
rect 4042 1804 4044 1808
rect 4048 1804 4050 1808
rect 4042 1802 4050 1804
rect 4066 1808 4074 1810
rect 4066 1804 4068 1808
rect 4072 1804 4074 1808
rect 4066 1802 4074 1804
rect 4090 1808 4098 1810
rect 4090 1804 4092 1808
rect 4096 1804 4098 1808
rect 4090 1802 4098 1804
rect 4114 1808 4122 1810
rect 4114 1804 4116 1808
rect 4120 1804 4122 1808
rect 4114 1802 4122 1804
rect 4138 1808 4146 1810
rect 4138 1804 4140 1808
rect 4144 1804 4146 1808
rect 4138 1802 4146 1804
rect 4162 1808 4170 1810
rect 4162 1804 4164 1808
rect 4168 1804 4170 1808
rect 4162 1802 4170 1804
rect 4186 1808 4194 1810
rect 4186 1804 4188 1808
rect 4192 1804 4194 1808
rect 4186 1802 4194 1804
rect 4210 1808 4218 1810
rect 4210 1804 4212 1808
rect 4216 1804 4218 1808
rect 4210 1802 4218 1804
rect 4234 1808 4242 1810
rect 4234 1804 4236 1808
rect 4240 1804 4242 1808
rect 4234 1802 4242 1804
rect 4258 1808 4266 1810
rect 4258 1804 4260 1808
rect 4264 1804 4266 1808
rect 4258 1802 4266 1804
rect 4282 1808 4290 1810
rect 4282 1804 4284 1808
rect 4288 1804 4290 1808
rect 4282 1802 4290 1804
rect 4498 1808 4506 1810
rect 4498 1804 4500 1808
rect 4504 1804 4506 1808
rect 4498 1802 4506 1804
rect 4522 1808 4530 1810
rect 4522 1804 4524 1808
rect 4528 1804 4530 1808
rect 4522 1802 4530 1804
rect 4546 1808 4554 1810
rect 4546 1804 4548 1808
rect 4552 1804 4554 1808
rect 4546 1802 4554 1804
rect 4570 1808 4578 1810
rect 4570 1804 4572 1808
rect 4576 1804 4578 1808
rect 4570 1802 4578 1804
rect 4594 1808 4602 1810
rect 4594 1804 4596 1808
rect 4600 1804 4602 1808
rect 4594 1802 4602 1804
rect 4618 1808 4626 1810
rect 4618 1804 4620 1808
rect 4624 1804 4626 1808
rect 4618 1802 4626 1804
rect 4642 1808 4650 1810
rect 4642 1804 4644 1808
rect 4648 1804 4650 1808
rect 4642 1802 4650 1804
rect 4666 1808 4674 1810
rect 4666 1804 4668 1808
rect 4672 1804 4674 1808
rect 4666 1802 4674 1804
rect 4690 1808 4698 1810
rect 4690 1804 4692 1808
rect 4696 1804 4698 1808
rect 4690 1802 4698 1804
rect 4714 1808 4722 1810
rect 4714 1804 4716 1808
rect 4720 1804 4722 1808
rect 4714 1802 4722 1804
rect 4738 1808 4746 1810
rect 4738 1804 4740 1808
rect 4744 1804 4746 1808
rect 4738 1802 4746 1804
rect 4762 1808 4770 1810
rect 4762 1804 4764 1808
rect 4768 1804 4770 1808
rect 4762 1802 4770 1804
rect 4786 1808 4794 1810
rect 4786 1804 4788 1808
rect 4792 1804 4794 1808
rect 4786 1802 4794 1804
rect 5698 1808 5706 1810
rect 5698 1804 5700 1808
rect 5704 1804 5706 1808
rect 5698 1802 5706 1804
rect 5722 1808 5730 1810
rect 5722 1804 5724 1808
rect 5728 1804 5730 1808
rect 5722 1802 5730 1804
rect 5746 1808 5754 1810
rect 5746 1804 5748 1808
rect 5752 1804 5754 1808
rect 5746 1802 5754 1804
rect 5770 1808 5778 1810
rect 5770 1804 5772 1808
rect 5776 1804 5778 1808
rect 5770 1802 5778 1804
rect 5794 1808 5802 1810
rect 5794 1804 5796 1808
rect 5800 1804 5802 1808
rect 5794 1802 5802 1804
rect 5818 1808 5826 1810
rect 5818 1804 5820 1808
rect 5824 1804 5826 1808
rect 5818 1802 5826 1804
rect 5842 1808 5850 1810
rect 5842 1804 5844 1808
rect 5848 1804 5850 1808
rect 5842 1802 5850 1804
rect 5866 1808 5874 1810
rect 5866 1804 5868 1808
rect 5872 1804 5874 1808
rect 5866 1802 5874 1804
rect 5890 1808 5898 1810
rect 5890 1804 5892 1808
rect 5896 1804 5898 1808
rect 5890 1802 5898 1804
rect 5914 1808 5922 1810
rect 5914 1804 5916 1808
rect 5920 1804 5922 1808
rect 5914 1802 5922 1804
rect 5938 1808 5946 1810
rect 5938 1804 5940 1808
rect 5944 1804 5946 1808
rect 5938 1802 5946 1804
rect 5962 1808 5970 1810
rect 5962 1804 5964 1808
rect 5968 1804 5970 1808
rect 5962 1802 5970 1804
rect 5986 1808 5994 1810
rect 5986 1804 5988 1808
rect 5992 1804 5994 1808
rect 5986 1802 5994 1804
rect 6010 1808 6018 1810
rect 6010 1804 6012 1808
rect 6016 1804 6018 1808
rect 6010 1802 6018 1804
rect 6034 1808 6042 1810
rect 6034 1804 6036 1808
rect 6040 1804 6042 1808
rect 6034 1802 6042 1804
rect 6058 1808 6066 1810
rect 6058 1804 6060 1808
rect 6064 1804 6066 1808
rect 6058 1802 6066 1804
rect 6082 1808 6090 1810
rect 6082 1804 6084 1808
rect 6088 1804 6090 1808
rect 6082 1802 6090 1804
rect 6298 1808 6306 1810
rect 6298 1804 6300 1808
rect 6304 1804 6306 1808
rect 6298 1802 6306 1804
rect 6322 1808 6330 1810
rect 6322 1804 6324 1808
rect 6328 1804 6330 1808
rect 6322 1802 6330 1804
rect 6346 1808 6354 1810
rect 6346 1804 6348 1808
rect 6352 1804 6354 1808
rect 6346 1802 6354 1804
rect 6370 1808 6378 1810
rect 6370 1804 6372 1808
rect 6376 1804 6378 1808
rect 6370 1802 6378 1804
rect 6394 1808 6402 1810
rect 6394 1804 6396 1808
rect 6400 1804 6402 1808
rect 6394 1802 6402 1804
rect 6418 1808 6426 1810
rect 6418 1804 6420 1808
rect 6424 1804 6426 1808
rect 6418 1802 6426 1804
rect 6442 1808 6450 1810
rect 6442 1804 6444 1808
rect 6448 1804 6450 1808
rect 6442 1802 6450 1804
rect 6466 1808 6474 1810
rect 6466 1804 6468 1808
rect 6472 1804 6474 1808
rect 6466 1802 6474 1804
rect 6490 1808 6498 1810
rect 6490 1804 6492 1808
rect 6496 1804 6498 1808
rect 6490 1802 6498 1804
rect 6514 1808 6522 1810
rect 6514 1804 6516 1808
rect 6520 1804 6522 1808
rect 6514 1802 6522 1804
rect 6538 1808 6546 1810
rect 6538 1804 6540 1808
rect 6544 1804 6546 1808
rect 6538 1802 6546 1804
rect 6562 1808 6570 1810
rect 6562 1804 6564 1808
rect 6568 1804 6570 1808
rect 6562 1802 6570 1804
rect 6586 1808 6594 1810
rect 6586 1804 6588 1808
rect 6592 1804 6594 1808
rect 6586 1802 6594 1804
rect 6610 1808 6618 1810
rect 6610 1804 6612 1808
rect 6616 1804 6618 1808
rect 6610 1802 6618 1804
rect 6634 1808 6642 1810
rect 6634 1804 6636 1808
rect 6640 1804 6642 1808
rect 6634 1802 6642 1804
rect 6658 1808 6666 1810
rect 6658 1804 6660 1808
rect 6664 1804 6666 1808
rect 6658 1802 6666 1804
rect 6682 1808 6690 1810
rect 6682 1804 6684 1808
rect 6688 1804 6690 1808
rect 6682 1802 6690 1804
rect 6898 1808 6906 1810
rect 6898 1804 6900 1808
rect 6904 1804 6906 1808
rect 6898 1802 6906 1804
rect 6922 1808 6930 1810
rect 6922 1804 6924 1808
rect 6928 1804 6930 1808
rect 6922 1802 6930 1804
rect 6946 1808 6954 1810
rect 6946 1804 6948 1808
rect 6952 1804 6954 1808
rect 6946 1802 6954 1804
rect 6970 1808 6978 1810
rect 6970 1804 6972 1808
rect 6976 1804 6978 1808
rect 6970 1802 6978 1804
rect 6994 1808 7002 1810
rect 6994 1804 6996 1808
rect 7000 1804 7002 1808
rect 6994 1802 7002 1804
rect 7018 1808 7026 1810
rect 7018 1804 7020 1808
rect 7024 1804 7026 1808
rect 7018 1802 7026 1804
rect 7042 1808 7050 1810
rect 7042 1804 7044 1808
rect 7048 1804 7050 1808
rect 7042 1802 7050 1804
rect 7066 1808 7074 1810
rect 7066 1804 7068 1808
rect 7072 1804 7074 1808
rect 7066 1802 7074 1804
rect 7090 1808 7098 1810
rect 7090 1804 7092 1808
rect 7096 1804 7098 1808
rect 7090 1802 7098 1804
rect 7114 1808 7122 1810
rect 7114 1804 7116 1808
rect 7120 1804 7122 1808
rect 7114 1802 7122 1804
rect 7138 1808 7146 1810
rect 7138 1804 7140 1808
rect 7144 1804 7146 1808
rect 7138 1802 7146 1804
rect 7162 1808 7170 1810
rect 7162 1804 7164 1808
rect 7168 1804 7170 1808
rect 7162 1802 7170 1804
rect 7186 1808 7194 1810
rect 7186 1804 7188 1808
rect 7192 1804 7194 1808
rect 7186 1802 7194 1804
rect 2400 1796 2406 1798
rect 2404 1792 2406 1796
rect 2400 1790 2406 1792
rect 2422 1796 2430 1798
rect 2422 1792 2424 1796
rect 2428 1792 2430 1796
rect 2422 1790 2430 1792
rect 2446 1796 2454 1798
rect 2446 1792 2448 1796
rect 2452 1792 2454 1796
rect 2446 1790 2454 1792
rect 2470 1796 2478 1798
rect 2470 1792 2472 1796
rect 2476 1792 2478 1796
rect 2470 1790 2478 1792
rect 2494 1796 2502 1798
rect 2494 1792 2496 1796
rect 2500 1792 2502 1796
rect 2494 1790 2502 1792
rect 2710 1796 2718 1798
rect 2710 1792 2712 1796
rect 2716 1792 2718 1796
rect 2710 1790 2718 1792
rect 2734 1796 2742 1798
rect 2734 1792 2736 1796
rect 2740 1792 2742 1796
rect 2734 1790 2742 1792
rect 2758 1796 2766 1798
rect 2758 1792 2760 1796
rect 2764 1792 2766 1796
rect 2758 1790 2766 1792
rect 2782 1796 2790 1798
rect 2782 1792 2784 1796
rect 2788 1792 2790 1796
rect 2782 1790 2790 1792
rect 2806 1796 2814 1798
rect 2806 1792 2808 1796
rect 2812 1792 2814 1796
rect 2806 1790 2814 1792
rect 2830 1796 2838 1798
rect 2830 1792 2832 1796
rect 2836 1792 2838 1796
rect 2830 1790 2838 1792
rect 2854 1796 2862 1798
rect 2854 1792 2856 1796
rect 2860 1792 2862 1796
rect 2854 1790 2862 1792
rect 2878 1796 2886 1798
rect 2878 1792 2880 1796
rect 2884 1792 2886 1796
rect 2878 1790 2886 1792
rect 2902 1796 2910 1798
rect 2902 1792 2904 1796
rect 2908 1792 2910 1796
rect 2902 1790 2910 1792
rect 2926 1796 2934 1798
rect 2926 1792 2928 1796
rect 2932 1792 2934 1796
rect 2926 1790 2934 1792
rect 2950 1796 2958 1798
rect 2950 1792 2952 1796
rect 2956 1792 2958 1796
rect 2950 1790 2958 1792
rect 2974 1796 2982 1798
rect 2974 1792 2976 1796
rect 2980 1792 2982 1796
rect 2974 1790 2982 1792
rect 2998 1796 3006 1798
rect 2998 1792 3000 1796
rect 3004 1792 3006 1796
rect 2998 1790 3006 1792
rect 3022 1796 3030 1798
rect 3022 1792 3024 1796
rect 3028 1792 3030 1796
rect 3022 1790 3030 1792
rect 3046 1796 3054 1798
rect 3046 1792 3048 1796
rect 3052 1792 3054 1796
rect 3046 1790 3054 1792
rect 3070 1796 3078 1798
rect 3070 1792 3072 1796
rect 3076 1792 3078 1796
rect 3070 1790 3078 1792
rect 3094 1796 3102 1798
rect 3094 1792 3096 1796
rect 3100 1792 3102 1796
rect 3094 1790 3102 1792
rect 3310 1796 3318 1798
rect 3310 1792 3312 1796
rect 3316 1792 3318 1796
rect 3310 1790 3318 1792
rect 3334 1796 3342 1798
rect 3334 1792 3336 1796
rect 3340 1792 3342 1796
rect 3334 1790 3342 1792
rect 3358 1796 3366 1798
rect 3358 1792 3360 1796
rect 3364 1792 3366 1796
rect 3358 1790 3366 1792
rect 3382 1796 3390 1798
rect 3382 1792 3384 1796
rect 3388 1792 3390 1796
rect 3382 1790 3390 1792
rect 3406 1796 3414 1798
rect 3406 1792 3408 1796
rect 3412 1792 3414 1796
rect 3406 1790 3414 1792
rect 3430 1796 3438 1798
rect 3430 1792 3432 1796
rect 3436 1792 3438 1796
rect 3430 1790 3438 1792
rect 3454 1796 3462 1798
rect 3454 1792 3456 1796
rect 3460 1792 3462 1796
rect 3454 1790 3462 1792
rect 3478 1796 3486 1798
rect 3478 1792 3480 1796
rect 3484 1792 3486 1796
rect 3478 1790 3486 1792
rect 3502 1796 3510 1798
rect 3502 1792 3504 1796
rect 3508 1792 3510 1796
rect 3502 1790 3510 1792
rect 3526 1796 3534 1798
rect 3526 1792 3528 1796
rect 3532 1792 3534 1796
rect 3526 1790 3534 1792
rect 3550 1796 3558 1798
rect 3550 1792 3552 1796
rect 3556 1792 3558 1796
rect 3550 1790 3558 1792
rect 3574 1796 3582 1798
rect 3574 1792 3576 1796
rect 3580 1792 3582 1796
rect 3574 1790 3582 1792
rect 3598 1796 3606 1798
rect 3598 1792 3600 1796
rect 3604 1792 3606 1796
rect 3598 1790 3606 1792
rect 3622 1796 3630 1798
rect 3622 1792 3624 1796
rect 3628 1792 3630 1796
rect 3622 1790 3630 1792
rect 3646 1796 3654 1798
rect 3646 1792 3648 1796
rect 3652 1792 3654 1796
rect 3646 1790 3654 1792
rect 3670 1796 3678 1798
rect 3670 1792 3672 1796
rect 3676 1792 3678 1796
rect 3670 1790 3678 1792
rect 3694 1796 3702 1798
rect 3694 1792 3696 1796
rect 3700 1792 3702 1796
rect 3694 1790 3702 1792
rect 3910 1796 3918 1798
rect 3910 1792 3912 1796
rect 3916 1792 3918 1796
rect 3910 1790 3918 1792
rect 3934 1796 3942 1798
rect 3934 1792 3936 1796
rect 3940 1792 3942 1796
rect 3934 1790 3942 1792
rect 3958 1796 3966 1798
rect 3958 1792 3960 1796
rect 3964 1792 3966 1796
rect 3958 1790 3966 1792
rect 3982 1796 3990 1798
rect 3982 1792 3984 1796
rect 3988 1792 3990 1796
rect 3982 1790 3990 1792
rect 4006 1796 4014 1798
rect 4006 1792 4008 1796
rect 4012 1792 4014 1796
rect 4006 1790 4014 1792
rect 4030 1796 4038 1798
rect 4030 1792 4032 1796
rect 4036 1792 4038 1796
rect 4030 1790 4038 1792
rect 4054 1796 4062 1798
rect 4054 1792 4056 1796
rect 4060 1792 4062 1796
rect 4054 1790 4062 1792
rect 4078 1796 4086 1798
rect 4078 1792 4080 1796
rect 4084 1792 4086 1796
rect 4078 1790 4086 1792
rect 4102 1796 4110 1798
rect 4102 1792 4104 1796
rect 4108 1792 4110 1796
rect 4102 1790 4110 1792
rect 4126 1796 4134 1798
rect 4126 1792 4128 1796
rect 4132 1792 4134 1796
rect 4126 1790 4134 1792
rect 4150 1796 4158 1798
rect 4150 1792 4152 1796
rect 4156 1792 4158 1796
rect 4150 1790 4158 1792
rect 4174 1796 4182 1798
rect 4174 1792 4176 1796
rect 4180 1792 4182 1796
rect 4174 1790 4182 1792
rect 4198 1796 4206 1798
rect 4198 1792 4200 1796
rect 4204 1792 4206 1796
rect 4198 1790 4206 1792
rect 4222 1796 4230 1798
rect 4222 1792 4224 1796
rect 4228 1792 4230 1796
rect 4222 1790 4230 1792
rect 4246 1796 4254 1798
rect 4246 1792 4248 1796
rect 4252 1792 4254 1796
rect 4246 1790 4254 1792
rect 4270 1796 4278 1798
rect 4270 1792 4272 1796
rect 4276 1792 4278 1796
rect 4270 1790 4278 1792
rect 4294 1796 4302 1798
rect 4294 1792 4296 1796
rect 4300 1792 4302 1796
rect 4294 1790 4302 1792
rect 4510 1796 4518 1798
rect 4510 1792 4512 1796
rect 4516 1792 4518 1796
rect 4510 1790 4518 1792
rect 4534 1796 4542 1798
rect 4534 1792 4536 1796
rect 4540 1792 4542 1796
rect 4534 1790 4542 1792
rect 4558 1796 4566 1798
rect 4558 1792 4560 1796
rect 4564 1792 4566 1796
rect 4558 1790 4566 1792
rect 4582 1796 4590 1798
rect 4582 1792 4584 1796
rect 4588 1792 4590 1796
rect 4582 1790 4590 1792
rect 4606 1796 4614 1798
rect 4606 1792 4608 1796
rect 4612 1792 4614 1796
rect 4606 1790 4614 1792
rect 4630 1796 4638 1798
rect 4630 1792 4632 1796
rect 4636 1792 4638 1796
rect 4630 1790 4638 1792
rect 4654 1796 4662 1798
rect 4654 1792 4656 1796
rect 4660 1792 4662 1796
rect 4654 1790 4662 1792
rect 4678 1796 4686 1798
rect 4678 1792 4680 1796
rect 4684 1792 4686 1796
rect 4678 1790 4686 1792
rect 4702 1796 4710 1798
rect 4702 1792 4704 1796
rect 4708 1792 4710 1796
rect 4702 1790 4710 1792
rect 4726 1796 4734 1798
rect 4726 1792 4728 1796
rect 4732 1792 4734 1796
rect 4726 1790 4734 1792
rect 4750 1796 4758 1798
rect 4750 1792 4752 1796
rect 4756 1792 4758 1796
rect 4750 1790 4758 1792
rect 4774 1796 4782 1798
rect 4774 1792 4776 1796
rect 4780 1792 4782 1796
rect 4774 1790 4782 1792
rect 4798 1790 4800 1798
rect 5710 1796 5718 1798
rect 5710 1792 5712 1796
rect 5716 1792 5718 1796
rect 5710 1790 5718 1792
rect 5734 1796 5742 1798
rect 5734 1792 5736 1796
rect 5740 1792 5742 1796
rect 5734 1790 5742 1792
rect 5758 1796 5766 1798
rect 5758 1792 5760 1796
rect 5764 1792 5766 1796
rect 5758 1790 5766 1792
rect 5782 1796 5790 1798
rect 5782 1792 5784 1796
rect 5788 1792 5790 1796
rect 5782 1790 5790 1792
rect 5806 1796 5814 1798
rect 5806 1792 5808 1796
rect 5812 1792 5814 1796
rect 5806 1790 5814 1792
rect 5830 1796 5838 1798
rect 5830 1792 5832 1796
rect 5836 1792 5838 1796
rect 5830 1790 5838 1792
rect 5854 1796 5862 1798
rect 5854 1792 5856 1796
rect 5860 1792 5862 1796
rect 5854 1790 5862 1792
rect 5878 1796 5886 1798
rect 5878 1792 5880 1796
rect 5884 1792 5886 1796
rect 5878 1790 5886 1792
rect 5902 1796 5910 1798
rect 5902 1792 5904 1796
rect 5908 1792 5910 1796
rect 5902 1790 5910 1792
rect 5926 1796 5934 1798
rect 5926 1792 5928 1796
rect 5932 1792 5934 1796
rect 5926 1790 5934 1792
rect 5950 1796 5958 1798
rect 5950 1792 5952 1796
rect 5956 1792 5958 1796
rect 5950 1790 5958 1792
rect 5974 1796 5982 1798
rect 5974 1792 5976 1796
rect 5980 1792 5982 1796
rect 5974 1790 5982 1792
rect 5998 1796 6006 1798
rect 5998 1792 6000 1796
rect 6004 1792 6006 1796
rect 5998 1790 6006 1792
rect 6022 1796 6030 1798
rect 6022 1792 6024 1796
rect 6028 1792 6030 1796
rect 6022 1790 6030 1792
rect 6046 1796 6054 1798
rect 6046 1792 6048 1796
rect 6052 1792 6054 1796
rect 6046 1790 6054 1792
rect 6070 1796 6078 1798
rect 6070 1792 6072 1796
rect 6076 1792 6078 1796
rect 6070 1790 6078 1792
rect 6094 1796 6102 1798
rect 6094 1792 6096 1796
rect 6100 1792 6102 1796
rect 6094 1790 6102 1792
rect 6310 1796 6318 1798
rect 6310 1792 6312 1796
rect 6316 1792 6318 1796
rect 6310 1790 6318 1792
rect 6334 1796 6342 1798
rect 6334 1792 6336 1796
rect 6340 1792 6342 1796
rect 6334 1790 6342 1792
rect 6358 1796 6366 1798
rect 6358 1792 6360 1796
rect 6364 1792 6366 1796
rect 6358 1790 6366 1792
rect 6382 1796 6390 1798
rect 6382 1792 6384 1796
rect 6388 1792 6390 1796
rect 6382 1790 6390 1792
rect 6406 1796 6414 1798
rect 6406 1792 6408 1796
rect 6412 1792 6414 1796
rect 6406 1790 6414 1792
rect 6430 1796 6438 1798
rect 6430 1792 6432 1796
rect 6436 1792 6438 1796
rect 6430 1790 6438 1792
rect 6454 1796 6462 1798
rect 6454 1792 6456 1796
rect 6460 1792 6462 1796
rect 6454 1790 6462 1792
rect 6478 1796 6486 1798
rect 6478 1792 6480 1796
rect 6484 1792 6486 1796
rect 6478 1790 6486 1792
rect 6502 1796 6510 1798
rect 6502 1792 6504 1796
rect 6508 1792 6510 1796
rect 6502 1790 6510 1792
rect 6526 1796 6534 1798
rect 6526 1792 6528 1796
rect 6532 1792 6534 1796
rect 6526 1790 6534 1792
rect 6550 1796 6558 1798
rect 6550 1792 6552 1796
rect 6556 1792 6558 1796
rect 6550 1790 6558 1792
rect 6574 1796 6582 1798
rect 6574 1792 6576 1796
rect 6580 1792 6582 1796
rect 6574 1790 6582 1792
rect 6598 1796 6606 1798
rect 6598 1792 6600 1796
rect 6604 1792 6606 1796
rect 6598 1790 6606 1792
rect 6622 1796 6630 1798
rect 6622 1792 6624 1796
rect 6628 1792 6630 1796
rect 6622 1790 6630 1792
rect 6646 1796 6654 1798
rect 6646 1792 6648 1796
rect 6652 1792 6654 1796
rect 6646 1790 6654 1792
rect 6670 1796 6678 1798
rect 6670 1792 6672 1796
rect 6676 1792 6678 1796
rect 6670 1790 6678 1792
rect 6694 1796 6702 1798
rect 6694 1792 6696 1796
rect 6700 1792 6702 1796
rect 6694 1790 6702 1792
rect 6910 1796 6918 1798
rect 6910 1792 6912 1796
rect 6916 1792 6918 1796
rect 6910 1790 6918 1792
rect 6934 1796 6942 1798
rect 6934 1792 6936 1796
rect 6940 1792 6942 1796
rect 6934 1790 6942 1792
rect 6958 1796 6966 1798
rect 6958 1792 6960 1796
rect 6964 1792 6966 1796
rect 6958 1790 6966 1792
rect 6982 1796 6990 1798
rect 6982 1792 6984 1796
rect 6988 1792 6990 1796
rect 6982 1790 6990 1792
rect 7006 1796 7014 1798
rect 7006 1792 7008 1796
rect 7012 1792 7014 1796
rect 7006 1790 7014 1792
rect 7030 1796 7038 1798
rect 7030 1792 7032 1796
rect 7036 1792 7038 1796
rect 7030 1790 7038 1792
rect 7054 1796 7062 1798
rect 7054 1792 7056 1796
rect 7060 1792 7062 1796
rect 7054 1790 7062 1792
rect 7078 1796 7086 1798
rect 7078 1792 7080 1796
rect 7084 1792 7086 1796
rect 7078 1790 7086 1792
rect 7102 1796 7110 1798
rect 7102 1792 7104 1796
rect 7108 1792 7110 1796
rect 7102 1790 7110 1792
rect 7126 1796 7134 1798
rect 7126 1792 7128 1796
rect 7132 1792 7134 1796
rect 7126 1790 7134 1792
rect 7150 1796 7158 1798
rect 7150 1792 7152 1796
rect 7156 1792 7158 1796
rect 7150 1790 7158 1792
rect 7174 1796 7182 1798
rect 7174 1792 7176 1796
rect 7180 1792 7182 1796
rect 7174 1790 7182 1792
rect 7198 1790 7200 1798
rect 2410 1784 2418 1786
rect 2410 1780 2412 1784
rect 2416 1780 2418 1784
rect 2410 1778 2418 1780
rect 2434 1784 2442 1786
rect 2434 1780 2436 1784
rect 2440 1780 2442 1784
rect 2434 1778 2442 1780
rect 2458 1784 2466 1786
rect 2458 1780 2460 1784
rect 2464 1780 2466 1784
rect 2458 1778 2466 1780
rect 2482 1784 2490 1786
rect 2482 1780 2484 1784
rect 2488 1780 2490 1784
rect 2482 1778 2490 1780
rect 2698 1784 2706 1786
rect 2698 1780 2700 1784
rect 2704 1780 2706 1784
rect 2698 1778 2706 1780
rect 2722 1784 2730 1786
rect 2722 1780 2724 1784
rect 2728 1780 2730 1784
rect 2722 1778 2730 1780
rect 2746 1784 2754 1786
rect 2746 1780 2748 1784
rect 2752 1780 2754 1784
rect 2746 1778 2754 1780
rect 2770 1784 2778 1786
rect 2770 1780 2772 1784
rect 2776 1780 2778 1784
rect 2770 1778 2778 1780
rect 2794 1784 2802 1786
rect 2794 1780 2796 1784
rect 2800 1780 2802 1784
rect 2794 1778 2802 1780
rect 2818 1784 2826 1786
rect 2818 1780 2820 1784
rect 2824 1780 2826 1784
rect 2818 1778 2826 1780
rect 2842 1784 2850 1786
rect 2842 1780 2844 1784
rect 2848 1780 2850 1784
rect 2842 1778 2850 1780
rect 2866 1784 2874 1786
rect 2866 1780 2868 1784
rect 2872 1780 2874 1784
rect 2866 1778 2874 1780
rect 2890 1784 2898 1786
rect 2890 1780 2892 1784
rect 2896 1780 2898 1784
rect 2890 1778 2898 1780
rect 2914 1784 2922 1786
rect 2914 1780 2916 1784
rect 2920 1780 2922 1784
rect 2914 1778 2922 1780
rect 2938 1784 2946 1786
rect 2938 1780 2940 1784
rect 2944 1780 2946 1784
rect 2938 1778 2946 1780
rect 2962 1784 2970 1786
rect 2962 1780 2964 1784
rect 2968 1780 2970 1784
rect 2962 1778 2970 1780
rect 2986 1784 2994 1786
rect 2986 1780 2988 1784
rect 2992 1780 2994 1784
rect 2986 1778 2994 1780
rect 3010 1784 3018 1786
rect 3010 1780 3012 1784
rect 3016 1780 3018 1784
rect 3010 1778 3018 1780
rect 3034 1784 3042 1786
rect 3034 1780 3036 1784
rect 3040 1780 3042 1784
rect 3034 1778 3042 1780
rect 3058 1784 3066 1786
rect 3058 1780 3060 1784
rect 3064 1780 3066 1784
rect 3058 1778 3066 1780
rect 3082 1784 3090 1786
rect 3082 1780 3084 1784
rect 3088 1780 3090 1784
rect 3082 1778 3090 1780
rect 3298 1784 3306 1786
rect 3298 1780 3300 1784
rect 3304 1780 3306 1784
rect 3298 1778 3306 1780
rect 3322 1784 3330 1786
rect 3322 1780 3324 1784
rect 3328 1780 3330 1784
rect 3322 1778 3330 1780
rect 3346 1784 3354 1786
rect 3346 1780 3348 1784
rect 3352 1780 3354 1784
rect 3346 1778 3354 1780
rect 3370 1784 3378 1786
rect 3370 1780 3372 1784
rect 3376 1780 3378 1784
rect 3370 1778 3378 1780
rect 3394 1784 3402 1786
rect 3394 1780 3396 1784
rect 3400 1780 3402 1784
rect 3394 1778 3402 1780
rect 3418 1784 3426 1786
rect 3418 1780 3420 1784
rect 3424 1780 3426 1784
rect 3418 1778 3426 1780
rect 3442 1784 3450 1786
rect 3442 1780 3444 1784
rect 3448 1780 3450 1784
rect 3442 1778 3450 1780
rect 3466 1784 3474 1786
rect 3466 1780 3468 1784
rect 3472 1780 3474 1784
rect 3466 1778 3474 1780
rect 3490 1784 3498 1786
rect 3490 1780 3492 1784
rect 3496 1780 3498 1784
rect 3490 1778 3498 1780
rect 3514 1784 3522 1786
rect 3514 1780 3516 1784
rect 3520 1780 3522 1784
rect 3514 1778 3522 1780
rect 3538 1784 3546 1786
rect 3538 1780 3540 1784
rect 3544 1780 3546 1784
rect 3538 1778 3546 1780
rect 3562 1784 3570 1786
rect 3562 1780 3564 1784
rect 3568 1780 3570 1784
rect 3562 1778 3570 1780
rect 3586 1784 3594 1786
rect 3586 1780 3588 1784
rect 3592 1780 3594 1784
rect 3586 1778 3594 1780
rect 3610 1784 3618 1786
rect 3610 1780 3612 1784
rect 3616 1780 3618 1784
rect 3610 1778 3618 1780
rect 3634 1784 3642 1786
rect 3634 1780 3636 1784
rect 3640 1780 3642 1784
rect 3634 1778 3642 1780
rect 3658 1784 3666 1786
rect 3658 1780 3660 1784
rect 3664 1780 3666 1784
rect 3658 1778 3666 1780
rect 3682 1784 3690 1786
rect 3682 1780 3684 1784
rect 3688 1780 3690 1784
rect 3682 1778 3690 1780
rect 3898 1784 3906 1786
rect 3898 1780 3900 1784
rect 3904 1780 3906 1784
rect 3898 1778 3906 1780
rect 3922 1784 3930 1786
rect 3922 1780 3924 1784
rect 3928 1780 3930 1784
rect 3922 1778 3930 1780
rect 3946 1784 3954 1786
rect 3946 1780 3948 1784
rect 3952 1780 3954 1784
rect 3946 1778 3954 1780
rect 3970 1784 3978 1786
rect 3970 1780 3972 1784
rect 3976 1780 3978 1784
rect 3970 1778 3978 1780
rect 3994 1784 4002 1786
rect 3994 1780 3996 1784
rect 4000 1780 4002 1784
rect 3994 1778 4002 1780
rect 4018 1784 4026 1786
rect 4018 1780 4020 1784
rect 4024 1780 4026 1784
rect 4018 1778 4026 1780
rect 4042 1784 4050 1786
rect 4042 1780 4044 1784
rect 4048 1780 4050 1784
rect 4042 1778 4050 1780
rect 4066 1784 4074 1786
rect 4066 1780 4068 1784
rect 4072 1780 4074 1784
rect 4066 1778 4074 1780
rect 4090 1784 4098 1786
rect 4090 1780 4092 1784
rect 4096 1780 4098 1784
rect 4090 1778 4098 1780
rect 4114 1784 4122 1786
rect 4114 1780 4116 1784
rect 4120 1780 4122 1784
rect 4114 1778 4122 1780
rect 4138 1784 4146 1786
rect 4138 1780 4140 1784
rect 4144 1780 4146 1784
rect 4138 1778 4146 1780
rect 4162 1784 4170 1786
rect 4162 1780 4164 1784
rect 4168 1780 4170 1784
rect 4162 1778 4170 1780
rect 4186 1784 4194 1786
rect 4186 1780 4188 1784
rect 4192 1780 4194 1784
rect 4186 1778 4194 1780
rect 4210 1784 4218 1786
rect 4210 1780 4212 1784
rect 4216 1780 4218 1784
rect 4210 1778 4218 1780
rect 4234 1784 4242 1786
rect 4234 1780 4236 1784
rect 4240 1780 4242 1784
rect 4234 1778 4242 1780
rect 4258 1784 4266 1786
rect 4258 1780 4260 1784
rect 4264 1780 4266 1784
rect 4258 1778 4266 1780
rect 4282 1784 4290 1786
rect 4282 1780 4284 1784
rect 4288 1780 4290 1784
rect 4282 1778 4290 1780
rect 4498 1784 4506 1786
rect 4498 1780 4500 1784
rect 4504 1780 4506 1784
rect 4498 1778 4506 1780
rect 4522 1784 4530 1786
rect 4522 1780 4524 1784
rect 4528 1780 4530 1784
rect 4522 1778 4530 1780
rect 4546 1784 4554 1786
rect 4546 1780 4548 1784
rect 4552 1780 4554 1784
rect 4546 1778 4554 1780
rect 4570 1784 4578 1786
rect 4570 1780 4572 1784
rect 4576 1780 4578 1784
rect 4570 1778 4578 1780
rect 4594 1784 4602 1786
rect 4594 1780 4596 1784
rect 4600 1780 4602 1784
rect 4594 1778 4602 1780
rect 4618 1784 4626 1786
rect 4618 1780 4620 1784
rect 4624 1780 4626 1784
rect 4618 1778 4626 1780
rect 4642 1784 4650 1786
rect 4642 1780 4644 1784
rect 4648 1780 4650 1784
rect 4642 1778 4650 1780
rect 4666 1784 4674 1786
rect 4666 1780 4668 1784
rect 4672 1780 4674 1784
rect 4666 1778 4674 1780
rect 4690 1784 4698 1786
rect 4690 1780 4692 1784
rect 4696 1780 4698 1784
rect 4690 1778 4698 1780
rect 4714 1784 4722 1786
rect 4714 1780 4716 1784
rect 4720 1780 4722 1784
rect 4714 1778 4722 1780
rect 4738 1784 4746 1786
rect 4738 1780 4740 1784
rect 4744 1780 4746 1784
rect 4738 1778 4746 1780
rect 4762 1784 4770 1786
rect 4762 1780 4764 1784
rect 4768 1780 4770 1784
rect 4762 1778 4770 1780
rect 4786 1784 4794 1786
rect 4786 1780 4788 1784
rect 4792 1780 4794 1784
rect 4786 1778 4794 1780
rect 5698 1784 5706 1786
rect 5698 1780 5700 1784
rect 5704 1780 5706 1784
rect 5698 1778 5706 1780
rect 5722 1784 5730 1786
rect 5722 1780 5724 1784
rect 5728 1780 5730 1784
rect 5722 1778 5730 1780
rect 5746 1784 5754 1786
rect 5746 1780 5748 1784
rect 5752 1780 5754 1784
rect 5746 1778 5754 1780
rect 5770 1784 5778 1786
rect 5770 1780 5772 1784
rect 5776 1780 5778 1784
rect 5770 1778 5778 1780
rect 5794 1784 5802 1786
rect 5794 1780 5796 1784
rect 5800 1780 5802 1784
rect 5794 1778 5802 1780
rect 5818 1784 5826 1786
rect 5818 1780 5820 1784
rect 5824 1780 5826 1784
rect 5818 1778 5826 1780
rect 5842 1784 5850 1786
rect 5842 1780 5844 1784
rect 5848 1780 5850 1784
rect 5842 1778 5850 1780
rect 5866 1784 5874 1786
rect 5866 1780 5868 1784
rect 5872 1780 5874 1784
rect 5866 1778 5874 1780
rect 5890 1784 5898 1786
rect 5890 1780 5892 1784
rect 5896 1780 5898 1784
rect 5890 1778 5898 1780
rect 5914 1784 5922 1786
rect 5914 1780 5916 1784
rect 5920 1780 5922 1784
rect 5914 1778 5922 1780
rect 5938 1784 5946 1786
rect 5938 1780 5940 1784
rect 5944 1780 5946 1784
rect 5938 1778 5946 1780
rect 5962 1784 5970 1786
rect 5962 1780 5964 1784
rect 5968 1780 5970 1784
rect 5962 1778 5970 1780
rect 5986 1784 5994 1786
rect 5986 1780 5988 1784
rect 5992 1780 5994 1784
rect 5986 1778 5994 1780
rect 6010 1784 6018 1786
rect 6010 1780 6012 1784
rect 6016 1780 6018 1784
rect 6010 1778 6018 1780
rect 6034 1784 6042 1786
rect 6034 1780 6036 1784
rect 6040 1780 6042 1784
rect 6034 1778 6042 1780
rect 6058 1784 6066 1786
rect 6058 1780 6060 1784
rect 6064 1780 6066 1784
rect 6058 1778 6066 1780
rect 6082 1784 6090 1786
rect 6082 1780 6084 1784
rect 6088 1780 6090 1784
rect 6082 1778 6090 1780
rect 6298 1784 6306 1786
rect 6298 1780 6300 1784
rect 6304 1780 6306 1784
rect 6298 1778 6306 1780
rect 6322 1784 6330 1786
rect 6322 1780 6324 1784
rect 6328 1780 6330 1784
rect 6322 1778 6330 1780
rect 6346 1784 6354 1786
rect 6346 1780 6348 1784
rect 6352 1780 6354 1784
rect 6346 1778 6354 1780
rect 6370 1784 6378 1786
rect 6370 1780 6372 1784
rect 6376 1780 6378 1784
rect 6370 1778 6378 1780
rect 6394 1784 6402 1786
rect 6394 1780 6396 1784
rect 6400 1780 6402 1784
rect 6394 1778 6402 1780
rect 6418 1784 6426 1786
rect 6418 1780 6420 1784
rect 6424 1780 6426 1784
rect 6418 1778 6426 1780
rect 6442 1784 6450 1786
rect 6442 1780 6444 1784
rect 6448 1780 6450 1784
rect 6442 1778 6450 1780
rect 6466 1784 6474 1786
rect 6466 1780 6468 1784
rect 6472 1780 6474 1784
rect 6466 1778 6474 1780
rect 6490 1784 6498 1786
rect 6490 1780 6492 1784
rect 6496 1780 6498 1784
rect 6490 1778 6498 1780
rect 6514 1784 6522 1786
rect 6514 1780 6516 1784
rect 6520 1780 6522 1784
rect 6514 1778 6522 1780
rect 6538 1784 6546 1786
rect 6538 1780 6540 1784
rect 6544 1780 6546 1784
rect 6538 1778 6546 1780
rect 6562 1784 6570 1786
rect 6562 1780 6564 1784
rect 6568 1780 6570 1784
rect 6562 1778 6570 1780
rect 6586 1784 6594 1786
rect 6586 1780 6588 1784
rect 6592 1780 6594 1784
rect 6586 1778 6594 1780
rect 6610 1784 6618 1786
rect 6610 1780 6612 1784
rect 6616 1780 6618 1784
rect 6610 1778 6618 1780
rect 6634 1784 6642 1786
rect 6634 1780 6636 1784
rect 6640 1780 6642 1784
rect 6634 1778 6642 1780
rect 6658 1784 6666 1786
rect 6658 1780 6660 1784
rect 6664 1780 6666 1784
rect 6658 1778 6666 1780
rect 6682 1784 6690 1786
rect 6682 1780 6684 1784
rect 6688 1780 6690 1784
rect 6682 1778 6690 1780
rect 6898 1784 6906 1786
rect 6898 1780 6900 1784
rect 6904 1780 6906 1784
rect 6898 1778 6906 1780
rect 6922 1784 6930 1786
rect 6922 1780 6924 1784
rect 6928 1780 6930 1784
rect 6922 1778 6930 1780
rect 6946 1784 6954 1786
rect 6946 1780 6948 1784
rect 6952 1780 6954 1784
rect 6946 1778 6954 1780
rect 6970 1784 6978 1786
rect 6970 1780 6972 1784
rect 6976 1780 6978 1784
rect 6970 1778 6978 1780
rect 6994 1784 7002 1786
rect 6994 1780 6996 1784
rect 7000 1780 7002 1784
rect 6994 1778 7002 1780
rect 7018 1784 7026 1786
rect 7018 1780 7020 1784
rect 7024 1780 7026 1784
rect 7018 1778 7026 1780
rect 7042 1784 7050 1786
rect 7042 1780 7044 1784
rect 7048 1780 7050 1784
rect 7042 1778 7050 1780
rect 7066 1784 7074 1786
rect 7066 1780 7068 1784
rect 7072 1780 7074 1784
rect 7066 1778 7074 1780
rect 7090 1784 7098 1786
rect 7090 1780 7092 1784
rect 7096 1780 7098 1784
rect 7090 1778 7098 1780
rect 7114 1784 7122 1786
rect 7114 1780 7116 1784
rect 7120 1780 7122 1784
rect 7114 1778 7122 1780
rect 7138 1784 7146 1786
rect 7138 1780 7140 1784
rect 7144 1780 7146 1784
rect 7138 1778 7146 1780
rect 7162 1784 7170 1786
rect 7162 1780 7164 1784
rect 7168 1780 7170 1784
rect 7162 1778 7170 1780
rect 7186 1784 7194 1786
rect 7186 1780 7188 1784
rect 7192 1780 7194 1784
rect 7186 1778 7194 1780
rect 2400 1772 2406 1774
rect 2404 1768 2406 1772
rect 2400 1766 2406 1768
rect 2422 1772 2430 1774
rect 2422 1768 2424 1772
rect 2428 1768 2430 1772
rect 2422 1766 2430 1768
rect 2446 1772 2454 1774
rect 2446 1768 2448 1772
rect 2452 1768 2454 1772
rect 2446 1766 2454 1768
rect 2470 1772 2478 1774
rect 2470 1768 2472 1772
rect 2476 1768 2478 1772
rect 2470 1766 2478 1768
rect 2494 1772 2502 1774
rect 2494 1768 2496 1772
rect 2500 1768 2502 1772
rect 2494 1766 2502 1768
rect 2710 1772 2718 1774
rect 2710 1768 2712 1772
rect 2716 1768 2718 1772
rect 2710 1766 2718 1768
rect 2734 1772 2742 1774
rect 2734 1768 2736 1772
rect 2740 1768 2742 1772
rect 2734 1766 2742 1768
rect 2758 1772 2766 1774
rect 2758 1768 2760 1772
rect 2764 1768 2766 1772
rect 2758 1766 2766 1768
rect 2782 1772 2790 1774
rect 2782 1768 2784 1772
rect 2788 1768 2790 1772
rect 2782 1766 2790 1768
rect 2806 1772 2814 1774
rect 2806 1768 2808 1772
rect 2812 1768 2814 1772
rect 2806 1766 2814 1768
rect 2830 1772 2838 1774
rect 2830 1768 2832 1772
rect 2836 1768 2838 1772
rect 2830 1766 2838 1768
rect 2854 1772 2862 1774
rect 2854 1768 2856 1772
rect 2860 1768 2862 1772
rect 2854 1766 2862 1768
rect 2878 1772 2886 1774
rect 2878 1768 2880 1772
rect 2884 1768 2886 1772
rect 2878 1766 2886 1768
rect 2902 1772 2910 1774
rect 2902 1768 2904 1772
rect 2908 1768 2910 1772
rect 2902 1766 2910 1768
rect 2926 1772 2934 1774
rect 2926 1768 2928 1772
rect 2932 1768 2934 1772
rect 2926 1766 2934 1768
rect 2950 1772 2958 1774
rect 2950 1768 2952 1772
rect 2956 1768 2958 1772
rect 2950 1766 2958 1768
rect 2974 1772 2982 1774
rect 2974 1768 2976 1772
rect 2980 1768 2982 1772
rect 2974 1766 2982 1768
rect 2998 1772 3006 1774
rect 2998 1768 3000 1772
rect 3004 1768 3006 1772
rect 2998 1766 3006 1768
rect 3022 1772 3030 1774
rect 3022 1768 3024 1772
rect 3028 1768 3030 1772
rect 3022 1766 3030 1768
rect 3046 1772 3054 1774
rect 3046 1768 3048 1772
rect 3052 1768 3054 1772
rect 3046 1766 3054 1768
rect 3070 1772 3078 1774
rect 3070 1768 3072 1772
rect 3076 1768 3078 1772
rect 3070 1766 3078 1768
rect 3094 1772 3102 1774
rect 3094 1768 3096 1772
rect 3100 1768 3102 1772
rect 3094 1766 3102 1768
rect 3310 1772 3318 1774
rect 3310 1768 3312 1772
rect 3316 1768 3318 1772
rect 3310 1766 3318 1768
rect 3334 1772 3342 1774
rect 3334 1768 3336 1772
rect 3340 1768 3342 1772
rect 3334 1766 3342 1768
rect 3358 1772 3366 1774
rect 3358 1768 3360 1772
rect 3364 1768 3366 1772
rect 3358 1766 3366 1768
rect 3382 1772 3390 1774
rect 3382 1768 3384 1772
rect 3388 1768 3390 1772
rect 3382 1766 3390 1768
rect 3406 1772 3414 1774
rect 3406 1768 3408 1772
rect 3412 1768 3414 1772
rect 3406 1766 3414 1768
rect 3430 1772 3438 1774
rect 3430 1768 3432 1772
rect 3436 1768 3438 1772
rect 3430 1766 3438 1768
rect 3454 1772 3462 1774
rect 3454 1768 3456 1772
rect 3460 1768 3462 1772
rect 3454 1766 3462 1768
rect 3478 1772 3486 1774
rect 3478 1768 3480 1772
rect 3484 1768 3486 1772
rect 3478 1766 3486 1768
rect 3502 1772 3510 1774
rect 3502 1768 3504 1772
rect 3508 1768 3510 1772
rect 3502 1766 3510 1768
rect 3526 1772 3534 1774
rect 3526 1768 3528 1772
rect 3532 1768 3534 1772
rect 3526 1766 3534 1768
rect 3550 1772 3558 1774
rect 3550 1768 3552 1772
rect 3556 1768 3558 1772
rect 3550 1766 3558 1768
rect 3574 1772 3582 1774
rect 3574 1768 3576 1772
rect 3580 1768 3582 1772
rect 3574 1766 3582 1768
rect 3598 1772 3606 1774
rect 3598 1768 3600 1772
rect 3604 1768 3606 1772
rect 3598 1766 3606 1768
rect 3622 1772 3630 1774
rect 3622 1768 3624 1772
rect 3628 1768 3630 1772
rect 3622 1766 3630 1768
rect 3646 1772 3654 1774
rect 3646 1768 3648 1772
rect 3652 1768 3654 1772
rect 3646 1766 3654 1768
rect 3670 1772 3678 1774
rect 3670 1768 3672 1772
rect 3676 1768 3678 1772
rect 3670 1766 3678 1768
rect 3694 1772 3702 1774
rect 3694 1768 3696 1772
rect 3700 1768 3702 1772
rect 3694 1766 3702 1768
rect 3910 1772 3918 1774
rect 3910 1768 3912 1772
rect 3916 1768 3918 1772
rect 3910 1766 3918 1768
rect 3934 1772 3942 1774
rect 3934 1768 3936 1772
rect 3940 1768 3942 1772
rect 3934 1766 3942 1768
rect 3958 1772 3966 1774
rect 3958 1768 3960 1772
rect 3964 1768 3966 1772
rect 3958 1766 3966 1768
rect 3982 1772 3990 1774
rect 3982 1768 3984 1772
rect 3988 1768 3990 1772
rect 3982 1766 3990 1768
rect 4006 1772 4014 1774
rect 4006 1768 4008 1772
rect 4012 1768 4014 1772
rect 4006 1766 4014 1768
rect 4030 1772 4038 1774
rect 4030 1768 4032 1772
rect 4036 1768 4038 1772
rect 4030 1766 4038 1768
rect 4054 1772 4062 1774
rect 4054 1768 4056 1772
rect 4060 1768 4062 1772
rect 4054 1766 4062 1768
rect 4078 1772 4086 1774
rect 4078 1768 4080 1772
rect 4084 1768 4086 1772
rect 4078 1766 4086 1768
rect 4102 1772 4110 1774
rect 4102 1768 4104 1772
rect 4108 1768 4110 1772
rect 4102 1766 4110 1768
rect 4126 1772 4134 1774
rect 4126 1768 4128 1772
rect 4132 1768 4134 1772
rect 4126 1766 4134 1768
rect 4150 1772 4158 1774
rect 4150 1768 4152 1772
rect 4156 1768 4158 1772
rect 4150 1766 4158 1768
rect 4174 1772 4182 1774
rect 4174 1768 4176 1772
rect 4180 1768 4182 1772
rect 4174 1766 4182 1768
rect 4198 1772 4206 1774
rect 4198 1768 4200 1772
rect 4204 1768 4206 1772
rect 4198 1766 4206 1768
rect 4222 1772 4230 1774
rect 4222 1768 4224 1772
rect 4228 1768 4230 1772
rect 4222 1766 4230 1768
rect 4246 1772 4254 1774
rect 4246 1768 4248 1772
rect 4252 1768 4254 1772
rect 4246 1766 4254 1768
rect 4270 1772 4278 1774
rect 4270 1768 4272 1772
rect 4276 1768 4278 1772
rect 4270 1766 4278 1768
rect 4294 1772 4302 1774
rect 4294 1768 4296 1772
rect 4300 1768 4302 1772
rect 4294 1766 4302 1768
rect 4510 1772 4518 1774
rect 4510 1768 4512 1772
rect 4516 1768 4518 1772
rect 4510 1766 4518 1768
rect 4534 1772 4542 1774
rect 4534 1768 4536 1772
rect 4540 1768 4542 1772
rect 4534 1766 4542 1768
rect 4558 1772 4566 1774
rect 4558 1768 4560 1772
rect 4564 1768 4566 1772
rect 4558 1766 4566 1768
rect 4582 1772 4590 1774
rect 4582 1768 4584 1772
rect 4588 1768 4590 1772
rect 4582 1766 4590 1768
rect 4606 1772 4614 1774
rect 4606 1768 4608 1772
rect 4612 1768 4614 1772
rect 4606 1766 4614 1768
rect 4630 1772 4638 1774
rect 4630 1768 4632 1772
rect 4636 1768 4638 1772
rect 4630 1766 4638 1768
rect 4654 1772 4662 1774
rect 4654 1768 4656 1772
rect 4660 1768 4662 1772
rect 4654 1766 4662 1768
rect 4678 1772 4686 1774
rect 4678 1768 4680 1772
rect 4684 1768 4686 1772
rect 4678 1766 4686 1768
rect 4702 1772 4710 1774
rect 4702 1768 4704 1772
rect 4708 1768 4710 1772
rect 4702 1766 4710 1768
rect 4726 1772 4734 1774
rect 4726 1768 4728 1772
rect 4732 1768 4734 1772
rect 4726 1766 4734 1768
rect 4750 1772 4758 1774
rect 4750 1768 4752 1772
rect 4756 1768 4758 1772
rect 4750 1766 4758 1768
rect 4774 1772 4782 1774
rect 4774 1768 4776 1772
rect 4780 1768 4782 1772
rect 4774 1766 4782 1768
rect 4798 1766 4800 1774
rect 5710 1772 5718 1774
rect 5710 1768 5712 1772
rect 5716 1768 5718 1772
rect 5710 1766 5718 1768
rect 5734 1772 5742 1774
rect 5734 1768 5736 1772
rect 5740 1768 5742 1772
rect 5734 1766 5742 1768
rect 5758 1772 5766 1774
rect 5758 1768 5760 1772
rect 5764 1768 5766 1772
rect 5758 1766 5766 1768
rect 5782 1772 5790 1774
rect 5782 1768 5784 1772
rect 5788 1768 5790 1772
rect 5782 1766 5790 1768
rect 5806 1772 5814 1774
rect 5806 1768 5808 1772
rect 5812 1768 5814 1772
rect 5806 1766 5814 1768
rect 5830 1772 5838 1774
rect 5830 1768 5832 1772
rect 5836 1768 5838 1772
rect 5830 1766 5838 1768
rect 5854 1772 5862 1774
rect 5854 1768 5856 1772
rect 5860 1768 5862 1772
rect 5854 1766 5862 1768
rect 5878 1772 5886 1774
rect 5878 1768 5880 1772
rect 5884 1768 5886 1772
rect 5878 1766 5886 1768
rect 5902 1772 5910 1774
rect 5902 1768 5904 1772
rect 5908 1768 5910 1772
rect 5902 1766 5910 1768
rect 5926 1772 5934 1774
rect 5926 1768 5928 1772
rect 5932 1768 5934 1772
rect 5926 1766 5934 1768
rect 5950 1772 5958 1774
rect 5950 1768 5952 1772
rect 5956 1768 5958 1772
rect 5950 1766 5958 1768
rect 5974 1772 5982 1774
rect 5974 1768 5976 1772
rect 5980 1768 5982 1772
rect 5974 1766 5982 1768
rect 5998 1772 6006 1774
rect 5998 1768 6000 1772
rect 6004 1768 6006 1772
rect 5998 1766 6006 1768
rect 6022 1772 6030 1774
rect 6022 1768 6024 1772
rect 6028 1768 6030 1772
rect 6022 1766 6030 1768
rect 6046 1772 6054 1774
rect 6046 1768 6048 1772
rect 6052 1768 6054 1772
rect 6046 1766 6054 1768
rect 6070 1772 6078 1774
rect 6070 1768 6072 1772
rect 6076 1768 6078 1772
rect 6070 1766 6078 1768
rect 6094 1772 6102 1774
rect 6094 1768 6096 1772
rect 6100 1768 6102 1772
rect 6094 1766 6102 1768
rect 6310 1772 6318 1774
rect 6310 1768 6312 1772
rect 6316 1768 6318 1772
rect 6310 1766 6318 1768
rect 6334 1772 6342 1774
rect 6334 1768 6336 1772
rect 6340 1768 6342 1772
rect 6334 1766 6342 1768
rect 6358 1772 6366 1774
rect 6358 1768 6360 1772
rect 6364 1768 6366 1772
rect 6358 1766 6366 1768
rect 6382 1772 6390 1774
rect 6382 1768 6384 1772
rect 6388 1768 6390 1772
rect 6382 1766 6390 1768
rect 6406 1772 6414 1774
rect 6406 1768 6408 1772
rect 6412 1768 6414 1772
rect 6406 1766 6414 1768
rect 6430 1772 6438 1774
rect 6430 1768 6432 1772
rect 6436 1768 6438 1772
rect 6430 1766 6438 1768
rect 6454 1772 6462 1774
rect 6454 1768 6456 1772
rect 6460 1768 6462 1772
rect 6454 1766 6462 1768
rect 6478 1772 6486 1774
rect 6478 1768 6480 1772
rect 6484 1768 6486 1772
rect 6478 1766 6486 1768
rect 6502 1772 6510 1774
rect 6502 1768 6504 1772
rect 6508 1768 6510 1772
rect 6502 1766 6510 1768
rect 6526 1772 6534 1774
rect 6526 1768 6528 1772
rect 6532 1768 6534 1772
rect 6526 1766 6534 1768
rect 6550 1772 6558 1774
rect 6550 1768 6552 1772
rect 6556 1768 6558 1772
rect 6550 1766 6558 1768
rect 6574 1772 6582 1774
rect 6574 1768 6576 1772
rect 6580 1768 6582 1772
rect 6574 1766 6582 1768
rect 6598 1772 6606 1774
rect 6598 1768 6600 1772
rect 6604 1768 6606 1772
rect 6598 1766 6606 1768
rect 6622 1772 6630 1774
rect 6622 1768 6624 1772
rect 6628 1768 6630 1772
rect 6622 1766 6630 1768
rect 6646 1772 6654 1774
rect 6646 1768 6648 1772
rect 6652 1768 6654 1772
rect 6646 1766 6654 1768
rect 6670 1772 6678 1774
rect 6670 1768 6672 1772
rect 6676 1768 6678 1772
rect 6670 1766 6678 1768
rect 6694 1772 6702 1774
rect 6694 1768 6696 1772
rect 6700 1768 6702 1772
rect 6694 1766 6702 1768
rect 6910 1772 6918 1774
rect 6910 1768 6912 1772
rect 6916 1768 6918 1772
rect 6910 1766 6918 1768
rect 6934 1772 6942 1774
rect 6934 1768 6936 1772
rect 6940 1768 6942 1772
rect 6934 1766 6942 1768
rect 6958 1772 6966 1774
rect 6958 1768 6960 1772
rect 6964 1768 6966 1772
rect 6958 1766 6966 1768
rect 6982 1772 6990 1774
rect 6982 1768 6984 1772
rect 6988 1768 6990 1772
rect 6982 1766 6990 1768
rect 7006 1772 7014 1774
rect 7006 1768 7008 1772
rect 7012 1768 7014 1772
rect 7006 1766 7014 1768
rect 7030 1772 7038 1774
rect 7030 1768 7032 1772
rect 7036 1768 7038 1772
rect 7030 1766 7038 1768
rect 7054 1772 7062 1774
rect 7054 1768 7056 1772
rect 7060 1768 7062 1772
rect 7054 1766 7062 1768
rect 7078 1772 7086 1774
rect 7078 1768 7080 1772
rect 7084 1768 7086 1772
rect 7078 1766 7086 1768
rect 7102 1772 7110 1774
rect 7102 1768 7104 1772
rect 7108 1768 7110 1772
rect 7102 1766 7110 1768
rect 7126 1772 7134 1774
rect 7126 1768 7128 1772
rect 7132 1768 7134 1772
rect 7126 1766 7134 1768
rect 7150 1772 7158 1774
rect 7150 1768 7152 1772
rect 7156 1768 7158 1772
rect 7150 1766 7158 1768
rect 7174 1772 7182 1774
rect 7174 1768 7176 1772
rect 7180 1768 7182 1772
rect 7174 1766 7182 1768
rect 7198 1766 7200 1774
rect 2410 1760 2418 1762
rect 2410 1756 2412 1760
rect 2416 1756 2418 1760
rect 2410 1754 2418 1756
rect 2434 1760 2442 1762
rect 2434 1756 2436 1760
rect 2440 1756 2442 1760
rect 2434 1754 2442 1756
rect 2458 1760 2466 1762
rect 2458 1756 2460 1760
rect 2464 1756 2466 1760
rect 2458 1754 2466 1756
rect 2482 1760 2490 1762
rect 2482 1756 2484 1760
rect 2488 1756 2490 1760
rect 2482 1754 2490 1756
rect 2698 1760 2706 1762
rect 2698 1756 2700 1760
rect 2704 1756 2706 1760
rect 2698 1754 2706 1756
rect 2722 1760 2730 1762
rect 2722 1756 2724 1760
rect 2728 1756 2730 1760
rect 2722 1754 2730 1756
rect 2746 1760 2754 1762
rect 2746 1756 2748 1760
rect 2752 1756 2754 1760
rect 2746 1754 2754 1756
rect 2770 1760 2778 1762
rect 2770 1756 2772 1760
rect 2776 1756 2778 1760
rect 2770 1754 2778 1756
rect 2794 1760 2802 1762
rect 2794 1756 2796 1760
rect 2800 1756 2802 1760
rect 2794 1754 2802 1756
rect 2818 1760 2826 1762
rect 2818 1756 2820 1760
rect 2824 1756 2826 1760
rect 2818 1754 2826 1756
rect 2842 1760 2850 1762
rect 2842 1756 2844 1760
rect 2848 1756 2850 1760
rect 2842 1754 2850 1756
rect 2866 1760 2874 1762
rect 2866 1756 2868 1760
rect 2872 1756 2874 1760
rect 2866 1754 2874 1756
rect 2890 1760 2898 1762
rect 2890 1756 2892 1760
rect 2896 1756 2898 1760
rect 2890 1754 2898 1756
rect 2914 1760 2922 1762
rect 2914 1756 2916 1760
rect 2920 1756 2922 1760
rect 2914 1754 2922 1756
rect 2938 1760 2946 1762
rect 2938 1756 2940 1760
rect 2944 1756 2946 1760
rect 2938 1754 2946 1756
rect 2962 1760 2970 1762
rect 2962 1756 2964 1760
rect 2968 1756 2970 1760
rect 2962 1754 2970 1756
rect 2986 1760 2994 1762
rect 2986 1756 2988 1760
rect 2992 1756 2994 1760
rect 2986 1754 2994 1756
rect 3010 1760 3018 1762
rect 3010 1756 3012 1760
rect 3016 1756 3018 1760
rect 3010 1754 3018 1756
rect 3034 1760 3042 1762
rect 3034 1756 3036 1760
rect 3040 1756 3042 1760
rect 3034 1754 3042 1756
rect 3058 1760 3066 1762
rect 3058 1756 3060 1760
rect 3064 1756 3066 1760
rect 3058 1754 3066 1756
rect 3082 1760 3090 1762
rect 3082 1756 3084 1760
rect 3088 1756 3090 1760
rect 3082 1754 3090 1756
rect 3298 1760 3306 1762
rect 3298 1756 3300 1760
rect 3304 1756 3306 1760
rect 3298 1754 3306 1756
rect 3322 1760 3330 1762
rect 3322 1756 3324 1760
rect 3328 1756 3330 1760
rect 3322 1754 3330 1756
rect 3346 1760 3354 1762
rect 3346 1756 3348 1760
rect 3352 1756 3354 1760
rect 3346 1754 3354 1756
rect 3370 1760 3378 1762
rect 3370 1756 3372 1760
rect 3376 1756 3378 1760
rect 3370 1754 3378 1756
rect 3394 1760 3402 1762
rect 3394 1756 3396 1760
rect 3400 1756 3402 1760
rect 3394 1754 3402 1756
rect 3418 1760 3426 1762
rect 3418 1756 3420 1760
rect 3424 1756 3426 1760
rect 3418 1754 3426 1756
rect 3442 1760 3450 1762
rect 3442 1756 3444 1760
rect 3448 1756 3450 1760
rect 3442 1754 3450 1756
rect 3466 1760 3474 1762
rect 3466 1756 3468 1760
rect 3472 1756 3474 1760
rect 3466 1754 3474 1756
rect 3490 1760 3498 1762
rect 3490 1756 3492 1760
rect 3496 1756 3498 1760
rect 3490 1754 3498 1756
rect 3514 1760 3522 1762
rect 3514 1756 3516 1760
rect 3520 1756 3522 1760
rect 3514 1754 3522 1756
rect 3538 1760 3546 1762
rect 3538 1756 3540 1760
rect 3544 1756 3546 1760
rect 3538 1754 3546 1756
rect 3562 1760 3570 1762
rect 3562 1756 3564 1760
rect 3568 1756 3570 1760
rect 3562 1754 3570 1756
rect 3586 1760 3594 1762
rect 3586 1756 3588 1760
rect 3592 1756 3594 1760
rect 3586 1754 3594 1756
rect 3610 1760 3618 1762
rect 3610 1756 3612 1760
rect 3616 1756 3618 1760
rect 3610 1754 3618 1756
rect 3634 1760 3642 1762
rect 3634 1756 3636 1760
rect 3640 1756 3642 1760
rect 3634 1754 3642 1756
rect 3658 1760 3666 1762
rect 3658 1756 3660 1760
rect 3664 1756 3666 1760
rect 3658 1754 3666 1756
rect 3682 1760 3690 1762
rect 3682 1756 3684 1760
rect 3688 1756 3690 1760
rect 3682 1754 3690 1756
rect 3898 1760 3906 1762
rect 3898 1756 3900 1760
rect 3904 1756 3906 1760
rect 3898 1754 3906 1756
rect 3922 1760 3930 1762
rect 3922 1756 3924 1760
rect 3928 1756 3930 1760
rect 3922 1754 3930 1756
rect 3946 1760 3954 1762
rect 3946 1756 3948 1760
rect 3952 1756 3954 1760
rect 3946 1754 3954 1756
rect 3970 1760 3978 1762
rect 3970 1756 3972 1760
rect 3976 1756 3978 1760
rect 3970 1754 3978 1756
rect 3994 1760 4002 1762
rect 3994 1756 3996 1760
rect 4000 1756 4002 1760
rect 3994 1754 4002 1756
rect 4018 1760 4026 1762
rect 4018 1756 4020 1760
rect 4024 1756 4026 1760
rect 4018 1754 4026 1756
rect 4042 1760 4050 1762
rect 4042 1756 4044 1760
rect 4048 1756 4050 1760
rect 4042 1754 4050 1756
rect 4066 1760 4074 1762
rect 4066 1756 4068 1760
rect 4072 1756 4074 1760
rect 4066 1754 4074 1756
rect 4090 1760 4098 1762
rect 4090 1756 4092 1760
rect 4096 1756 4098 1760
rect 4090 1754 4098 1756
rect 4114 1760 4122 1762
rect 4114 1756 4116 1760
rect 4120 1756 4122 1760
rect 4114 1754 4122 1756
rect 4138 1760 4146 1762
rect 4138 1756 4140 1760
rect 4144 1756 4146 1760
rect 4138 1754 4146 1756
rect 4162 1760 4170 1762
rect 4162 1756 4164 1760
rect 4168 1756 4170 1760
rect 4162 1754 4170 1756
rect 4186 1760 4194 1762
rect 4186 1756 4188 1760
rect 4192 1756 4194 1760
rect 4186 1754 4194 1756
rect 4210 1760 4218 1762
rect 4210 1756 4212 1760
rect 4216 1756 4218 1760
rect 4210 1754 4218 1756
rect 4234 1760 4242 1762
rect 4234 1756 4236 1760
rect 4240 1756 4242 1760
rect 4234 1754 4242 1756
rect 4258 1760 4266 1762
rect 4258 1756 4260 1760
rect 4264 1756 4266 1760
rect 4258 1754 4266 1756
rect 4282 1760 4290 1762
rect 4282 1756 4284 1760
rect 4288 1756 4290 1760
rect 4282 1754 4290 1756
rect 4498 1760 4506 1762
rect 4498 1756 4500 1760
rect 4504 1756 4506 1760
rect 4498 1754 4506 1756
rect 4522 1760 4530 1762
rect 4522 1756 4524 1760
rect 4528 1756 4530 1760
rect 4522 1754 4530 1756
rect 4546 1760 4554 1762
rect 4546 1756 4548 1760
rect 4552 1756 4554 1760
rect 4546 1754 4554 1756
rect 4570 1760 4578 1762
rect 4570 1756 4572 1760
rect 4576 1756 4578 1760
rect 4570 1754 4578 1756
rect 4594 1760 4602 1762
rect 4594 1756 4596 1760
rect 4600 1756 4602 1760
rect 4594 1754 4602 1756
rect 4618 1760 4626 1762
rect 4618 1756 4620 1760
rect 4624 1756 4626 1760
rect 4618 1754 4626 1756
rect 4642 1760 4650 1762
rect 4642 1756 4644 1760
rect 4648 1756 4650 1760
rect 4642 1754 4650 1756
rect 4666 1760 4674 1762
rect 4666 1756 4668 1760
rect 4672 1756 4674 1760
rect 4666 1754 4674 1756
rect 4690 1760 4698 1762
rect 4690 1756 4692 1760
rect 4696 1756 4698 1760
rect 4690 1754 4698 1756
rect 4714 1760 4722 1762
rect 4714 1756 4716 1760
rect 4720 1756 4722 1760
rect 4714 1754 4722 1756
rect 4738 1760 4746 1762
rect 4738 1756 4740 1760
rect 4744 1756 4746 1760
rect 4738 1754 4746 1756
rect 4762 1760 4770 1762
rect 4762 1756 4764 1760
rect 4768 1756 4770 1760
rect 4762 1754 4770 1756
rect 4786 1760 4794 1762
rect 4786 1756 4788 1760
rect 4792 1756 4794 1760
rect 4786 1754 4794 1756
rect 5698 1760 5706 1762
rect 5698 1756 5700 1760
rect 5704 1756 5706 1760
rect 5698 1754 5706 1756
rect 5722 1760 5730 1762
rect 5722 1756 5724 1760
rect 5728 1756 5730 1760
rect 5722 1754 5730 1756
rect 5746 1760 5754 1762
rect 5746 1756 5748 1760
rect 5752 1756 5754 1760
rect 5746 1754 5754 1756
rect 5770 1760 5778 1762
rect 5770 1756 5772 1760
rect 5776 1756 5778 1760
rect 5770 1754 5778 1756
rect 5794 1760 5802 1762
rect 5794 1756 5796 1760
rect 5800 1756 5802 1760
rect 5794 1754 5802 1756
rect 5818 1760 5826 1762
rect 5818 1756 5820 1760
rect 5824 1756 5826 1760
rect 5818 1754 5826 1756
rect 5842 1760 5850 1762
rect 5842 1756 5844 1760
rect 5848 1756 5850 1760
rect 5842 1754 5850 1756
rect 5866 1760 5874 1762
rect 5866 1756 5868 1760
rect 5872 1756 5874 1760
rect 5866 1754 5874 1756
rect 5890 1760 5898 1762
rect 5890 1756 5892 1760
rect 5896 1756 5898 1760
rect 5890 1754 5898 1756
rect 5914 1760 5922 1762
rect 5914 1756 5916 1760
rect 5920 1756 5922 1760
rect 5914 1754 5922 1756
rect 5938 1760 5946 1762
rect 5938 1756 5940 1760
rect 5944 1756 5946 1760
rect 5938 1754 5946 1756
rect 5962 1760 5970 1762
rect 5962 1756 5964 1760
rect 5968 1756 5970 1760
rect 5962 1754 5970 1756
rect 5986 1760 5994 1762
rect 5986 1756 5988 1760
rect 5992 1756 5994 1760
rect 5986 1754 5994 1756
rect 6010 1760 6018 1762
rect 6010 1756 6012 1760
rect 6016 1756 6018 1760
rect 6010 1754 6018 1756
rect 6034 1760 6042 1762
rect 6034 1756 6036 1760
rect 6040 1756 6042 1760
rect 6034 1754 6042 1756
rect 6058 1760 6066 1762
rect 6058 1756 6060 1760
rect 6064 1756 6066 1760
rect 6058 1754 6066 1756
rect 6082 1760 6090 1762
rect 6082 1756 6084 1760
rect 6088 1756 6090 1760
rect 6082 1754 6090 1756
rect 6298 1760 6306 1762
rect 6298 1756 6300 1760
rect 6304 1756 6306 1760
rect 6298 1754 6306 1756
rect 6322 1760 6330 1762
rect 6322 1756 6324 1760
rect 6328 1756 6330 1760
rect 6322 1754 6330 1756
rect 6346 1760 6354 1762
rect 6346 1756 6348 1760
rect 6352 1756 6354 1760
rect 6346 1754 6354 1756
rect 6370 1760 6378 1762
rect 6370 1756 6372 1760
rect 6376 1756 6378 1760
rect 6370 1754 6378 1756
rect 6394 1760 6402 1762
rect 6394 1756 6396 1760
rect 6400 1756 6402 1760
rect 6394 1754 6402 1756
rect 6418 1760 6426 1762
rect 6418 1756 6420 1760
rect 6424 1756 6426 1760
rect 6418 1754 6426 1756
rect 6442 1760 6450 1762
rect 6442 1756 6444 1760
rect 6448 1756 6450 1760
rect 6442 1754 6450 1756
rect 6466 1760 6474 1762
rect 6466 1756 6468 1760
rect 6472 1756 6474 1760
rect 6466 1754 6474 1756
rect 6490 1760 6498 1762
rect 6490 1756 6492 1760
rect 6496 1756 6498 1760
rect 6490 1754 6498 1756
rect 6514 1760 6522 1762
rect 6514 1756 6516 1760
rect 6520 1756 6522 1760
rect 6514 1754 6522 1756
rect 6538 1760 6546 1762
rect 6538 1756 6540 1760
rect 6544 1756 6546 1760
rect 6538 1754 6546 1756
rect 6562 1760 6570 1762
rect 6562 1756 6564 1760
rect 6568 1756 6570 1760
rect 6562 1754 6570 1756
rect 6586 1760 6594 1762
rect 6586 1756 6588 1760
rect 6592 1756 6594 1760
rect 6586 1754 6594 1756
rect 6610 1760 6618 1762
rect 6610 1756 6612 1760
rect 6616 1756 6618 1760
rect 6610 1754 6618 1756
rect 6634 1760 6642 1762
rect 6634 1756 6636 1760
rect 6640 1756 6642 1760
rect 6634 1754 6642 1756
rect 6658 1760 6666 1762
rect 6658 1756 6660 1760
rect 6664 1756 6666 1760
rect 6658 1754 6666 1756
rect 6682 1760 6690 1762
rect 6682 1756 6684 1760
rect 6688 1756 6690 1760
rect 6682 1754 6690 1756
rect 6898 1760 6906 1762
rect 6898 1756 6900 1760
rect 6904 1756 6906 1760
rect 6898 1754 6906 1756
rect 6922 1760 6930 1762
rect 6922 1756 6924 1760
rect 6928 1756 6930 1760
rect 6922 1754 6930 1756
rect 6946 1760 6954 1762
rect 6946 1756 6948 1760
rect 6952 1756 6954 1760
rect 6946 1754 6954 1756
rect 6970 1760 6978 1762
rect 6970 1756 6972 1760
rect 6976 1756 6978 1760
rect 6970 1754 6978 1756
rect 6994 1760 7002 1762
rect 6994 1756 6996 1760
rect 7000 1756 7002 1760
rect 6994 1754 7002 1756
rect 7018 1760 7026 1762
rect 7018 1756 7020 1760
rect 7024 1756 7026 1760
rect 7018 1754 7026 1756
rect 7042 1760 7050 1762
rect 7042 1756 7044 1760
rect 7048 1756 7050 1760
rect 7042 1754 7050 1756
rect 7066 1760 7074 1762
rect 7066 1756 7068 1760
rect 7072 1756 7074 1760
rect 7066 1754 7074 1756
rect 7090 1760 7098 1762
rect 7090 1756 7092 1760
rect 7096 1756 7098 1760
rect 7090 1754 7098 1756
rect 7114 1760 7122 1762
rect 7114 1756 7116 1760
rect 7120 1756 7122 1760
rect 7114 1754 7122 1756
rect 7138 1760 7146 1762
rect 7138 1756 7140 1760
rect 7144 1756 7146 1760
rect 7138 1754 7146 1756
rect 7162 1760 7170 1762
rect 7162 1756 7164 1760
rect 7168 1756 7170 1760
rect 7162 1754 7170 1756
rect 7186 1760 7194 1762
rect 7186 1756 7188 1760
rect 7192 1756 7194 1760
rect 7186 1754 7194 1756
rect 2400 1748 2406 1750
rect 2404 1744 2406 1748
rect 2400 1742 2406 1744
rect 2422 1748 2430 1750
rect 2422 1744 2424 1748
rect 2428 1744 2430 1748
rect 2422 1742 2430 1744
rect 2446 1748 2454 1750
rect 2446 1744 2448 1748
rect 2452 1744 2454 1748
rect 2446 1742 2454 1744
rect 2470 1748 2478 1750
rect 2470 1744 2472 1748
rect 2476 1744 2478 1748
rect 2470 1742 2478 1744
rect 2494 1748 2502 1750
rect 2494 1744 2496 1748
rect 2500 1744 2502 1748
rect 2494 1742 2502 1744
rect 2710 1748 2718 1750
rect 2710 1744 2712 1748
rect 2716 1744 2718 1748
rect 2710 1742 2718 1744
rect 2734 1748 2742 1750
rect 2734 1744 2736 1748
rect 2740 1744 2742 1748
rect 2734 1742 2742 1744
rect 2758 1748 2766 1750
rect 2758 1744 2760 1748
rect 2764 1744 2766 1748
rect 2758 1742 2766 1744
rect 2782 1748 2790 1750
rect 2782 1744 2784 1748
rect 2788 1744 2790 1748
rect 2782 1742 2790 1744
rect 2806 1748 2814 1750
rect 2806 1744 2808 1748
rect 2812 1744 2814 1748
rect 2806 1742 2814 1744
rect 2830 1748 2838 1750
rect 2830 1744 2832 1748
rect 2836 1744 2838 1748
rect 2830 1742 2838 1744
rect 2854 1748 2862 1750
rect 2854 1744 2856 1748
rect 2860 1744 2862 1748
rect 2854 1742 2862 1744
rect 2878 1748 2886 1750
rect 2878 1744 2880 1748
rect 2884 1744 2886 1748
rect 2878 1742 2886 1744
rect 2902 1748 2910 1750
rect 2902 1744 2904 1748
rect 2908 1744 2910 1748
rect 2902 1742 2910 1744
rect 2926 1748 2934 1750
rect 2926 1744 2928 1748
rect 2932 1744 2934 1748
rect 2926 1742 2934 1744
rect 2950 1748 2958 1750
rect 2950 1744 2952 1748
rect 2956 1744 2958 1748
rect 2950 1742 2958 1744
rect 2974 1748 2982 1750
rect 2974 1744 2976 1748
rect 2980 1744 2982 1748
rect 2974 1742 2982 1744
rect 2998 1748 3006 1750
rect 2998 1744 3000 1748
rect 3004 1744 3006 1748
rect 2998 1742 3006 1744
rect 3022 1748 3030 1750
rect 3022 1744 3024 1748
rect 3028 1744 3030 1748
rect 3022 1742 3030 1744
rect 3046 1748 3054 1750
rect 3046 1744 3048 1748
rect 3052 1744 3054 1748
rect 3046 1742 3054 1744
rect 3070 1748 3078 1750
rect 3070 1744 3072 1748
rect 3076 1744 3078 1748
rect 3070 1742 3078 1744
rect 3094 1748 3102 1750
rect 3094 1744 3096 1748
rect 3100 1744 3102 1748
rect 3094 1742 3102 1744
rect 3310 1748 3318 1750
rect 3310 1744 3312 1748
rect 3316 1744 3318 1748
rect 3310 1742 3318 1744
rect 3334 1748 3342 1750
rect 3334 1744 3336 1748
rect 3340 1744 3342 1748
rect 3334 1742 3342 1744
rect 3358 1748 3366 1750
rect 3358 1744 3360 1748
rect 3364 1744 3366 1748
rect 3358 1742 3366 1744
rect 3382 1748 3390 1750
rect 3382 1744 3384 1748
rect 3388 1744 3390 1748
rect 3382 1742 3390 1744
rect 3406 1748 3414 1750
rect 3406 1744 3408 1748
rect 3412 1744 3414 1748
rect 3406 1742 3414 1744
rect 3430 1748 3438 1750
rect 3430 1744 3432 1748
rect 3436 1744 3438 1748
rect 3430 1742 3438 1744
rect 3454 1748 3462 1750
rect 3454 1744 3456 1748
rect 3460 1744 3462 1748
rect 3454 1742 3462 1744
rect 3478 1748 3486 1750
rect 3478 1744 3480 1748
rect 3484 1744 3486 1748
rect 3478 1742 3486 1744
rect 3502 1748 3510 1750
rect 3502 1744 3504 1748
rect 3508 1744 3510 1748
rect 3502 1742 3510 1744
rect 3526 1748 3534 1750
rect 3526 1744 3528 1748
rect 3532 1744 3534 1748
rect 3526 1742 3534 1744
rect 3550 1748 3558 1750
rect 3550 1744 3552 1748
rect 3556 1744 3558 1748
rect 3550 1742 3558 1744
rect 3574 1748 3582 1750
rect 3574 1744 3576 1748
rect 3580 1744 3582 1748
rect 3574 1742 3582 1744
rect 3598 1748 3606 1750
rect 3598 1744 3600 1748
rect 3604 1744 3606 1748
rect 3598 1742 3606 1744
rect 3622 1748 3630 1750
rect 3622 1744 3624 1748
rect 3628 1744 3630 1748
rect 3622 1742 3630 1744
rect 3646 1748 3654 1750
rect 3646 1744 3648 1748
rect 3652 1744 3654 1748
rect 3646 1742 3654 1744
rect 3670 1748 3678 1750
rect 3670 1744 3672 1748
rect 3676 1744 3678 1748
rect 3670 1742 3678 1744
rect 3694 1748 3702 1750
rect 3694 1744 3696 1748
rect 3700 1744 3702 1748
rect 3694 1742 3702 1744
rect 3910 1748 3918 1750
rect 3910 1744 3912 1748
rect 3916 1744 3918 1748
rect 3910 1742 3918 1744
rect 3934 1748 3942 1750
rect 3934 1744 3936 1748
rect 3940 1744 3942 1748
rect 3934 1742 3942 1744
rect 3958 1748 3966 1750
rect 3958 1744 3960 1748
rect 3964 1744 3966 1748
rect 3958 1742 3966 1744
rect 3982 1748 3990 1750
rect 3982 1744 3984 1748
rect 3988 1744 3990 1748
rect 3982 1742 3990 1744
rect 4006 1748 4014 1750
rect 4006 1744 4008 1748
rect 4012 1744 4014 1748
rect 4006 1742 4014 1744
rect 4030 1748 4038 1750
rect 4030 1744 4032 1748
rect 4036 1744 4038 1748
rect 4030 1742 4038 1744
rect 4054 1748 4062 1750
rect 4054 1744 4056 1748
rect 4060 1744 4062 1748
rect 4054 1742 4062 1744
rect 4078 1748 4086 1750
rect 4078 1744 4080 1748
rect 4084 1744 4086 1748
rect 4078 1742 4086 1744
rect 4102 1748 4110 1750
rect 4102 1744 4104 1748
rect 4108 1744 4110 1748
rect 4102 1742 4110 1744
rect 4126 1748 4134 1750
rect 4126 1744 4128 1748
rect 4132 1744 4134 1748
rect 4126 1742 4134 1744
rect 4150 1748 4158 1750
rect 4150 1744 4152 1748
rect 4156 1744 4158 1748
rect 4150 1742 4158 1744
rect 4174 1748 4182 1750
rect 4174 1744 4176 1748
rect 4180 1744 4182 1748
rect 4174 1742 4182 1744
rect 4198 1748 4206 1750
rect 4198 1744 4200 1748
rect 4204 1744 4206 1748
rect 4198 1742 4206 1744
rect 4222 1748 4230 1750
rect 4222 1744 4224 1748
rect 4228 1744 4230 1748
rect 4222 1742 4230 1744
rect 4246 1748 4254 1750
rect 4246 1744 4248 1748
rect 4252 1744 4254 1748
rect 4246 1742 4254 1744
rect 4270 1748 4278 1750
rect 4270 1744 4272 1748
rect 4276 1744 4278 1748
rect 4270 1742 4278 1744
rect 4294 1748 4302 1750
rect 4294 1744 4296 1748
rect 4300 1744 4302 1748
rect 4294 1742 4302 1744
rect 4510 1748 4518 1750
rect 4510 1744 4512 1748
rect 4516 1744 4518 1748
rect 4510 1742 4518 1744
rect 4534 1748 4542 1750
rect 4534 1744 4536 1748
rect 4540 1744 4542 1748
rect 4534 1742 4542 1744
rect 4558 1748 4566 1750
rect 4558 1744 4560 1748
rect 4564 1744 4566 1748
rect 4558 1742 4566 1744
rect 4582 1748 4590 1750
rect 4582 1744 4584 1748
rect 4588 1744 4590 1748
rect 4582 1742 4590 1744
rect 4606 1748 4614 1750
rect 4606 1744 4608 1748
rect 4612 1744 4614 1748
rect 4606 1742 4614 1744
rect 4630 1748 4638 1750
rect 4630 1744 4632 1748
rect 4636 1744 4638 1748
rect 4630 1742 4638 1744
rect 4654 1748 4662 1750
rect 4654 1744 4656 1748
rect 4660 1744 4662 1748
rect 4654 1742 4662 1744
rect 4678 1748 4686 1750
rect 4678 1744 4680 1748
rect 4684 1744 4686 1748
rect 4678 1742 4686 1744
rect 4702 1748 4710 1750
rect 4702 1744 4704 1748
rect 4708 1744 4710 1748
rect 4702 1742 4710 1744
rect 4726 1748 4734 1750
rect 4726 1744 4728 1748
rect 4732 1744 4734 1748
rect 4726 1742 4734 1744
rect 4750 1748 4758 1750
rect 4750 1744 4752 1748
rect 4756 1744 4758 1748
rect 4750 1742 4758 1744
rect 4774 1748 4782 1750
rect 4774 1744 4776 1748
rect 4780 1744 4782 1748
rect 4774 1742 4782 1744
rect 4798 1742 4800 1750
rect 5710 1748 5718 1750
rect 5710 1744 5712 1748
rect 5716 1744 5718 1748
rect 5710 1742 5718 1744
rect 5734 1748 5742 1750
rect 5734 1744 5736 1748
rect 5740 1744 5742 1748
rect 5734 1742 5742 1744
rect 5758 1748 5766 1750
rect 5758 1744 5760 1748
rect 5764 1744 5766 1748
rect 5758 1742 5766 1744
rect 5782 1748 5790 1750
rect 5782 1744 5784 1748
rect 5788 1744 5790 1748
rect 5782 1742 5790 1744
rect 5806 1748 5814 1750
rect 5806 1744 5808 1748
rect 5812 1744 5814 1748
rect 5806 1742 5814 1744
rect 5830 1748 5838 1750
rect 5830 1744 5832 1748
rect 5836 1744 5838 1748
rect 5830 1742 5838 1744
rect 5854 1748 5862 1750
rect 5854 1744 5856 1748
rect 5860 1744 5862 1748
rect 5854 1742 5862 1744
rect 5878 1748 5886 1750
rect 5878 1744 5880 1748
rect 5884 1744 5886 1748
rect 5878 1742 5886 1744
rect 5902 1748 5910 1750
rect 5902 1744 5904 1748
rect 5908 1744 5910 1748
rect 5902 1742 5910 1744
rect 5926 1748 5934 1750
rect 5926 1744 5928 1748
rect 5932 1744 5934 1748
rect 5926 1742 5934 1744
rect 5950 1748 5958 1750
rect 5950 1744 5952 1748
rect 5956 1744 5958 1748
rect 5950 1742 5958 1744
rect 5974 1748 5982 1750
rect 5974 1744 5976 1748
rect 5980 1744 5982 1748
rect 5974 1742 5982 1744
rect 5998 1748 6006 1750
rect 5998 1744 6000 1748
rect 6004 1744 6006 1748
rect 5998 1742 6006 1744
rect 6022 1748 6030 1750
rect 6022 1744 6024 1748
rect 6028 1744 6030 1748
rect 6022 1742 6030 1744
rect 6046 1748 6054 1750
rect 6046 1744 6048 1748
rect 6052 1744 6054 1748
rect 6046 1742 6054 1744
rect 6070 1748 6078 1750
rect 6070 1744 6072 1748
rect 6076 1744 6078 1748
rect 6070 1742 6078 1744
rect 6094 1748 6102 1750
rect 6094 1744 6096 1748
rect 6100 1744 6102 1748
rect 6094 1742 6102 1744
rect 6310 1748 6318 1750
rect 6310 1744 6312 1748
rect 6316 1744 6318 1748
rect 6310 1742 6318 1744
rect 6334 1748 6342 1750
rect 6334 1744 6336 1748
rect 6340 1744 6342 1748
rect 6334 1742 6342 1744
rect 6358 1748 6366 1750
rect 6358 1744 6360 1748
rect 6364 1744 6366 1748
rect 6358 1742 6366 1744
rect 6382 1748 6390 1750
rect 6382 1744 6384 1748
rect 6388 1744 6390 1748
rect 6382 1742 6390 1744
rect 6406 1748 6414 1750
rect 6406 1744 6408 1748
rect 6412 1744 6414 1748
rect 6406 1742 6414 1744
rect 6430 1748 6438 1750
rect 6430 1744 6432 1748
rect 6436 1744 6438 1748
rect 6430 1742 6438 1744
rect 6454 1748 6462 1750
rect 6454 1744 6456 1748
rect 6460 1744 6462 1748
rect 6454 1742 6462 1744
rect 6478 1748 6486 1750
rect 6478 1744 6480 1748
rect 6484 1744 6486 1748
rect 6478 1742 6486 1744
rect 6502 1748 6510 1750
rect 6502 1744 6504 1748
rect 6508 1744 6510 1748
rect 6502 1742 6510 1744
rect 6526 1748 6534 1750
rect 6526 1744 6528 1748
rect 6532 1744 6534 1748
rect 6526 1742 6534 1744
rect 6550 1748 6558 1750
rect 6550 1744 6552 1748
rect 6556 1744 6558 1748
rect 6550 1742 6558 1744
rect 6574 1748 6582 1750
rect 6574 1744 6576 1748
rect 6580 1744 6582 1748
rect 6574 1742 6582 1744
rect 6598 1748 6606 1750
rect 6598 1744 6600 1748
rect 6604 1744 6606 1748
rect 6598 1742 6606 1744
rect 6622 1748 6630 1750
rect 6622 1744 6624 1748
rect 6628 1744 6630 1748
rect 6622 1742 6630 1744
rect 6646 1748 6654 1750
rect 6646 1744 6648 1748
rect 6652 1744 6654 1748
rect 6646 1742 6654 1744
rect 6670 1748 6678 1750
rect 6670 1744 6672 1748
rect 6676 1744 6678 1748
rect 6670 1742 6678 1744
rect 6694 1748 6702 1750
rect 6694 1744 6696 1748
rect 6700 1744 6702 1748
rect 6694 1742 6702 1744
rect 6910 1748 6918 1750
rect 6910 1744 6912 1748
rect 6916 1744 6918 1748
rect 6910 1742 6918 1744
rect 6934 1748 6942 1750
rect 6934 1744 6936 1748
rect 6940 1744 6942 1748
rect 6934 1742 6942 1744
rect 6958 1748 6966 1750
rect 6958 1744 6960 1748
rect 6964 1744 6966 1748
rect 6958 1742 6966 1744
rect 6982 1748 6990 1750
rect 6982 1744 6984 1748
rect 6988 1744 6990 1748
rect 6982 1742 6990 1744
rect 7006 1748 7014 1750
rect 7006 1744 7008 1748
rect 7012 1744 7014 1748
rect 7006 1742 7014 1744
rect 7030 1748 7038 1750
rect 7030 1744 7032 1748
rect 7036 1744 7038 1748
rect 7030 1742 7038 1744
rect 7054 1748 7062 1750
rect 7054 1744 7056 1748
rect 7060 1744 7062 1748
rect 7054 1742 7062 1744
rect 7078 1748 7086 1750
rect 7078 1744 7080 1748
rect 7084 1744 7086 1748
rect 7078 1742 7086 1744
rect 7102 1748 7110 1750
rect 7102 1744 7104 1748
rect 7108 1744 7110 1748
rect 7102 1742 7110 1744
rect 7126 1748 7134 1750
rect 7126 1744 7128 1748
rect 7132 1744 7134 1748
rect 7126 1742 7134 1744
rect 7150 1748 7158 1750
rect 7150 1744 7152 1748
rect 7156 1744 7158 1748
rect 7150 1742 7158 1744
rect 7174 1748 7182 1750
rect 7174 1744 7176 1748
rect 7180 1744 7182 1748
rect 7174 1742 7182 1744
rect 7198 1742 7200 1750
rect 2410 1736 2418 1738
rect 2410 1732 2412 1736
rect 2416 1732 2418 1736
rect 2410 1730 2418 1732
rect 2434 1736 2442 1738
rect 2434 1732 2436 1736
rect 2440 1732 2442 1736
rect 2434 1730 2442 1732
rect 2458 1736 2466 1738
rect 2458 1732 2460 1736
rect 2464 1732 2466 1736
rect 2458 1730 2466 1732
rect 2482 1736 2490 1738
rect 2482 1732 2484 1736
rect 2488 1732 2490 1736
rect 2482 1730 2490 1732
rect 2698 1736 2706 1738
rect 2698 1732 2700 1736
rect 2704 1732 2706 1736
rect 2698 1730 2706 1732
rect 2722 1736 2730 1738
rect 2722 1732 2724 1736
rect 2728 1732 2730 1736
rect 2722 1730 2730 1732
rect 2746 1736 2754 1738
rect 2746 1732 2748 1736
rect 2752 1732 2754 1736
rect 2746 1730 2754 1732
rect 2770 1736 2778 1738
rect 2770 1732 2772 1736
rect 2776 1732 2778 1736
rect 2770 1730 2778 1732
rect 2794 1736 2802 1738
rect 2794 1732 2796 1736
rect 2800 1732 2802 1736
rect 2794 1730 2802 1732
rect 2818 1736 2826 1738
rect 2818 1732 2820 1736
rect 2824 1732 2826 1736
rect 2818 1730 2826 1732
rect 2842 1736 2850 1738
rect 2842 1732 2844 1736
rect 2848 1732 2850 1736
rect 2842 1730 2850 1732
rect 2866 1736 2874 1738
rect 2866 1732 2868 1736
rect 2872 1732 2874 1736
rect 2866 1730 2874 1732
rect 2890 1736 2898 1738
rect 2890 1732 2892 1736
rect 2896 1732 2898 1736
rect 2890 1730 2898 1732
rect 2914 1736 2922 1738
rect 2914 1732 2916 1736
rect 2920 1732 2922 1736
rect 2914 1730 2922 1732
rect 2938 1736 2946 1738
rect 2938 1732 2940 1736
rect 2944 1732 2946 1736
rect 2938 1730 2946 1732
rect 2962 1736 2970 1738
rect 2962 1732 2964 1736
rect 2968 1732 2970 1736
rect 2962 1730 2970 1732
rect 2986 1736 2994 1738
rect 2986 1732 2988 1736
rect 2992 1732 2994 1736
rect 2986 1730 2994 1732
rect 3010 1736 3018 1738
rect 3010 1732 3012 1736
rect 3016 1732 3018 1736
rect 3010 1730 3018 1732
rect 3034 1736 3042 1738
rect 3034 1732 3036 1736
rect 3040 1732 3042 1736
rect 3034 1730 3042 1732
rect 3058 1736 3066 1738
rect 3058 1732 3060 1736
rect 3064 1732 3066 1736
rect 3058 1730 3066 1732
rect 3082 1736 3090 1738
rect 3082 1732 3084 1736
rect 3088 1732 3090 1736
rect 3082 1730 3090 1732
rect 3298 1736 3306 1738
rect 3298 1732 3300 1736
rect 3304 1732 3306 1736
rect 3298 1730 3306 1732
rect 3322 1736 3330 1738
rect 3322 1732 3324 1736
rect 3328 1732 3330 1736
rect 3322 1730 3330 1732
rect 3346 1736 3354 1738
rect 3346 1732 3348 1736
rect 3352 1732 3354 1736
rect 3346 1730 3354 1732
rect 3370 1736 3378 1738
rect 3370 1732 3372 1736
rect 3376 1732 3378 1736
rect 3370 1730 3378 1732
rect 3394 1736 3402 1738
rect 3394 1732 3396 1736
rect 3400 1732 3402 1736
rect 3394 1730 3402 1732
rect 3418 1736 3426 1738
rect 3418 1732 3420 1736
rect 3424 1732 3426 1736
rect 3418 1730 3426 1732
rect 3442 1736 3450 1738
rect 3442 1732 3444 1736
rect 3448 1732 3450 1736
rect 3442 1730 3450 1732
rect 3466 1736 3474 1738
rect 3466 1732 3468 1736
rect 3472 1732 3474 1736
rect 3466 1730 3474 1732
rect 3490 1736 3498 1738
rect 3490 1732 3492 1736
rect 3496 1732 3498 1736
rect 3490 1730 3498 1732
rect 3514 1736 3522 1738
rect 3514 1732 3516 1736
rect 3520 1732 3522 1736
rect 3514 1730 3522 1732
rect 3538 1736 3546 1738
rect 3538 1732 3540 1736
rect 3544 1732 3546 1736
rect 3538 1730 3546 1732
rect 3562 1736 3570 1738
rect 3562 1732 3564 1736
rect 3568 1732 3570 1736
rect 3562 1730 3570 1732
rect 3586 1736 3594 1738
rect 3586 1732 3588 1736
rect 3592 1732 3594 1736
rect 3586 1730 3594 1732
rect 3610 1736 3618 1738
rect 3610 1732 3612 1736
rect 3616 1732 3618 1736
rect 3610 1730 3618 1732
rect 3634 1736 3642 1738
rect 3634 1732 3636 1736
rect 3640 1732 3642 1736
rect 3634 1730 3642 1732
rect 3658 1736 3666 1738
rect 3658 1732 3660 1736
rect 3664 1732 3666 1736
rect 3658 1730 3666 1732
rect 3682 1736 3690 1738
rect 3682 1732 3684 1736
rect 3688 1732 3690 1736
rect 3682 1730 3690 1732
rect 3898 1736 3906 1738
rect 3898 1732 3900 1736
rect 3904 1732 3906 1736
rect 3898 1730 3906 1732
rect 3922 1736 3930 1738
rect 3922 1732 3924 1736
rect 3928 1732 3930 1736
rect 3922 1730 3930 1732
rect 3946 1736 3954 1738
rect 3946 1732 3948 1736
rect 3952 1732 3954 1736
rect 3946 1730 3954 1732
rect 3970 1736 3978 1738
rect 3970 1732 3972 1736
rect 3976 1732 3978 1736
rect 3970 1730 3978 1732
rect 3994 1736 4002 1738
rect 3994 1732 3996 1736
rect 4000 1732 4002 1736
rect 3994 1730 4002 1732
rect 4018 1736 4026 1738
rect 4018 1732 4020 1736
rect 4024 1732 4026 1736
rect 4018 1730 4026 1732
rect 4042 1736 4050 1738
rect 4042 1732 4044 1736
rect 4048 1732 4050 1736
rect 4042 1730 4050 1732
rect 4066 1736 4074 1738
rect 4066 1732 4068 1736
rect 4072 1732 4074 1736
rect 4066 1730 4074 1732
rect 4090 1736 4098 1738
rect 4090 1732 4092 1736
rect 4096 1732 4098 1736
rect 4090 1730 4098 1732
rect 4114 1736 4122 1738
rect 4114 1732 4116 1736
rect 4120 1732 4122 1736
rect 4114 1730 4122 1732
rect 4138 1736 4146 1738
rect 4138 1732 4140 1736
rect 4144 1732 4146 1736
rect 4138 1730 4146 1732
rect 4162 1736 4170 1738
rect 4162 1732 4164 1736
rect 4168 1732 4170 1736
rect 4162 1730 4170 1732
rect 4186 1736 4194 1738
rect 4186 1732 4188 1736
rect 4192 1732 4194 1736
rect 4186 1730 4194 1732
rect 4210 1736 4218 1738
rect 4210 1732 4212 1736
rect 4216 1732 4218 1736
rect 4210 1730 4218 1732
rect 4234 1736 4242 1738
rect 4234 1732 4236 1736
rect 4240 1732 4242 1736
rect 4234 1730 4242 1732
rect 4258 1736 4266 1738
rect 4258 1732 4260 1736
rect 4264 1732 4266 1736
rect 4258 1730 4266 1732
rect 4282 1736 4290 1738
rect 4282 1732 4284 1736
rect 4288 1732 4290 1736
rect 4282 1730 4290 1732
rect 4498 1736 4506 1738
rect 4498 1732 4500 1736
rect 4504 1732 4506 1736
rect 4498 1730 4506 1732
rect 4522 1736 4530 1738
rect 4522 1732 4524 1736
rect 4528 1732 4530 1736
rect 4522 1730 4530 1732
rect 4546 1736 4554 1738
rect 4546 1732 4548 1736
rect 4552 1732 4554 1736
rect 4546 1730 4554 1732
rect 4570 1736 4578 1738
rect 4570 1732 4572 1736
rect 4576 1732 4578 1736
rect 4570 1730 4578 1732
rect 4594 1736 4602 1738
rect 4594 1732 4596 1736
rect 4600 1732 4602 1736
rect 4594 1730 4602 1732
rect 4618 1736 4626 1738
rect 4618 1732 4620 1736
rect 4624 1732 4626 1736
rect 4618 1730 4626 1732
rect 4642 1736 4650 1738
rect 4642 1732 4644 1736
rect 4648 1732 4650 1736
rect 4642 1730 4650 1732
rect 4666 1736 4674 1738
rect 4666 1732 4668 1736
rect 4672 1732 4674 1736
rect 4666 1730 4674 1732
rect 4690 1736 4698 1738
rect 4690 1732 4692 1736
rect 4696 1732 4698 1736
rect 4690 1730 4698 1732
rect 4714 1736 4722 1738
rect 4714 1732 4716 1736
rect 4720 1732 4722 1736
rect 4714 1730 4722 1732
rect 4738 1736 4746 1738
rect 4738 1732 4740 1736
rect 4744 1732 4746 1736
rect 4738 1730 4746 1732
rect 4762 1736 4770 1738
rect 4762 1732 4764 1736
rect 4768 1732 4770 1736
rect 4762 1730 4770 1732
rect 4786 1736 4794 1738
rect 4786 1732 4788 1736
rect 4792 1732 4794 1736
rect 4786 1730 4794 1732
rect 5698 1736 5706 1738
rect 5698 1732 5700 1736
rect 5704 1732 5706 1736
rect 5698 1730 5706 1732
rect 5722 1736 5730 1738
rect 5722 1732 5724 1736
rect 5728 1732 5730 1736
rect 5722 1730 5730 1732
rect 5746 1736 5754 1738
rect 5746 1732 5748 1736
rect 5752 1732 5754 1736
rect 5746 1730 5754 1732
rect 5770 1736 5778 1738
rect 5770 1732 5772 1736
rect 5776 1732 5778 1736
rect 5770 1730 5778 1732
rect 5794 1736 5802 1738
rect 5794 1732 5796 1736
rect 5800 1732 5802 1736
rect 5794 1730 5802 1732
rect 5818 1736 5826 1738
rect 5818 1732 5820 1736
rect 5824 1732 5826 1736
rect 5818 1730 5826 1732
rect 5842 1736 5850 1738
rect 5842 1732 5844 1736
rect 5848 1732 5850 1736
rect 5842 1730 5850 1732
rect 5866 1736 5874 1738
rect 5866 1732 5868 1736
rect 5872 1732 5874 1736
rect 5866 1730 5874 1732
rect 5890 1736 5898 1738
rect 5890 1732 5892 1736
rect 5896 1732 5898 1736
rect 5890 1730 5898 1732
rect 5914 1736 5922 1738
rect 5914 1732 5916 1736
rect 5920 1732 5922 1736
rect 5914 1730 5922 1732
rect 5938 1736 5946 1738
rect 5938 1732 5940 1736
rect 5944 1732 5946 1736
rect 5938 1730 5946 1732
rect 5962 1736 5970 1738
rect 5962 1732 5964 1736
rect 5968 1732 5970 1736
rect 5962 1730 5970 1732
rect 5986 1736 5994 1738
rect 5986 1732 5988 1736
rect 5992 1732 5994 1736
rect 5986 1730 5994 1732
rect 6010 1736 6018 1738
rect 6010 1732 6012 1736
rect 6016 1732 6018 1736
rect 6010 1730 6018 1732
rect 6034 1736 6042 1738
rect 6034 1732 6036 1736
rect 6040 1732 6042 1736
rect 6034 1730 6042 1732
rect 6058 1736 6066 1738
rect 6058 1732 6060 1736
rect 6064 1732 6066 1736
rect 6058 1730 6066 1732
rect 6082 1736 6090 1738
rect 6082 1732 6084 1736
rect 6088 1732 6090 1736
rect 6082 1730 6090 1732
rect 6298 1736 6306 1738
rect 6298 1732 6300 1736
rect 6304 1732 6306 1736
rect 6298 1730 6306 1732
rect 6322 1736 6330 1738
rect 6322 1732 6324 1736
rect 6328 1732 6330 1736
rect 6322 1730 6330 1732
rect 6346 1736 6354 1738
rect 6346 1732 6348 1736
rect 6352 1732 6354 1736
rect 6346 1730 6354 1732
rect 6370 1736 6378 1738
rect 6370 1732 6372 1736
rect 6376 1732 6378 1736
rect 6370 1730 6378 1732
rect 6394 1736 6402 1738
rect 6394 1732 6396 1736
rect 6400 1732 6402 1736
rect 6394 1730 6402 1732
rect 6418 1736 6426 1738
rect 6418 1732 6420 1736
rect 6424 1732 6426 1736
rect 6418 1730 6426 1732
rect 6442 1736 6450 1738
rect 6442 1732 6444 1736
rect 6448 1732 6450 1736
rect 6442 1730 6450 1732
rect 6466 1736 6474 1738
rect 6466 1732 6468 1736
rect 6472 1732 6474 1736
rect 6466 1730 6474 1732
rect 6490 1736 6498 1738
rect 6490 1732 6492 1736
rect 6496 1732 6498 1736
rect 6490 1730 6498 1732
rect 6514 1736 6522 1738
rect 6514 1732 6516 1736
rect 6520 1732 6522 1736
rect 6514 1730 6522 1732
rect 6538 1736 6546 1738
rect 6538 1732 6540 1736
rect 6544 1732 6546 1736
rect 6538 1730 6546 1732
rect 6562 1736 6570 1738
rect 6562 1732 6564 1736
rect 6568 1732 6570 1736
rect 6562 1730 6570 1732
rect 6586 1736 6594 1738
rect 6586 1732 6588 1736
rect 6592 1732 6594 1736
rect 6586 1730 6594 1732
rect 6610 1736 6618 1738
rect 6610 1732 6612 1736
rect 6616 1732 6618 1736
rect 6610 1730 6618 1732
rect 6634 1736 6642 1738
rect 6634 1732 6636 1736
rect 6640 1732 6642 1736
rect 6634 1730 6642 1732
rect 6658 1736 6666 1738
rect 6658 1732 6660 1736
rect 6664 1732 6666 1736
rect 6658 1730 6666 1732
rect 6682 1736 6690 1738
rect 6682 1732 6684 1736
rect 6688 1732 6690 1736
rect 6682 1730 6690 1732
rect 6898 1736 6906 1738
rect 6898 1732 6900 1736
rect 6904 1732 6906 1736
rect 6898 1730 6906 1732
rect 6922 1736 6930 1738
rect 6922 1732 6924 1736
rect 6928 1732 6930 1736
rect 6922 1730 6930 1732
rect 6946 1736 6954 1738
rect 6946 1732 6948 1736
rect 6952 1732 6954 1736
rect 6946 1730 6954 1732
rect 6970 1736 6978 1738
rect 6970 1732 6972 1736
rect 6976 1732 6978 1736
rect 6970 1730 6978 1732
rect 6994 1736 7002 1738
rect 6994 1732 6996 1736
rect 7000 1732 7002 1736
rect 6994 1730 7002 1732
rect 7018 1736 7026 1738
rect 7018 1732 7020 1736
rect 7024 1732 7026 1736
rect 7018 1730 7026 1732
rect 7042 1736 7050 1738
rect 7042 1732 7044 1736
rect 7048 1732 7050 1736
rect 7042 1730 7050 1732
rect 7066 1736 7074 1738
rect 7066 1732 7068 1736
rect 7072 1732 7074 1736
rect 7066 1730 7074 1732
rect 7090 1736 7098 1738
rect 7090 1732 7092 1736
rect 7096 1732 7098 1736
rect 7090 1730 7098 1732
rect 7114 1736 7122 1738
rect 7114 1732 7116 1736
rect 7120 1732 7122 1736
rect 7114 1730 7122 1732
rect 7138 1736 7146 1738
rect 7138 1732 7140 1736
rect 7144 1732 7146 1736
rect 7138 1730 7146 1732
rect 7162 1736 7170 1738
rect 7162 1732 7164 1736
rect 7168 1732 7170 1736
rect 7162 1730 7170 1732
rect 7186 1736 7194 1738
rect 7186 1732 7188 1736
rect 7192 1732 7194 1736
rect 7186 1730 7194 1732
rect 2400 1724 2406 1726
rect 2404 1720 2406 1724
rect 2400 1718 2406 1720
rect 2422 1724 2430 1726
rect 2422 1720 2424 1724
rect 2428 1720 2430 1724
rect 2422 1718 2430 1720
rect 2446 1724 2454 1726
rect 2446 1720 2448 1724
rect 2452 1720 2454 1724
rect 2446 1718 2454 1720
rect 2470 1724 2478 1726
rect 2470 1720 2472 1724
rect 2476 1720 2478 1724
rect 2470 1718 2478 1720
rect 2494 1724 2502 1726
rect 2494 1720 2496 1724
rect 2500 1720 2502 1724
rect 2494 1718 2502 1720
rect 2710 1724 2718 1726
rect 2710 1720 2712 1724
rect 2716 1720 2718 1724
rect 2710 1718 2718 1720
rect 2734 1724 2742 1726
rect 2734 1720 2736 1724
rect 2740 1720 2742 1724
rect 2734 1718 2742 1720
rect 2758 1724 2766 1726
rect 2758 1720 2760 1724
rect 2764 1720 2766 1724
rect 2758 1718 2766 1720
rect 2782 1724 2790 1726
rect 2782 1720 2784 1724
rect 2788 1720 2790 1724
rect 2782 1718 2790 1720
rect 2806 1724 2814 1726
rect 2806 1720 2808 1724
rect 2812 1720 2814 1724
rect 2806 1718 2814 1720
rect 2830 1724 2838 1726
rect 2830 1720 2832 1724
rect 2836 1720 2838 1724
rect 2830 1718 2838 1720
rect 2854 1724 2862 1726
rect 2854 1720 2856 1724
rect 2860 1720 2862 1724
rect 2854 1718 2862 1720
rect 2878 1724 2886 1726
rect 2878 1720 2880 1724
rect 2884 1720 2886 1724
rect 2878 1718 2886 1720
rect 2902 1724 2910 1726
rect 2902 1720 2904 1724
rect 2908 1720 2910 1724
rect 2902 1718 2910 1720
rect 2926 1724 2934 1726
rect 2926 1720 2928 1724
rect 2932 1720 2934 1724
rect 2926 1718 2934 1720
rect 2950 1724 2958 1726
rect 2950 1720 2952 1724
rect 2956 1720 2958 1724
rect 2950 1718 2958 1720
rect 2974 1724 2982 1726
rect 2974 1720 2976 1724
rect 2980 1720 2982 1724
rect 2974 1718 2982 1720
rect 2998 1724 3006 1726
rect 2998 1720 3000 1724
rect 3004 1720 3006 1724
rect 2998 1718 3006 1720
rect 3022 1724 3030 1726
rect 3022 1720 3024 1724
rect 3028 1720 3030 1724
rect 3022 1718 3030 1720
rect 3046 1724 3054 1726
rect 3046 1720 3048 1724
rect 3052 1720 3054 1724
rect 3046 1718 3054 1720
rect 3070 1724 3078 1726
rect 3070 1720 3072 1724
rect 3076 1720 3078 1724
rect 3070 1718 3078 1720
rect 3094 1724 3102 1726
rect 3094 1720 3096 1724
rect 3100 1720 3102 1724
rect 3094 1718 3102 1720
rect 3310 1724 3318 1726
rect 3310 1720 3312 1724
rect 3316 1720 3318 1724
rect 3310 1718 3318 1720
rect 3334 1724 3342 1726
rect 3334 1720 3336 1724
rect 3340 1720 3342 1724
rect 3334 1718 3342 1720
rect 3358 1724 3366 1726
rect 3358 1720 3360 1724
rect 3364 1720 3366 1724
rect 3358 1718 3366 1720
rect 3382 1724 3390 1726
rect 3382 1720 3384 1724
rect 3388 1720 3390 1724
rect 3382 1718 3390 1720
rect 3406 1724 3414 1726
rect 3406 1720 3408 1724
rect 3412 1720 3414 1724
rect 3406 1718 3414 1720
rect 3430 1724 3438 1726
rect 3430 1720 3432 1724
rect 3436 1720 3438 1724
rect 3430 1718 3438 1720
rect 3454 1724 3462 1726
rect 3454 1720 3456 1724
rect 3460 1720 3462 1724
rect 3454 1718 3462 1720
rect 3478 1724 3486 1726
rect 3478 1720 3480 1724
rect 3484 1720 3486 1724
rect 3478 1718 3486 1720
rect 3502 1724 3510 1726
rect 3502 1720 3504 1724
rect 3508 1720 3510 1724
rect 3502 1718 3510 1720
rect 3526 1724 3534 1726
rect 3526 1720 3528 1724
rect 3532 1720 3534 1724
rect 3526 1718 3534 1720
rect 3550 1724 3558 1726
rect 3550 1720 3552 1724
rect 3556 1720 3558 1724
rect 3550 1718 3558 1720
rect 3574 1724 3582 1726
rect 3574 1720 3576 1724
rect 3580 1720 3582 1724
rect 3574 1718 3582 1720
rect 3598 1724 3606 1726
rect 3598 1720 3600 1724
rect 3604 1720 3606 1724
rect 3598 1718 3606 1720
rect 3622 1724 3630 1726
rect 3622 1720 3624 1724
rect 3628 1720 3630 1724
rect 3622 1718 3630 1720
rect 3646 1724 3654 1726
rect 3646 1720 3648 1724
rect 3652 1720 3654 1724
rect 3646 1718 3654 1720
rect 3670 1724 3678 1726
rect 3670 1720 3672 1724
rect 3676 1720 3678 1724
rect 3670 1718 3678 1720
rect 3694 1724 3702 1726
rect 3694 1720 3696 1724
rect 3700 1720 3702 1724
rect 3694 1718 3702 1720
rect 3910 1724 3918 1726
rect 3910 1720 3912 1724
rect 3916 1720 3918 1724
rect 3910 1718 3918 1720
rect 3934 1724 3942 1726
rect 3934 1720 3936 1724
rect 3940 1720 3942 1724
rect 3934 1718 3942 1720
rect 3958 1724 3966 1726
rect 3958 1720 3960 1724
rect 3964 1720 3966 1724
rect 3958 1718 3966 1720
rect 3982 1724 3990 1726
rect 3982 1720 3984 1724
rect 3988 1720 3990 1724
rect 3982 1718 3990 1720
rect 4006 1724 4014 1726
rect 4006 1720 4008 1724
rect 4012 1720 4014 1724
rect 4006 1718 4014 1720
rect 4030 1724 4038 1726
rect 4030 1720 4032 1724
rect 4036 1720 4038 1724
rect 4030 1718 4038 1720
rect 4054 1724 4062 1726
rect 4054 1720 4056 1724
rect 4060 1720 4062 1724
rect 4054 1718 4062 1720
rect 4078 1724 4086 1726
rect 4078 1720 4080 1724
rect 4084 1720 4086 1724
rect 4078 1718 4086 1720
rect 4102 1724 4110 1726
rect 4102 1720 4104 1724
rect 4108 1720 4110 1724
rect 4102 1718 4110 1720
rect 4126 1724 4134 1726
rect 4126 1720 4128 1724
rect 4132 1720 4134 1724
rect 4126 1718 4134 1720
rect 4150 1724 4158 1726
rect 4150 1720 4152 1724
rect 4156 1720 4158 1724
rect 4150 1718 4158 1720
rect 4174 1724 4182 1726
rect 4174 1720 4176 1724
rect 4180 1720 4182 1724
rect 4174 1718 4182 1720
rect 4198 1724 4206 1726
rect 4198 1720 4200 1724
rect 4204 1720 4206 1724
rect 4198 1718 4206 1720
rect 4222 1724 4230 1726
rect 4222 1720 4224 1724
rect 4228 1720 4230 1724
rect 4222 1718 4230 1720
rect 4246 1724 4254 1726
rect 4246 1720 4248 1724
rect 4252 1720 4254 1724
rect 4246 1718 4254 1720
rect 4270 1724 4278 1726
rect 4270 1720 4272 1724
rect 4276 1720 4278 1724
rect 4270 1718 4278 1720
rect 4294 1724 4302 1726
rect 4294 1720 4296 1724
rect 4300 1720 4302 1724
rect 4294 1718 4302 1720
rect 4510 1724 4518 1726
rect 4510 1720 4512 1724
rect 4516 1720 4518 1724
rect 4510 1718 4518 1720
rect 4534 1724 4542 1726
rect 4534 1720 4536 1724
rect 4540 1720 4542 1724
rect 4534 1718 4542 1720
rect 4558 1724 4566 1726
rect 4558 1720 4560 1724
rect 4564 1720 4566 1724
rect 4558 1718 4566 1720
rect 4582 1724 4590 1726
rect 4582 1720 4584 1724
rect 4588 1720 4590 1724
rect 4582 1718 4590 1720
rect 4606 1724 4614 1726
rect 4606 1720 4608 1724
rect 4612 1720 4614 1724
rect 4606 1718 4614 1720
rect 4630 1724 4638 1726
rect 4630 1720 4632 1724
rect 4636 1720 4638 1724
rect 4630 1718 4638 1720
rect 4654 1724 4662 1726
rect 4654 1720 4656 1724
rect 4660 1720 4662 1724
rect 4654 1718 4662 1720
rect 4678 1724 4686 1726
rect 4678 1720 4680 1724
rect 4684 1720 4686 1724
rect 4678 1718 4686 1720
rect 4702 1724 4710 1726
rect 4702 1720 4704 1724
rect 4708 1720 4710 1724
rect 4702 1718 4710 1720
rect 4726 1724 4734 1726
rect 4726 1720 4728 1724
rect 4732 1720 4734 1724
rect 4726 1718 4734 1720
rect 4750 1724 4758 1726
rect 4750 1720 4752 1724
rect 4756 1720 4758 1724
rect 4750 1718 4758 1720
rect 4774 1724 4782 1726
rect 4774 1720 4776 1724
rect 4780 1720 4782 1724
rect 4774 1718 4782 1720
rect 4798 1718 4800 1726
rect 5710 1724 5718 1726
rect 5710 1720 5712 1724
rect 5716 1720 5718 1724
rect 5710 1718 5718 1720
rect 5734 1724 5742 1726
rect 5734 1720 5736 1724
rect 5740 1720 5742 1724
rect 5734 1718 5742 1720
rect 5758 1724 5766 1726
rect 5758 1720 5760 1724
rect 5764 1720 5766 1724
rect 5758 1718 5766 1720
rect 5782 1724 5790 1726
rect 5782 1720 5784 1724
rect 5788 1720 5790 1724
rect 5782 1718 5790 1720
rect 5806 1724 5814 1726
rect 5806 1720 5808 1724
rect 5812 1720 5814 1724
rect 5806 1718 5814 1720
rect 5830 1724 5838 1726
rect 5830 1720 5832 1724
rect 5836 1720 5838 1724
rect 5830 1718 5838 1720
rect 5854 1724 5862 1726
rect 5854 1720 5856 1724
rect 5860 1720 5862 1724
rect 5854 1718 5862 1720
rect 5878 1724 5886 1726
rect 5878 1720 5880 1724
rect 5884 1720 5886 1724
rect 5878 1718 5886 1720
rect 5902 1724 5910 1726
rect 5902 1720 5904 1724
rect 5908 1720 5910 1724
rect 5902 1718 5910 1720
rect 5926 1724 5934 1726
rect 5926 1720 5928 1724
rect 5932 1720 5934 1724
rect 5926 1718 5934 1720
rect 5950 1724 5958 1726
rect 5950 1720 5952 1724
rect 5956 1720 5958 1724
rect 5950 1718 5958 1720
rect 5974 1724 5982 1726
rect 5974 1720 5976 1724
rect 5980 1720 5982 1724
rect 5974 1718 5982 1720
rect 5998 1724 6006 1726
rect 5998 1720 6000 1724
rect 6004 1720 6006 1724
rect 5998 1718 6006 1720
rect 6022 1724 6030 1726
rect 6022 1720 6024 1724
rect 6028 1720 6030 1724
rect 6022 1718 6030 1720
rect 6046 1724 6054 1726
rect 6046 1720 6048 1724
rect 6052 1720 6054 1724
rect 6046 1718 6054 1720
rect 6070 1724 6078 1726
rect 6070 1720 6072 1724
rect 6076 1720 6078 1724
rect 6070 1718 6078 1720
rect 6094 1724 6102 1726
rect 6094 1720 6096 1724
rect 6100 1720 6102 1724
rect 6094 1718 6102 1720
rect 6310 1724 6318 1726
rect 6310 1720 6312 1724
rect 6316 1720 6318 1724
rect 6310 1718 6318 1720
rect 6334 1724 6342 1726
rect 6334 1720 6336 1724
rect 6340 1720 6342 1724
rect 6334 1718 6342 1720
rect 6358 1724 6366 1726
rect 6358 1720 6360 1724
rect 6364 1720 6366 1724
rect 6358 1718 6366 1720
rect 6382 1724 6390 1726
rect 6382 1720 6384 1724
rect 6388 1720 6390 1724
rect 6382 1718 6390 1720
rect 6406 1724 6414 1726
rect 6406 1720 6408 1724
rect 6412 1720 6414 1724
rect 6406 1718 6414 1720
rect 6430 1724 6438 1726
rect 6430 1720 6432 1724
rect 6436 1720 6438 1724
rect 6430 1718 6438 1720
rect 6454 1724 6462 1726
rect 6454 1720 6456 1724
rect 6460 1720 6462 1724
rect 6454 1718 6462 1720
rect 6478 1724 6486 1726
rect 6478 1720 6480 1724
rect 6484 1720 6486 1724
rect 6478 1718 6486 1720
rect 6502 1724 6510 1726
rect 6502 1720 6504 1724
rect 6508 1720 6510 1724
rect 6502 1718 6510 1720
rect 6526 1724 6534 1726
rect 6526 1720 6528 1724
rect 6532 1720 6534 1724
rect 6526 1718 6534 1720
rect 6550 1724 6558 1726
rect 6550 1720 6552 1724
rect 6556 1720 6558 1724
rect 6550 1718 6558 1720
rect 6574 1724 6582 1726
rect 6574 1720 6576 1724
rect 6580 1720 6582 1724
rect 6574 1718 6582 1720
rect 6598 1724 6606 1726
rect 6598 1720 6600 1724
rect 6604 1720 6606 1724
rect 6598 1718 6606 1720
rect 6622 1724 6630 1726
rect 6622 1720 6624 1724
rect 6628 1720 6630 1724
rect 6622 1718 6630 1720
rect 6646 1724 6654 1726
rect 6646 1720 6648 1724
rect 6652 1720 6654 1724
rect 6646 1718 6654 1720
rect 6670 1724 6678 1726
rect 6670 1720 6672 1724
rect 6676 1720 6678 1724
rect 6670 1718 6678 1720
rect 6694 1724 6702 1726
rect 6694 1720 6696 1724
rect 6700 1720 6702 1724
rect 6694 1718 6702 1720
rect 6910 1724 6918 1726
rect 6910 1720 6912 1724
rect 6916 1720 6918 1724
rect 6910 1718 6918 1720
rect 6934 1724 6942 1726
rect 6934 1720 6936 1724
rect 6940 1720 6942 1724
rect 6934 1718 6942 1720
rect 6958 1724 6966 1726
rect 6958 1720 6960 1724
rect 6964 1720 6966 1724
rect 6958 1718 6966 1720
rect 6982 1724 6990 1726
rect 6982 1720 6984 1724
rect 6988 1720 6990 1724
rect 6982 1718 6990 1720
rect 7006 1724 7014 1726
rect 7006 1720 7008 1724
rect 7012 1720 7014 1724
rect 7006 1718 7014 1720
rect 7030 1724 7038 1726
rect 7030 1720 7032 1724
rect 7036 1720 7038 1724
rect 7030 1718 7038 1720
rect 7054 1724 7062 1726
rect 7054 1720 7056 1724
rect 7060 1720 7062 1724
rect 7054 1718 7062 1720
rect 7078 1724 7086 1726
rect 7078 1720 7080 1724
rect 7084 1720 7086 1724
rect 7078 1718 7086 1720
rect 7102 1724 7110 1726
rect 7102 1720 7104 1724
rect 7108 1720 7110 1724
rect 7102 1718 7110 1720
rect 7126 1724 7134 1726
rect 7126 1720 7128 1724
rect 7132 1720 7134 1724
rect 7126 1718 7134 1720
rect 7150 1724 7158 1726
rect 7150 1720 7152 1724
rect 7156 1720 7158 1724
rect 7150 1718 7158 1720
rect 7174 1724 7182 1726
rect 7174 1720 7176 1724
rect 7180 1720 7182 1724
rect 7174 1718 7182 1720
rect 7198 1718 7200 1726
rect 2410 1712 2418 1714
rect 2410 1708 2412 1712
rect 2416 1708 2418 1712
rect 2410 1706 2418 1708
rect 2434 1712 2442 1714
rect 2434 1708 2436 1712
rect 2440 1708 2442 1712
rect 2434 1706 2442 1708
rect 2458 1712 2466 1714
rect 2458 1708 2460 1712
rect 2464 1708 2466 1712
rect 2458 1706 2466 1708
rect 2482 1712 2490 1714
rect 2482 1708 2484 1712
rect 2488 1708 2490 1712
rect 2482 1706 2490 1708
rect 2698 1712 2706 1714
rect 2698 1708 2700 1712
rect 2704 1708 2706 1712
rect 2698 1706 2706 1708
rect 2722 1712 2730 1714
rect 2722 1708 2724 1712
rect 2728 1708 2730 1712
rect 2722 1706 2730 1708
rect 2746 1712 2754 1714
rect 2746 1708 2748 1712
rect 2752 1708 2754 1712
rect 2746 1706 2754 1708
rect 2770 1712 2778 1714
rect 2770 1708 2772 1712
rect 2776 1708 2778 1712
rect 2770 1706 2778 1708
rect 2794 1712 2802 1714
rect 2794 1708 2796 1712
rect 2800 1708 2802 1712
rect 2794 1706 2802 1708
rect 2818 1712 2826 1714
rect 2818 1708 2820 1712
rect 2824 1708 2826 1712
rect 2818 1706 2826 1708
rect 2842 1712 2850 1714
rect 2842 1708 2844 1712
rect 2848 1708 2850 1712
rect 2842 1706 2850 1708
rect 2866 1712 2874 1714
rect 2866 1708 2868 1712
rect 2872 1708 2874 1712
rect 2866 1706 2874 1708
rect 2890 1712 2898 1714
rect 2890 1708 2892 1712
rect 2896 1708 2898 1712
rect 2890 1706 2898 1708
rect 2914 1712 2922 1714
rect 2914 1708 2916 1712
rect 2920 1708 2922 1712
rect 2914 1706 2922 1708
rect 2938 1712 2946 1714
rect 2938 1708 2940 1712
rect 2944 1708 2946 1712
rect 2938 1706 2946 1708
rect 2962 1712 2970 1714
rect 2962 1708 2964 1712
rect 2968 1708 2970 1712
rect 2962 1706 2970 1708
rect 2986 1712 2994 1714
rect 2986 1708 2988 1712
rect 2992 1708 2994 1712
rect 2986 1706 2994 1708
rect 3010 1712 3018 1714
rect 3010 1708 3012 1712
rect 3016 1708 3018 1712
rect 3010 1706 3018 1708
rect 3034 1712 3042 1714
rect 3034 1708 3036 1712
rect 3040 1708 3042 1712
rect 3034 1706 3042 1708
rect 3058 1712 3066 1714
rect 3058 1708 3060 1712
rect 3064 1708 3066 1712
rect 3058 1706 3066 1708
rect 3082 1712 3090 1714
rect 3082 1708 3084 1712
rect 3088 1708 3090 1712
rect 3082 1706 3090 1708
rect 3298 1712 3306 1714
rect 3298 1708 3300 1712
rect 3304 1708 3306 1712
rect 3298 1706 3306 1708
rect 3322 1712 3330 1714
rect 3322 1708 3324 1712
rect 3328 1708 3330 1712
rect 3322 1706 3330 1708
rect 3346 1712 3354 1714
rect 3346 1708 3348 1712
rect 3352 1708 3354 1712
rect 3346 1706 3354 1708
rect 3370 1712 3378 1714
rect 3370 1708 3372 1712
rect 3376 1708 3378 1712
rect 3370 1706 3378 1708
rect 3394 1712 3402 1714
rect 3394 1708 3396 1712
rect 3400 1708 3402 1712
rect 3394 1706 3402 1708
rect 3418 1712 3426 1714
rect 3418 1708 3420 1712
rect 3424 1708 3426 1712
rect 3418 1706 3426 1708
rect 3442 1712 3450 1714
rect 3442 1708 3444 1712
rect 3448 1708 3450 1712
rect 3442 1706 3450 1708
rect 3466 1712 3474 1714
rect 3466 1708 3468 1712
rect 3472 1708 3474 1712
rect 3466 1706 3474 1708
rect 3490 1712 3498 1714
rect 3490 1708 3492 1712
rect 3496 1708 3498 1712
rect 3490 1706 3498 1708
rect 3514 1712 3522 1714
rect 3514 1708 3516 1712
rect 3520 1708 3522 1712
rect 3514 1706 3522 1708
rect 3538 1712 3546 1714
rect 3538 1708 3540 1712
rect 3544 1708 3546 1712
rect 3538 1706 3546 1708
rect 3562 1712 3570 1714
rect 3562 1708 3564 1712
rect 3568 1708 3570 1712
rect 3562 1706 3570 1708
rect 3586 1712 3594 1714
rect 3586 1708 3588 1712
rect 3592 1708 3594 1712
rect 3586 1706 3594 1708
rect 3610 1712 3618 1714
rect 3610 1708 3612 1712
rect 3616 1708 3618 1712
rect 3610 1706 3618 1708
rect 3634 1712 3642 1714
rect 3634 1708 3636 1712
rect 3640 1708 3642 1712
rect 3634 1706 3642 1708
rect 3658 1712 3666 1714
rect 3658 1708 3660 1712
rect 3664 1708 3666 1712
rect 3658 1706 3666 1708
rect 3682 1712 3690 1714
rect 3682 1708 3684 1712
rect 3688 1708 3690 1712
rect 3682 1706 3690 1708
rect 3898 1712 3906 1714
rect 3898 1708 3900 1712
rect 3904 1708 3906 1712
rect 3898 1706 3906 1708
rect 3922 1712 3930 1714
rect 3922 1708 3924 1712
rect 3928 1708 3930 1712
rect 3922 1706 3930 1708
rect 3946 1712 3954 1714
rect 3946 1708 3948 1712
rect 3952 1708 3954 1712
rect 3946 1706 3954 1708
rect 3970 1712 3978 1714
rect 3970 1708 3972 1712
rect 3976 1708 3978 1712
rect 3970 1706 3978 1708
rect 3994 1712 4002 1714
rect 3994 1708 3996 1712
rect 4000 1708 4002 1712
rect 3994 1706 4002 1708
rect 4018 1712 4026 1714
rect 4018 1708 4020 1712
rect 4024 1708 4026 1712
rect 4018 1706 4026 1708
rect 4042 1712 4050 1714
rect 4042 1708 4044 1712
rect 4048 1708 4050 1712
rect 4042 1706 4050 1708
rect 4066 1712 4074 1714
rect 4066 1708 4068 1712
rect 4072 1708 4074 1712
rect 4066 1706 4074 1708
rect 4090 1712 4098 1714
rect 4090 1708 4092 1712
rect 4096 1708 4098 1712
rect 4090 1706 4098 1708
rect 4114 1712 4122 1714
rect 4114 1708 4116 1712
rect 4120 1708 4122 1712
rect 4114 1706 4122 1708
rect 4138 1712 4146 1714
rect 4138 1708 4140 1712
rect 4144 1708 4146 1712
rect 4138 1706 4146 1708
rect 4162 1712 4170 1714
rect 4162 1708 4164 1712
rect 4168 1708 4170 1712
rect 4162 1706 4170 1708
rect 4186 1712 4194 1714
rect 4186 1708 4188 1712
rect 4192 1708 4194 1712
rect 4186 1706 4194 1708
rect 4210 1712 4218 1714
rect 4210 1708 4212 1712
rect 4216 1708 4218 1712
rect 4210 1706 4218 1708
rect 4234 1712 4242 1714
rect 4234 1708 4236 1712
rect 4240 1708 4242 1712
rect 4234 1706 4242 1708
rect 4258 1712 4266 1714
rect 4258 1708 4260 1712
rect 4264 1708 4266 1712
rect 4258 1706 4266 1708
rect 4282 1712 4290 1714
rect 4282 1708 4284 1712
rect 4288 1708 4290 1712
rect 4282 1706 4290 1708
rect 4498 1712 4506 1714
rect 4498 1708 4500 1712
rect 4504 1708 4506 1712
rect 4498 1706 4506 1708
rect 4522 1712 4530 1714
rect 4522 1708 4524 1712
rect 4528 1708 4530 1712
rect 4522 1706 4530 1708
rect 4546 1712 4554 1714
rect 4546 1708 4548 1712
rect 4552 1708 4554 1712
rect 4546 1706 4554 1708
rect 4570 1712 4578 1714
rect 4570 1708 4572 1712
rect 4576 1708 4578 1712
rect 4570 1706 4578 1708
rect 4594 1712 4602 1714
rect 4594 1708 4596 1712
rect 4600 1708 4602 1712
rect 4594 1706 4602 1708
rect 4618 1712 4626 1714
rect 4618 1708 4620 1712
rect 4624 1708 4626 1712
rect 4618 1706 4626 1708
rect 4642 1712 4650 1714
rect 4642 1708 4644 1712
rect 4648 1708 4650 1712
rect 4642 1706 4650 1708
rect 4666 1712 4674 1714
rect 4666 1708 4668 1712
rect 4672 1708 4674 1712
rect 4666 1706 4674 1708
rect 4690 1712 4698 1714
rect 4690 1708 4692 1712
rect 4696 1708 4698 1712
rect 4690 1706 4698 1708
rect 4714 1712 4722 1714
rect 4714 1708 4716 1712
rect 4720 1708 4722 1712
rect 4714 1706 4722 1708
rect 4738 1712 4746 1714
rect 4738 1708 4740 1712
rect 4744 1708 4746 1712
rect 4738 1706 4746 1708
rect 4762 1712 4770 1714
rect 4762 1708 4764 1712
rect 4768 1708 4770 1712
rect 4762 1706 4770 1708
rect 4786 1712 4794 1714
rect 4786 1708 4788 1712
rect 4792 1708 4794 1712
rect 4786 1706 4794 1708
rect 5698 1712 5706 1714
rect 5698 1708 5700 1712
rect 5704 1708 5706 1712
rect 5698 1706 5706 1708
rect 5722 1712 5730 1714
rect 5722 1708 5724 1712
rect 5728 1708 5730 1712
rect 5722 1706 5730 1708
rect 5746 1712 5754 1714
rect 5746 1708 5748 1712
rect 5752 1708 5754 1712
rect 5746 1706 5754 1708
rect 5770 1712 5778 1714
rect 5770 1708 5772 1712
rect 5776 1708 5778 1712
rect 5770 1706 5778 1708
rect 5794 1712 5802 1714
rect 5794 1708 5796 1712
rect 5800 1708 5802 1712
rect 5794 1706 5802 1708
rect 5818 1712 5826 1714
rect 5818 1708 5820 1712
rect 5824 1708 5826 1712
rect 5818 1706 5826 1708
rect 5842 1712 5850 1714
rect 5842 1708 5844 1712
rect 5848 1708 5850 1712
rect 5842 1706 5850 1708
rect 5866 1712 5874 1714
rect 5866 1708 5868 1712
rect 5872 1708 5874 1712
rect 5866 1706 5874 1708
rect 5890 1712 5898 1714
rect 5890 1708 5892 1712
rect 5896 1708 5898 1712
rect 5890 1706 5898 1708
rect 5914 1712 5922 1714
rect 5914 1708 5916 1712
rect 5920 1708 5922 1712
rect 5914 1706 5922 1708
rect 5938 1712 5946 1714
rect 5938 1708 5940 1712
rect 5944 1708 5946 1712
rect 5938 1706 5946 1708
rect 5962 1712 5970 1714
rect 5962 1708 5964 1712
rect 5968 1708 5970 1712
rect 5962 1706 5970 1708
rect 5986 1712 5994 1714
rect 5986 1708 5988 1712
rect 5992 1708 5994 1712
rect 5986 1706 5994 1708
rect 6010 1712 6018 1714
rect 6010 1708 6012 1712
rect 6016 1708 6018 1712
rect 6010 1706 6018 1708
rect 6034 1712 6042 1714
rect 6034 1708 6036 1712
rect 6040 1708 6042 1712
rect 6034 1706 6042 1708
rect 6058 1712 6066 1714
rect 6058 1708 6060 1712
rect 6064 1708 6066 1712
rect 6058 1706 6066 1708
rect 6082 1712 6090 1714
rect 6082 1708 6084 1712
rect 6088 1708 6090 1712
rect 6082 1706 6090 1708
rect 6298 1712 6306 1714
rect 6298 1708 6300 1712
rect 6304 1708 6306 1712
rect 6298 1706 6306 1708
rect 6322 1712 6330 1714
rect 6322 1708 6324 1712
rect 6328 1708 6330 1712
rect 6322 1706 6330 1708
rect 6346 1712 6354 1714
rect 6346 1708 6348 1712
rect 6352 1708 6354 1712
rect 6346 1706 6354 1708
rect 6370 1712 6378 1714
rect 6370 1708 6372 1712
rect 6376 1708 6378 1712
rect 6370 1706 6378 1708
rect 6394 1712 6402 1714
rect 6394 1708 6396 1712
rect 6400 1708 6402 1712
rect 6394 1706 6402 1708
rect 6418 1712 6426 1714
rect 6418 1708 6420 1712
rect 6424 1708 6426 1712
rect 6418 1706 6426 1708
rect 6442 1712 6450 1714
rect 6442 1708 6444 1712
rect 6448 1708 6450 1712
rect 6442 1706 6450 1708
rect 6466 1712 6474 1714
rect 6466 1708 6468 1712
rect 6472 1708 6474 1712
rect 6466 1706 6474 1708
rect 6490 1712 6498 1714
rect 6490 1708 6492 1712
rect 6496 1708 6498 1712
rect 6490 1706 6498 1708
rect 6514 1712 6522 1714
rect 6514 1708 6516 1712
rect 6520 1708 6522 1712
rect 6514 1706 6522 1708
rect 6538 1712 6546 1714
rect 6538 1708 6540 1712
rect 6544 1708 6546 1712
rect 6538 1706 6546 1708
rect 6562 1712 6570 1714
rect 6562 1708 6564 1712
rect 6568 1708 6570 1712
rect 6562 1706 6570 1708
rect 6586 1712 6594 1714
rect 6586 1708 6588 1712
rect 6592 1708 6594 1712
rect 6586 1706 6594 1708
rect 6610 1712 6618 1714
rect 6610 1708 6612 1712
rect 6616 1708 6618 1712
rect 6610 1706 6618 1708
rect 6634 1712 6642 1714
rect 6634 1708 6636 1712
rect 6640 1708 6642 1712
rect 6634 1706 6642 1708
rect 6658 1712 6666 1714
rect 6658 1708 6660 1712
rect 6664 1708 6666 1712
rect 6658 1706 6666 1708
rect 6682 1712 6690 1714
rect 6682 1708 6684 1712
rect 6688 1708 6690 1712
rect 6682 1706 6690 1708
rect 6898 1712 6906 1714
rect 6898 1708 6900 1712
rect 6904 1708 6906 1712
rect 6898 1706 6906 1708
rect 6922 1712 6930 1714
rect 6922 1708 6924 1712
rect 6928 1708 6930 1712
rect 6922 1706 6930 1708
rect 6946 1712 6954 1714
rect 6946 1708 6948 1712
rect 6952 1708 6954 1712
rect 6946 1706 6954 1708
rect 6970 1712 6978 1714
rect 6970 1708 6972 1712
rect 6976 1708 6978 1712
rect 6970 1706 6978 1708
rect 6994 1712 7002 1714
rect 6994 1708 6996 1712
rect 7000 1708 7002 1712
rect 6994 1706 7002 1708
rect 7018 1712 7026 1714
rect 7018 1708 7020 1712
rect 7024 1708 7026 1712
rect 7018 1706 7026 1708
rect 7042 1712 7050 1714
rect 7042 1708 7044 1712
rect 7048 1708 7050 1712
rect 7042 1706 7050 1708
rect 7066 1712 7074 1714
rect 7066 1708 7068 1712
rect 7072 1708 7074 1712
rect 7066 1706 7074 1708
rect 7090 1712 7098 1714
rect 7090 1708 7092 1712
rect 7096 1708 7098 1712
rect 7090 1706 7098 1708
rect 7114 1712 7122 1714
rect 7114 1708 7116 1712
rect 7120 1708 7122 1712
rect 7114 1706 7122 1708
rect 7138 1712 7146 1714
rect 7138 1708 7140 1712
rect 7144 1708 7146 1712
rect 7138 1706 7146 1708
rect 7162 1712 7170 1714
rect 7162 1708 7164 1712
rect 7168 1708 7170 1712
rect 7162 1706 7170 1708
rect 7186 1712 7194 1714
rect 7186 1708 7188 1712
rect 7192 1708 7194 1712
rect 7186 1706 7194 1708
rect 2400 1700 2406 1702
rect 2404 1696 2406 1700
rect 2400 1694 2406 1696
rect 2422 1700 2430 1702
rect 2422 1696 2424 1700
rect 2428 1696 2430 1700
rect 2422 1694 2430 1696
rect 2446 1700 2454 1702
rect 2446 1696 2448 1700
rect 2452 1696 2454 1700
rect 2446 1694 2454 1696
rect 2470 1700 2478 1702
rect 2470 1696 2472 1700
rect 2476 1696 2478 1700
rect 2470 1694 2478 1696
rect 2494 1700 2502 1702
rect 2494 1696 2496 1700
rect 2500 1696 2502 1700
rect 2494 1694 2502 1696
rect 2710 1700 2718 1702
rect 2710 1696 2712 1700
rect 2716 1696 2718 1700
rect 2710 1694 2718 1696
rect 2734 1700 2742 1702
rect 2734 1696 2736 1700
rect 2740 1696 2742 1700
rect 2734 1694 2742 1696
rect 2758 1700 2766 1702
rect 2758 1696 2760 1700
rect 2764 1696 2766 1700
rect 2758 1694 2766 1696
rect 2782 1700 2790 1702
rect 2782 1696 2784 1700
rect 2788 1696 2790 1700
rect 2782 1694 2790 1696
rect 2806 1700 2814 1702
rect 2806 1696 2808 1700
rect 2812 1696 2814 1700
rect 2806 1694 2814 1696
rect 2830 1700 2838 1702
rect 2830 1696 2832 1700
rect 2836 1696 2838 1700
rect 2830 1694 2838 1696
rect 2854 1700 2862 1702
rect 2854 1696 2856 1700
rect 2860 1696 2862 1700
rect 2854 1694 2862 1696
rect 2878 1700 2886 1702
rect 2878 1696 2880 1700
rect 2884 1696 2886 1700
rect 2878 1694 2886 1696
rect 2902 1700 2910 1702
rect 2902 1696 2904 1700
rect 2908 1696 2910 1700
rect 2902 1694 2910 1696
rect 2926 1700 2934 1702
rect 2926 1696 2928 1700
rect 2932 1696 2934 1700
rect 2926 1694 2934 1696
rect 2950 1700 2958 1702
rect 2950 1696 2952 1700
rect 2956 1696 2958 1700
rect 2950 1694 2958 1696
rect 2974 1700 2982 1702
rect 2974 1696 2976 1700
rect 2980 1696 2982 1700
rect 2974 1694 2982 1696
rect 2998 1700 3006 1702
rect 2998 1696 3000 1700
rect 3004 1696 3006 1700
rect 2998 1694 3006 1696
rect 3022 1700 3030 1702
rect 3022 1696 3024 1700
rect 3028 1696 3030 1700
rect 3022 1694 3030 1696
rect 3046 1700 3054 1702
rect 3046 1696 3048 1700
rect 3052 1696 3054 1700
rect 3046 1694 3054 1696
rect 3070 1700 3078 1702
rect 3070 1696 3072 1700
rect 3076 1696 3078 1700
rect 3070 1694 3078 1696
rect 3094 1700 3102 1702
rect 3094 1696 3096 1700
rect 3100 1696 3102 1700
rect 3094 1694 3102 1696
rect 3310 1700 3318 1702
rect 3310 1696 3312 1700
rect 3316 1696 3318 1700
rect 3310 1694 3318 1696
rect 3334 1700 3342 1702
rect 3334 1696 3336 1700
rect 3340 1696 3342 1700
rect 3334 1694 3342 1696
rect 3358 1700 3366 1702
rect 3358 1696 3360 1700
rect 3364 1696 3366 1700
rect 3358 1694 3366 1696
rect 3382 1700 3390 1702
rect 3382 1696 3384 1700
rect 3388 1696 3390 1700
rect 3382 1694 3390 1696
rect 3406 1700 3414 1702
rect 3406 1696 3408 1700
rect 3412 1696 3414 1700
rect 3406 1694 3414 1696
rect 3430 1700 3438 1702
rect 3430 1696 3432 1700
rect 3436 1696 3438 1700
rect 3430 1694 3438 1696
rect 3454 1700 3462 1702
rect 3454 1696 3456 1700
rect 3460 1696 3462 1700
rect 3454 1694 3462 1696
rect 3478 1700 3486 1702
rect 3478 1696 3480 1700
rect 3484 1696 3486 1700
rect 3478 1694 3486 1696
rect 3502 1700 3510 1702
rect 3502 1696 3504 1700
rect 3508 1696 3510 1700
rect 3502 1694 3510 1696
rect 3526 1700 3534 1702
rect 3526 1696 3528 1700
rect 3532 1696 3534 1700
rect 3526 1694 3534 1696
rect 3550 1700 3558 1702
rect 3550 1696 3552 1700
rect 3556 1696 3558 1700
rect 3550 1694 3558 1696
rect 3574 1700 3582 1702
rect 3574 1696 3576 1700
rect 3580 1696 3582 1700
rect 3574 1694 3582 1696
rect 3598 1700 3606 1702
rect 3598 1696 3600 1700
rect 3604 1696 3606 1700
rect 3598 1694 3606 1696
rect 3622 1700 3630 1702
rect 3622 1696 3624 1700
rect 3628 1696 3630 1700
rect 3622 1694 3630 1696
rect 3646 1700 3654 1702
rect 3646 1696 3648 1700
rect 3652 1696 3654 1700
rect 3646 1694 3654 1696
rect 3670 1700 3678 1702
rect 3670 1696 3672 1700
rect 3676 1696 3678 1700
rect 3670 1694 3678 1696
rect 3694 1700 3702 1702
rect 3694 1696 3696 1700
rect 3700 1696 3702 1700
rect 3694 1694 3702 1696
rect 3910 1700 3918 1702
rect 3910 1696 3912 1700
rect 3916 1696 3918 1700
rect 3910 1694 3918 1696
rect 3934 1700 3942 1702
rect 3934 1696 3936 1700
rect 3940 1696 3942 1700
rect 3934 1694 3942 1696
rect 3958 1700 3966 1702
rect 3958 1696 3960 1700
rect 3964 1696 3966 1700
rect 3958 1694 3966 1696
rect 3982 1700 3990 1702
rect 3982 1696 3984 1700
rect 3988 1696 3990 1700
rect 3982 1694 3990 1696
rect 4006 1700 4014 1702
rect 4006 1696 4008 1700
rect 4012 1696 4014 1700
rect 4006 1694 4014 1696
rect 4030 1700 4038 1702
rect 4030 1696 4032 1700
rect 4036 1696 4038 1700
rect 4030 1694 4038 1696
rect 4054 1700 4062 1702
rect 4054 1696 4056 1700
rect 4060 1696 4062 1700
rect 4054 1694 4062 1696
rect 4078 1700 4086 1702
rect 4078 1696 4080 1700
rect 4084 1696 4086 1700
rect 4078 1694 4086 1696
rect 4102 1700 4110 1702
rect 4102 1696 4104 1700
rect 4108 1696 4110 1700
rect 4102 1694 4110 1696
rect 4126 1700 4134 1702
rect 4126 1696 4128 1700
rect 4132 1696 4134 1700
rect 4126 1694 4134 1696
rect 4150 1700 4158 1702
rect 4150 1696 4152 1700
rect 4156 1696 4158 1700
rect 4150 1694 4158 1696
rect 4174 1700 4182 1702
rect 4174 1696 4176 1700
rect 4180 1696 4182 1700
rect 4174 1694 4182 1696
rect 4198 1700 4206 1702
rect 4198 1696 4200 1700
rect 4204 1696 4206 1700
rect 4198 1694 4206 1696
rect 4222 1700 4230 1702
rect 4222 1696 4224 1700
rect 4228 1696 4230 1700
rect 4222 1694 4230 1696
rect 4246 1700 4254 1702
rect 4246 1696 4248 1700
rect 4252 1696 4254 1700
rect 4246 1694 4254 1696
rect 4270 1700 4278 1702
rect 4270 1696 4272 1700
rect 4276 1696 4278 1700
rect 4270 1694 4278 1696
rect 4294 1700 4302 1702
rect 4294 1696 4296 1700
rect 4300 1696 4302 1700
rect 4294 1694 4302 1696
rect 4510 1700 4518 1702
rect 4510 1696 4512 1700
rect 4516 1696 4518 1700
rect 4510 1694 4518 1696
rect 4534 1700 4542 1702
rect 4534 1696 4536 1700
rect 4540 1696 4542 1700
rect 4534 1694 4542 1696
rect 4558 1700 4566 1702
rect 4558 1696 4560 1700
rect 4564 1696 4566 1700
rect 4558 1694 4566 1696
rect 4582 1700 4590 1702
rect 4582 1696 4584 1700
rect 4588 1696 4590 1700
rect 4582 1694 4590 1696
rect 4606 1700 4614 1702
rect 4606 1696 4608 1700
rect 4612 1696 4614 1700
rect 4606 1694 4614 1696
rect 4630 1700 4638 1702
rect 4630 1696 4632 1700
rect 4636 1696 4638 1700
rect 4630 1694 4638 1696
rect 4654 1700 4662 1702
rect 4654 1696 4656 1700
rect 4660 1696 4662 1700
rect 4654 1694 4662 1696
rect 4678 1700 4686 1702
rect 4678 1696 4680 1700
rect 4684 1696 4686 1700
rect 4678 1694 4686 1696
rect 4702 1700 4710 1702
rect 4702 1696 4704 1700
rect 4708 1696 4710 1700
rect 4702 1694 4710 1696
rect 4726 1700 4734 1702
rect 4726 1696 4728 1700
rect 4732 1696 4734 1700
rect 4726 1694 4734 1696
rect 4750 1700 4758 1702
rect 4750 1696 4752 1700
rect 4756 1696 4758 1700
rect 4750 1694 4758 1696
rect 4774 1700 4782 1702
rect 4774 1696 4776 1700
rect 4780 1696 4782 1700
rect 4774 1694 4782 1696
rect 4798 1694 4800 1702
rect 5710 1700 5718 1702
rect 5710 1696 5712 1700
rect 5716 1696 5718 1700
rect 5710 1694 5718 1696
rect 5734 1700 5742 1702
rect 5734 1696 5736 1700
rect 5740 1696 5742 1700
rect 5734 1694 5742 1696
rect 5758 1700 5766 1702
rect 5758 1696 5760 1700
rect 5764 1696 5766 1700
rect 5758 1694 5766 1696
rect 5782 1700 5790 1702
rect 5782 1696 5784 1700
rect 5788 1696 5790 1700
rect 5782 1694 5790 1696
rect 5806 1700 5814 1702
rect 5806 1696 5808 1700
rect 5812 1696 5814 1700
rect 5806 1694 5814 1696
rect 5830 1700 5838 1702
rect 5830 1696 5832 1700
rect 5836 1696 5838 1700
rect 5830 1694 5838 1696
rect 5854 1700 5862 1702
rect 5854 1696 5856 1700
rect 5860 1696 5862 1700
rect 5854 1694 5862 1696
rect 5878 1700 5886 1702
rect 5878 1696 5880 1700
rect 5884 1696 5886 1700
rect 5878 1694 5886 1696
rect 5902 1700 5910 1702
rect 5902 1696 5904 1700
rect 5908 1696 5910 1700
rect 5902 1694 5910 1696
rect 5926 1700 5934 1702
rect 5926 1696 5928 1700
rect 5932 1696 5934 1700
rect 5926 1694 5934 1696
rect 5950 1700 5958 1702
rect 5950 1696 5952 1700
rect 5956 1696 5958 1700
rect 5950 1694 5958 1696
rect 5974 1700 5982 1702
rect 5974 1696 5976 1700
rect 5980 1696 5982 1700
rect 5974 1694 5982 1696
rect 5998 1700 6006 1702
rect 5998 1696 6000 1700
rect 6004 1696 6006 1700
rect 5998 1694 6006 1696
rect 6022 1700 6030 1702
rect 6022 1696 6024 1700
rect 6028 1696 6030 1700
rect 6022 1694 6030 1696
rect 6046 1700 6054 1702
rect 6046 1696 6048 1700
rect 6052 1696 6054 1700
rect 6046 1694 6054 1696
rect 6070 1700 6078 1702
rect 6070 1696 6072 1700
rect 6076 1696 6078 1700
rect 6070 1694 6078 1696
rect 6094 1700 6102 1702
rect 6094 1696 6096 1700
rect 6100 1696 6102 1700
rect 6094 1694 6102 1696
rect 6310 1700 6318 1702
rect 6310 1696 6312 1700
rect 6316 1696 6318 1700
rect 6310 1694 6318 1696
rect 6334 1700 6342 1702
rect 6334 1696 6336 1700
rect 6340 1696 6342 1700
rect 6334 1694 6342 1696
rect 6358 1700 6366 1702
rect 6358 1696 6360 1700
rect 6364 1696 6366 1700
rect 6358 1694 6366 1696
rect 6382 1700 6390 1702
rect 6382 1696 6384 1700
rect 6388 1696 6390 1700
rect 6382 1694 6390 1696
rect 6406 1700 6414 1702
rect 6406 1696 6408 1700
rect 6412 1696 6414 1700
rect 6406 1694 6414 1696
rect 6430 1700 6438 1702
rect 6430 1696 6432 1700
rect 6436 1696 6438 1700
rect 6430 1694 6438 1696
rect 6454 1700 6462 1702
rect 6454 1696 6456 1700
rect 6460 1696 6462 1700
rect 6454 1694 6462 1696
rect 6478 1700 6486 1702
rect 6478 1696 6480 1700
rect 6484 1696 6486 1700
rect 6478 1694 6486 1696
rect 6502 1700 6510 1702
rect 6502 1696 6504 1700
rect 6508 1696 6510 1700
rect 6502 1694 6510 1696
rect 6526 1700 6534 1702
rect 6526 1696 6528 1700
rect 6532 1696 6534 1700
rect 6526 1694 6534 1696
rect 6550 1700 6558 1702
rect 6550 1696 6552 1700
rect 6556 1696 6558 1700
rect 6550 1694 6558 1696
rect 6574 1700 6582 1702
rect 6574 1696 6576 1700
rect 6580 1696 6582 1700
rect 6574 1694 6582 1696
rect 6598 1700 6606 1702
rect 6598 1696 6600 1700
rect 6604 1696 6606 1700
rect 6598 1694 6606 1696
rect 6622 1700 6630 1702
rect 6622 1696 6624 1700
rect 6628 1696 6630 1700
rect 6622 1694 6630 1696
rect 6646 1700 6654 1702
rect 6646 1696 6648 1700
rect 6652 1696 6654 1700
rect 6646 1694 6654 1696
rect 6670 1700 6678 1702
rect 6670 1696 6672 1700
rect 6676 1696 6678 1700
rect 6670 1694 6678 1696
rect 6694 1700 6702 1702
rect 6694 1696 6696 1700
rect 6700 1696 6702 1700
rect 6694 1694 6702 1696
rect 6910 1700 6918 1702
rect 6910 1696 6912 1700
rect 6916 1696 6918 1700
rect 6910 1694 6918 1696
rect 6934 1700 6942 1702
rect 6934 1696 6936 1700
rect 6940 1696 6942 1700
rect 6934 1694 6942 1696
rect 6958 1700 6966 1702
rect 6958 1696 6960 1700
rect 6964 1696 6966 1700
rect 6958 1694 6966 1696
rect 6982 1700 6990 1702
rect 6982 1696 6984 1700
rect 6988 1696 6990 1700
rect 6982 1694 6990 1696
rect 7006 1700 7014 1702
rect 7006 1696 7008 1700
rect 7012 1696 7014 1700
rect 7006 1694 7014 1696
rect 7030 1700 7038 1702
rect 7030 1696 7032 1700
rect 7036 1696 7038 1700
rect 7030 1694 7038 1696
rect 7054 1700 7062 1702
rect 7054 1696 7056 1700
rect 7060 1696 7062 1700
rect 7054 1694 7062 1696
rect 7078 1700 7086 1702
rect 7078 1696 7080 1700
rect 7084 1696 7086 1700
rect 7078 1694 7086 1696
rect 7102 1700 7110 1702
rect 7102 1696 7104 1700
rect 7108 1696 7110 1700
rect 7102 1694 7110 1696
rect 7126 1700 7134 1702
rect 7126 1696 7128 1700
rect 7132 1696 7134 1700
rect 7126 1694 7134 1696
rect 7150 1700 7158 1702
rect 7150 1696 7152 1700
rect 7156 1696 7158 1700
rect 7150 1694 7158 1696
rect 7174 1700 7182 1702
rect 7174 1696 7176 1700
rect 7180 1696 7182 1700
rect 7174 1694 7182 1696
rect 7198 1694 7200 1702
rect 2410 1688 2418 1690
rect 2410 1684 2412 1688
rect 2416 1684 2418 1688
rect 2410 1682 2418 1684
rect 2434 1688 2442 1690
rect 2434 1684 2436 1688
rect 2440 1684 2442 1688
rect 2434 1682 2442 1684
rect 2458 1688 2466 1690
rect 2458 1684 2460 1688
rect 2464 1684 2466 1688
rect 2458 1682 2466 1684
rect 2482 1688 2490 1690
rect 2482 1684 2484 1688
rect 2488 1684 2490 1688
rect 2482 1682 2490 1684
rect 2698 1688 2706 1690
rect 2698 1684 2700 1688
rect 2704 1684 2706 1688
rect 2698 1682 2706 1684
rect 2722 1688 2730 1690
rect 2722 1684 2724 1688
rect 2728 1684 2730 1688
rect 2722 1682 2730 1684
rect 2746 1688 2754 1690
rect 2746 1684 2748 1688
rect 2752 1684 2754 1688
rect 2746 1682 2754 1684
rect 2770 1688 2778 1690
rect 2770 1684 2772 1688
rect 2776 1684 2778 1688
rect 2770 1682 2778 1684
rect 2794 1688 2802 1690
rect 2794 1684 2796 1688
rect 2800 1684 2802 1688
rect 2794 1682 2802 1684
rect 2818 1688 2826 1690
rect 2818 1684 2820 1688
rect 2824 1684 2826 1688
rect 2818 1682 2826 1684
rect 2842 1688 2850 1690
rect 2842 1684 2844 1688
rect 2848 1684 2850 1688
rect 2842 1682 2850 1684
rect 2866 1688 2874 1690
rect 2866 1684 2868 1688
rect 2872 1684 2874 1688
rect 2866 1682 2874 1684
rect 2890 1688 2898 1690
rect 2890 1684 2892 1688
rect 2896 1684 2898 1688
rect 2890 1682 2898 1684
rect 2914 1688 2922 1690
rect 2914 1684 2916 1688
rect 2920 1684 2922 1688
rect 2914 1682 2922 1684
rect 2938 1688 2946 1690
rect 2938 1684 2940 1688
rect 2944 1684 2946 1688
rect 2938 1682 2946 1684
rect 2962 1688 2970 1690
rect 2962 1684 2964 1688
rect 2968 1684 2970 1688
rect 2962 1682 2970 1684
rect 2986 1688 2994 1690
rect 2986 1684 2988 1688
rect 2992 1684 2994 1688
rect 2986 1682 2994 1684
rect 3010 1688 3018 1690
rect 3010 1684 3012 1688
rect 3016 1684 3018 1688
rect 3010 1682 3018 1684
rect 3034 1688 3042 1690
rect 3034 1684 3036 1688
rect 3040 1684 3042 1688
rect 3034 1682 3042 1684
rect 3058 1688 3066 1690
rect 3058 1684 3060 1688
rect 3064 1684 3066 1688
rect 3058 1682 3066 1684
rect 3082 1688 3090 1690
rect 3082 1684 3084 1688
rect 3088 1684 3090 1688
rect 3082 1682 3090 1684
rect 3298 1688 3306 1690
rect 3298 1684 3300 1688
rect 3304 1684 3306 1688
rect 3298 1682 3306 1684
rect 3322 1688 3330 1690
rect 3322 1684 3324 1688
rect 3328 1684 3330 1688
rect 3322 1682 3330 1684
rect 3346 1688 3354 1690
rect 3346 1684 3348 1688
rect 3352 1684 3354 1688
rect 3346 1682 3354 1684
rect 3370 1688 3378 1690
rect 3370 1684 3372 1688
rect 3376 1684 3378 1688
rect 3370 1682 3378 1684
rect 3394 1688 3402 1690
rect 3394 1684 3396 1688
rect 3400 1684 3402 1688
rect 3394 1682 3402 1684
rect 3418 1688 3426 1690
rect 3418 1684 3420 1688
rect 3424 1684 3426 1688
rect 3418 1682 3426 1684
rect 3442 1688 3450 1690
rect 3442 1684 3444 1688
rect 3448 1684 3450 1688
rect 3442 1682 3450 1684
rect 3466 1688 3474 1690
rect 3466 1684 3468 1688
rect 3472 1684 3474 1688
rect 3466 1682 3474 1684
rect 3490 1688 3498 1690
rect 3490 1684 3492 1688
rect 3496 1684 3498 1688
rect 3490 1682 3498 1684
rect 3514 1688 3522 1690
rect 3514 1684 3516 1688
rect 3520 1684 3522 1688
rect 3514 1682 3522 1684
rect 3538 1688 3546 1690
rect 3538 1684 3540 1688
rect 3544 1684 3546 1688
rect 3538 1682 3546 1684
rect 3562 1688 3570 1690
rect 3562 1684 3564 1688
rect 3568 1684 3570 1688
rect 3562 1682 3570 1684
rect 3586 1688 3594 1690
rect 3586 1684 3588 1688
rect 3592 1684 3594 1688
rect 3586 1682 3594 1684
rect 3610 1688 3618 1690
rect 3610 1684 3612 1688
rect 3616 1684 3618 1688
rect 3610 1682 3618 1684
rect 3634 1688 3642 1690
rect 3634 1684 3636 1688
rect 3640 1684 3642 1688
rect 3634 1682 3642 1684
rect 3658 1688 3666 1690
rect 3658 1684 3660 1688
rect 3664 1684 3666 1688
rect 3658 1682 3666 1684
rect 3682 1688 3690 1690
rect 3682 1684 3684 1688
rect 3688 1684 3690 1688
rect 3682 1682 3690 1684
rect 3898 1688 3906 1690
rect 3898 1684 3900 1688
rect 3904 1684 3906 1688
rect 3898 1682 3906 1684
rect 3922 1688 3930 1690
rect 3922 1684 3924 1688
rect 3928 1684 3930 1688
rect 3922 1682 3930 1684
rect 3946 1688 3954 1690
rect 3946 1684 3948 1688
rect 3952 1684 3954 1688
rect 3946 1682 3954 1684
rect 3970 1688 3978 1690
rect 3970 1684 3972 1688
rect 3976 1684 3978 1688
rect 3970 1682 3978 1684
rect 3994 1688 4002 1690
rect 3994 1684 3996 1688
rect 4000 1684 4002 1688
rect 3994 1682 4002 1684
rect 4018 1688 4026 1690
rect 4018 1684 4020 1688
rect 4024 1684 4026 1688
rect 4018 1682 4026 1684
rect 4042 1688 4050 1690
rect 4042 1684 4044 1688
rect 4048 1684 4050 1688
rect 4042 1682 4050 1684
rect 4066 1688 4074 1690
rect 4066 1684 4068 1688
rect 4072 1684 4074 1688
rect 4066 1682 4074 1684
rect 4090 1688 4098 1690
rect 4090 1684 4092 1688
rect 4096 1684 4098 1688
rect 4090 1682 4098 1684
rect 4114 1688 4122 1690
rect 4114 1684 4116 1688
rect 4120 1684 4122 1688
rect 4114 1682 4122 1684
rect 4138 1688 4146 1690
rect 4138 1684 4140 1688
rect 4144 1684 4146 1688
rect 4138 1682 4146 1684
rect 4162 1688 4170 1690
rect 4162 1684 4164 1688
rect 4168 1684 4170 1688
rect 4162 1682 4170 1684
rect 4186 1688 4194 1690
rect 4186 1684 4188 1688
rect 4192 1684 4194 1688
rect 4186 1682 4194 1684
rect 4210 1688 4218 1690
rect 4210 1684 4212 1688
rect 4216 1684 4218 1688
rect 4210 1682 4218 1684
rect 4234 1688 4242 1690
rect 4234 1684 4236 1688
rect 4240 1684 4242 1688
rect 4234 1682 4242 1684
rect 4258 1688 4266 1690
rect 4258 1684 4260 1688
rect 4264 1684 4266 1688
rect 4258 1682 4266 1684
rect 4282 1688 4290 1690
rect 4282 1684 4284 1688
rect 4288 1684 4290 1688
rect 4282 1682 4290 1684
rect 4498 1688 4506 1690
rect 4498 1684 4500 1688
rect 4504 1684 4506 1688
rect 4498 1682 4506 1684
rect 4522 1688 4530 1690
rect 4522 1684 4524 1688
rect 4528 1684 4530 1688
rect 4522 1682 4530 1684
rect 4546 1688 4554 1690
rect 4546 1684 4548 1688
rect 4552 1684 4554 1688
rect 4546 1682 4554 1684
rect 4570 1688 4578 1690
rect 4570 1684 4572 1688
rect 4576 1684 4578 1688
rect 4570 1682 4578 1684
rect 4594 1688 4602 1690
rect 4594 1684 4596 1688
rect 4600 1684 4602 1688
rect 4594 1682 4602 1684
rect 4618 1688 4626 1690
rect 4618 1684 4620 1688
rect 4624 1684 4626 1688
rect 4618 1682 4626 1684
rect 4642 1688 4650 1690
rect 4642 1684 4644 1688
rect 4648 1684 4650 1688
rect 4642 1682 4650 1684
rect 4666 1688 4674 1690
rect 4666 1684 4668 1688
rect 4672 1684 4674 1688
rect 4666 1682 4674 1684
rect 4690 1688 4698 1690
rect 4690 1684 4692 1688
rect 4696 1684 4698 1688
rect 4690 1682 4698 1684
rect 4714 1688 4722 1690
rect 4714 1684 4716 1688
rect 4720 1684 4722 1688
rect 4714 1682 4722 1684
rect 4738 1688 4746 1690
rect 4738 1684 4740 1688
rect 4744 1684 4746 1688
rect 4738 1682 4746 1684
rect 4762 1688 4770 1690
rect 4762 1684 4764 1688
rect 4768 1684 4770 1688
rect 4762 1682 4770 1684
rect 4786 1688 4794 1690
rect 4786 1684 4788 1688
rect 4792 1684 4794 1688
rect 4786 1682 4794 1684
rect 5698 1688 5706 1690
rect 5698 1684 5700 1688
rect 5704 1684 5706 1688
rect 5698 1682 5706 1684
rect 5722 1688 5730 1690
rect 5722 1684 5724 1688
rect 5728 1684 5730 1688
rect 5722 1682 5730 1684
rect 5746 1688 5754 1690
rect 5746 1684 5748 1688
rect 5752 1684 5754 1688
rect 5746 1682 5754 1684
rect 5770 1688 5778 1690
rect 5770 1684 5772 1688
rect 5776 1684 5778 1688
rect 5770 1682 5778 1684
rect 5794 1688 5802 1690
rect 5794 1684 5796 1688
rect 5800 1684 5802 1688
rect 5794 1682 5802 1684
rect 5818 1688 5826 1690
rect 5818 1684 5820 1688
rect 5824 1684 5826 1688
rect 5818 1682 5826 1684
rect 5842 1688 5850 1690
rect 5842 1684 5844 1688
rect 5848 1684 5850 1688
rect 5842 1682 5850 1684
rect 5866 1688 5874 1690
rect 5866 1684 5868 1688
rect 5872 1684 5874 1688
rect 5866 1682 5874 1684
rect 5890 1688 5898 1690
rect 5890 1684 5892 1688
rect 5896 1684 5898 1688
rect 5890 1682 5898 1684
rect 5914 1688 5922 1690
rect 5914 1684 5916 1688
rect 5920 1684 5922 1688
rect 5914 1682 5922 1684
rect 5938 1688 5946 1690
rect 5938 1684 5940 1688
rect 5944 1684 5946 1688
rect 5938 1682 5946 1684
rect 5962 1688 5970 1690
rect 5962 1684 5964 1688
rect 5968 1684 5970 1688
rect 5962 1682 5970 1684
rect 5986 1688 5994 1690
rect 5986 1684 5988 1688
rect 5992 1684 5994 1688
rect 5986 1682 5994 1684
rect 6010 1688 6018 1690
rect 6010 1684 6012 1688
rect 6016 1684 6018 1688
rect 6010 1682 6018 1684
rect 6034 1688 6042 1690
rect 6034 1684 6036 1688
rect 6040 1684 6042 1688
rect 6034 1682 6042 1684
rect 6058 1688 6066 1690
rect 6058 1684 6060 1688
rect 6064 1684 6066 1688
rect 6058 1682 6066 1684
rect 6082 1688 6090 1690
rect 6082 1684 6084 1688
rect 6088 1684 6090 1688
rect 6082 1682 6090 1684
rect 6298 1688 6306 1690
rect 6298 1684 6300 1688
rect 6304 1684 6306 1688
rect 6298 1682 6306 1684
rect 6322 1688 6330 1690
rect 6322 1684 6324 1688
rect 6328 1684 6330 1688
rect 6322 1682 6330 1684
rect 6346 1688 6354 1690
rect 6346 1684 6348 1688
rect 6352 1684 6354 1688
rect 6346 1682 6354 1684
rect 6370 1688 6378 1690
rect 6370 1684 6372 1688
rect 6376 1684 6378 1688
rect 6370 1682 6378 1684
rect 6394 1688 6402 1690
rect 6394 1684 6396 1688
rect 6400 1684 6402 1688
rect 6394 1682 6402 1684
rect 6418 1688 6426 1690
rect 6418 1684 6420 1688
rect 6424 1684 6426 1688
rect 6418 1682 6426 1684
rect 6442 1688 6450 1690
rect 6442 1684 6444 1688
rect 6448 1684 6450 1688
rect 6442 1682 6450 1684
rect 6466 1688 6474 1690
rect 6466 1684 6468 1688
rect 6472 1684 6474 1688
rect 6466 1682 6474 1684
rect 6490 1688 6498 1690
rect 6490 1684 6492 1688
rect 6496 1684 6498 1688
rect 6490 1682 6498 1684
rect 6514 1688 6522 1690
rect 6514 1684 6516 1688
rect 6520 1684 6522 1688
rect 6514 1682 6522 1684
rect 6538 1688 6546 1690
rect 6538 1684 6540 1688
rect 6544 1684 6546 1688
rect 6538 1682 6546 1684
rect 6562 1688 6570 1690
rect 6562 1684 6564 1688
rect 6568 1684 6570 1688
rect 6562 1682 6570 1684
rect 6586 1688 6594 1690
rect 6586 1684 6588 1688
rect 6592 1684 6594 1688
rect 6586 1682 6594 1684
rect 6610 1688 6618 1690
rect 6610 1684 6612 1688
rect 6616 1684 6618 1688
rect 6610 1682 6618 1684
rect 6634 1688 6642 1690
rect 6634 1684 6636 1688
rect 6640 1684 6642 1688
rect 6634 1682 6642 1684
rect 6658 1688 6666 1690
rect 6658 1684 6660 1688
rect 6664 1684 6666 1688
rect 6658 1682 6666 1684
rect 6682 1688 6690 1690
rect 6682 1684 6684 1688
rect 6688 1684 6690 1688
rect 6682 1682 6690 1684
rect 6898 1688 6906 1690
rect 6898 1684 6900 1688
rect 6904 1684 6906 1688
rect 6898 1682 6906 1684
rect 6922 1688 6930 1690
rect 6922 1684 6924 1688
rect 6928 1684 6930 1688
rect 6922 1682 6930 1684
rect 6946 1688 6954 1690
rect 6946 1684 6948 1688
rect 6952 1684 6954 1688
rect 6946 1682 6954 1684
rect 6970 1688 6978 1690
rect 6970 1684 6972 1688
rect 6976 1684 6978 1688
rect 6970 1682 6978 1684
rect 6994 1688 7002 1690
rect 6994 1684 6996 1688
rect 7000 1684 7002 1688
rect 6994 1682 7002 1684
rect 7018 1688 7026 1690
rect 7018 1684 7020 1688
rect 7024 1684 7026 1688
rect 7018 1682 7026 1684
rect 7042 1688 7050 1690
rect 7042 1684 7044 1688
rect 7048 1684 7050 1688
rect 7042 1682 7050 1684
rect 7066 1688 7074 1690
rect 7066 1684 7068 1688
rect 7072 1684 7074 1688
rect 7066 1682 7074 1684
rect 7090 1688 7098 1690
rect 7090 1684 7092 1688
rect 7096 1684 7098 1688
rect 7090 1682 7098 1684
rect 7114 1688 7122 1690
rect 7114 1684 7116 1688
rect 7120 1684 7122 1688
rect 7114 1682 7122 1684
rect 7138 1688 7146 1690
rect 7138 1684 7140 1688
rect 7144 1684 7146 1688
rect 7138 1682 7146 1684
rect 7162 1688 7170 1690
rect 7162 1684 7164 1688
rect 7168 1684 7170 1688
rect 7162 1682 7170 1684
rect 7186 1688 7194 1690
rect 7186 1684 7188 1688
rect 7192 1684 7194 1688
rect 7186 1682 7194 1684
rect 2400 1676 2406 1678
rect 2404 1672 2406 1676
rect 2400 1670 2406 1672
rect 2422 1676 2430 1678
rect 2422 1672 2424 1676
rect 2428 1672 2430 1676
rect 2422 1670 2430 1672
rect 2446 1676 2454 1678
rect 2446 1672 2448 1676
rect 2452 1672 2454 1676
rect 2446 1670 2454 1672
rect 2470 1676 2478 1678
rect 2470 1672 2472 1676
rect 2476 1672 2478 1676
rect 2470 1670 2478 1672
rect 2494 1676 2502 1678
rect 2494 1672 2496 1676
rect 2500 1672 2502 1676
rect 2494 1670 2502 1672
rect 2710 1676 2718 1678
rect 2710 1672 2712 1676
rect 2716 1672 2718 1676
rect 2710 1670 2718 1672
rect 2734 1676 2742 1678
rect 2734 1672 2736 1676
rect 2740 1672 2742 1676
rect 2734 1670 2742 1672
rect 2758 1676 2766 1678
rect 2758 1672 2760 1676
rect 2764 1672 2766 1676
rect 2758 1670 2766 1672
rect 2782 1676 2790 1678
rect 2782 1672 2784 1676
rect 2788 1672 2790 1676
rect 2782 1670 2790 1672
rect 2806 1676 2814 1678
rect 2806 1672 2808 1676
rect 2812 1672 2814 1676
rect 2806 1670 2814 1672
rect 2830 1676 2838 1678
rect 2830 1672 2832 1676
rect 2836 1672 2838 1676
rect 2830 1670 2838 1672
rect 2854 1676 2862 1678
rect 2854 1672 2856 1676
rect 2860 1672 2862 1676
rect 2854 1670 2862 1672
rect 2878 1676 2886 1678
rect 2878 1672 2880 1676
rect 2884 1672 2886 1676
rect 2878 1670 2886 1672
rect 2902 1676 2910 1678
rect 2902 1672 2904 1676
rect 2908 1672 2910 1676
rect 2902 1670 2910 1672
rect 2926 1676 2934 1678
rect 2926 1672 2928 1676
rect 2932 1672 2934 1676
rect 2926 1670 2934 1672
rect 2950 1676 2958 1678
rect 2950 1672 2952 1676
rect 2956 1672 2958 1676
rect 2950 1670 2958 1672
rect 2974 1676 2982 1678
rect 2974 1672 2976 1676
rect 2980 1672 2982 1676
rect 2974 1670 2982 1672
rect 2998 1676 3006 1678
rect 2998 1672 3000 1676
rect 3004 1672 3006 1676
rect 2998 1670 3006 1672
rect 3022 1676 3030 1678
rect 3022 1672 3024 1676
rect 3028 1672 3030 1676
rect 3022 1670 3030 1672
rect 3046 1676 3054 1678
rect 3046 1672 3048 1676
rect 3052 1672 3054 1676
rect 3046 1670 3054 1672
rect 3070 1676 3078 1678
rect 3070 1672 3072 1676
rect 3076 1672 3078 1676
rect 3070 1670 3078 1672
rect 3094 1676 3102 1678
rect 3094 1672 3096 1676
rect 3100 1672 3102 1676
rect 3094 1670 3102 1672
rect 3310 1676 3318 1678
rect 3310 1672 3312 1676
rect 3316 1672 3318 1676
rect 3310 1670 3318 1672
rect 3334 1676 3342 1678
rect 3334 1672 3336 1676
rect 3340 1672 3342 1676
rect 3334 1670 3342 1672
rect 3358 1676 3366 1678
rect 3358 1672 3360 1676
rect 3364 1672 3366 1676
rect 3358 1670 3366 1672
rect 3382 1676 3390 1678
rect 3382 1672 3384 1676
rect 3388 1672 3390 1676
rect 3382 1670 3390 1672
rect 3406 1676 3414 1678
rect 3406 1672 3408 1676
rect 3412 1672 3414 1676
rect 3406 1670 3414 1672
rect 3430 1676 3438 1678
rect 3430 1672 3432 1676
rect 3436 1672 3438 1676
rect 3430 1670 3438 1672
rect 3454 1676 3462 1678
rect 3454 1672 3456 1676
rect 3460 1672 3462 1676
rect 3454 1670 3462 1672
rect 3478 1676 3486 1678
rect 3478 1672 3480 1676
rect 3484 1672 3486 1676
rect 3478 1670 3486 1672
rect 3502 1676 3510 1678
rect 3502 1672 3504 1676
rect 3508 1672 3510 1676
rect 3502 1670 3510 1672
rect 3526 1676 3534 1678
rect 3526 1672 3528 1676
rect 3532 1672 3534 1676
rect 3526 1670 3534 1672
rect 3550 1676 3558 1678
rect 3550 1672 3552 1676
rect 3556 1672 3558 1676
rect 3550 1670 3558 1672
rect 3574 1676 3582 1678
rect 3574 1672 3576 1676
rect 3580 1672 3582 1676
rect 3574 1670 3582 1672
rect 3598 1676 3606 1678
rect 3598 1672 3600 1676
rect 3604 1672 3606 1676
rect 3598 1670 3606 1672
rect 3622 1676 3630 1678
rect 3622 1672 3624 1676
rect 3628 1672 3630 1676
rect 3622 1670 3630 1672
rect 3646 1676 3654 1678
rect 3646 1672 3648 1676
rect 3652 1672 3654 1676
rect 3646 1670 3654 1672
rect 3670 1676 3678 1678
rect 3670 1672 3672 1676
rect 3676 1672 3678 1676
rect 3670 1670 3678 1672
rect 3694 1676 3702 1678
rect 3694 1672 3696 1676
rect 3700 1672 3702 1676
rect 3694 1670 3702 1672
rect 3910 1676 3918 1678
rect 3910 1672 3912 1676
rect 3916 1672 3918 1676
rect 3910 1670 3918 1672
rect 3934 1676 3942 1678
rect 3934 1672 3936 1676
rect 3940 1672 3942 1676
rect 3934 1670 3942 1672
rect 3958 1676 3966 1678
rect 3958 1672 3960 1676
rect 3964 1672 3966 1676
rect 3958 1670 3966 1672
rect 3982 1676 3990 1678
rect 3982 1672 3984 1676
rect 3988 1672 3990 1676
rect 3982 1670 3990 1672
rect 4006 1676 4014 1678
rect 4006 1672 4008 1676
rect 4012 1672 4014 1676
rect 4006 1670 4014 1672
rect 4030 1676 4038 1678
rect 4030 1672 4032 1676
rect 4036 1672 4038 1676
rect 4030 1670 4038 1672
rect 4054 1676 4062 1678
rect 4054 1672 4056 1676
rect 4060 1672 4062 1676
rect 4054 1670 4062 1672
rect 4078 1676 4086 1678
rect 4078 1672 4080 1676
rect 4084 1672 4086 1676
rect 4078 1670 4086 1672
rect 4102 1676 4110 1678
rect 4102 1672 4104 1676
rect 4108 1672 4110 1676
rect 4102 1670 4110 1672
rect 4126 1676 4134 1678
rect 4126 1672 4128 1676
rect 4132 1672 4134 1676
rect 4126 1670 4134 1672
rect 4150 1676 4158 1678
rect 4150 1672 4152 1676
rect 4156 1672 4158 1676
rect 4150 1670 4158 1672
rect 4174 1676 4182 1678
rect 4174 1672 4176 1676
rect 4180 1672 4182 1676
rect 4174 1670 4182 1672
rect 4198 1676 4206 1678
rect 4198 1672 4200 1676
rect 4204 1672 4206 1676
rect 4198 1670 4206 1672
rect 4222 1676 4230 1678
rect 4222 1672 4224 1676
rect 4228 1672 4230 1676
rect 4222 1670 4230 1672
rect 4246 1676 4254 1678
rect 4246 1672 4248 1676
rect 4252 1672 4254 1676
rect 4246 1670 4254 1672
rect 4270 1676 4278 1678
rect 4270 1672 4272 1676
rect 4276 1672 4278 1676
rect 4270 1670 4278 1672
rect 4294 1676 4302 1678
rect 4294 1672 4296 1676
rect 4300 1672 4302 1676
rect 4294 1670 4302 1672
rect 4510 1676 4518 1678
rect 4510 1672 4512 1676
rect 4516 1672 4518 1676
rect 4510 1670 4518 1672
rect 4534 1676 4542 1678
rect 4534 1672 4536 1676
rect 4540 1672 4542 1676
rect 4534 1670 4542 1672
rect 4558 1676 4566 1678
rect 4558 1672 4560 1676
rect 4564 1672 4566 1676
rect 4558 1670 4566 1672
rect 4582 1676 4590 1678
rect 4582 1672 4584 1676
rect 4588 1672 4590 1676
rect 4582 1670 4590 1672
rect 4606 1676 4614 1678
rect 4606 1672 4608 1676
rect 4612 1672 4614 1676
rect 4606 1670 4614 1672
rect 4630 1676 4638 1678
rect 4630 1672 4632 1676
rect 4636 1672 4638 1676
rect 4630 1670 4638 1672
rect 4654 1676 4662 1678
rect 4654 1672 4656 1676
rect 4660 1672 4662 1676
rect 4654 1670 4662 1672
rect 4678 1676 4686 1678
rect 4678 1672 4680 1676
rect 4684 1672 4686 1676
rect 4678 1670 4686 1672
rect 4702 1676 4710 1678
rect 4702 1672 4704 1676
rect 4708 1672 4710 1676
rect 4702 1670 4710 1672
rect 4726 1676 4734 1678
rect 4726 1672 4728 1676
rect 4732 1672 4734 1676
rect 4726 1670 4734 1672
rect 4750 1676 4758 1678
rect 4750 1672 4752 1676
rect 4756 1672 4758 1676
rect 4750 1670 4758 1672
rect 4774 1676 4782 1678
rect 4774 1672 4776 1676
rect 4780 1672 4782 1676
rect 4774 1670 4782 1672
rect 4798 1670 4800 1678
rect 5710 1676 5718 1678
rect 5710 1672 5712 1676
rect 5716 1672 5718 1676
rect 5710 1670 5718 1672
rect 5734 1676 5742 1678
rect 5734 1672 5736 1676
rect 5740 1672 5742 1676
rect 5734 1670 5742 1672
rect 5758 1676 5766 1678
rect 5758 1672 5760 1676
rect 5764 1672 5766 1676
rect 5758 1670 5766 1672
rect 5782 1676 5790 1678
rect 5782 1672 5784 1676
rect 5788 1672 5790 1676
rect 5782 1670 5790 1672
rect 5806 1676 5814 1678
rect 5806 1672 5808 1676
rect 5812 1672 5814 1676
rect 5806 1670 5814 1672
rect 5830 1676 5838 1678
rect 5830 1672 5832 1676
rect 5836 1672 5838 1676
rect 5830 1670 5838 1672
rect 5854 1676 5862 1678
rect 5854 1672 5856 1676
rect 5860 1672 5862 1676
rect 5854 1670 5862 1672
rect 5878 1676 5886 1678
rect 5878 1672 5880 1676
rect 5884 1672 5886 1676
rect 5878 1670 5886 1672
rect 5902 1676 5910 1678
rect 5902 1672 5904 1676
rect 5908 1672 5910 1676
rect 5902 1670 5910 1672
rect 5926 1676 5934 1678
rect 5926 1672 5928 1676
rect 5932 1672 5934 1676
rect 5926 1670 5934 1672
rect 5950 1676 5958 1678
rect 5950 1672 5952 1676
rect 5956 1672 5958 1676
rect 5950 1670 5958 1672
rect 5974 1676 5982 1678
rect 5974 1672 5976 1676
rect 5980 1672 5982 1676
rect 5974 1670 5982 1672
rect 5998 1676 6006 1678
rect 5998 1672 6000 1676
rect 6004 1672 6006 1676
rect 5998 1670 6006 1672
rect 6022 1676 6030 1678
rect 6022 1672 6024 1676
rect 6028 1672 6030 1676
rect 6022 1670 6030 1672
rect 6046 1676 6054 1678
rect 6046 1672 6048 1676
rect 6052 1672 6054 1676
rect 6046 1670 6054 1672
rect 6070 1676 6078 1678
rect 6070 1672 6072 1676
rect 6076 1672 6078 1676
rect 6070 1670 6078 1672
rect 6094 1676 6102 1678
rect 6094 1672 6096 1676
rect 6100 1672 6102 1676
rect 6094 1670 6102 1672
rect 6310 1676 6318 1678
rect 6310 1672 6312 1676
rect 6316 1672 6318 1676
rect 6310 1670 6318 1672
rect 6334 1676 6342 1678
rect 6334 1672 6336 1676
rect 6340 1672 6342 1676
rect 6334 1670 6342 1672
rect 6358 1676 6366 1678
rect 6358 1672 6360 1676
rect 6364 1672 6366 1676
rect 6358 1670 6366 1672
rect 6382 1676 6390 1678
rect 6382 1672 6384 1676
rect 6388 1672 6390 1676
rect 6382 1670 6390 1672
rect 6406 1676 6414 1678
rect 6406 1672 6408 1676
rect 6412 1672 6414 1676
rect 6406 1670 6414 1672
rect 6430 1676 6438 1678
rect 6430 1672 6432 1676
rect 6436 1672 6438 1676
rect 6430 1670 6438 1672
rect 6454 1676 6462 1678
rect 6454 1672 6456 1676
rect 6460 1672 6462 1676
rect 6454 1670 6462 1672
rect 6478 1676 6486 1678
rect 6478 1672 6480 1676
rect 6484 1672 6486 1676
rect 6478 1670 6486 1672
rect 6502 1676 6510 1678
rect 6502 1672 6504 1676
rect 6508 1672 6510 1676
rect 6502 1670 6510 1672
rect 6526 1676 6534 1678
rect 6526 1672 6528 1676
rect 6532 1672 6534 1676
rect 6526 1670 6534 1672
rect 6550 1676 6558 1678
rect 6550 1672 6552 1676
rect 6556 1672 6558 1676
rect 6550 1670 6558 1672
rect 6574 1676 6582 1678
rect 6574 1672 6576 1676
rect 6580 1672 6582 1676
rect 6574 1670 6582 1672
rect 6598 1676 6606 1678
rect 6598 1672 6600 1676
rect 6604 1672 6606 1676
rect 6598 1670 6606 1672
rect 6622 1676 6630 1678
rect 6622 1672 6624 1676
rect 6628 1672 6630 1676
rect 6622 1670 6630 1672
rect 6646 1676 6654 1678
rect 6646 1672 6648 1676
rect 6652 1672 6654 1676
rect 6646 1670 6654 1672
rect 6670 1676 6678 1678
rect 6670 1672 6672 1676
rect 6676 1672 6678 1676
rect 6670 1670 6678 1672
rect 6694 1676 6702 1678
rect 6694 1672 6696 1676
rect 6700 1672 6702 1676
rect 6694 1670 6702 1672
rect 6910 1676 6918 1678
rect 6910 1672 6912 1676
rect 6916 1672 6918 1676
rect 6910 1670 6918 1672
rect 6934 1676 6942 1678
rect 6934 1672 6936 1676
rect 6940 1672 6942 1676
rect 6934 1670 6942 1672
rect 6958 1676 6966 1678
rect 6958 1672 6960 1676
rect 6964 1672 6966 1676
rect 6958 1670 6966 1672
rect 6982 1676 6990 1678
rect 6982 1672 6984 1676
rect 6988 1672 6990 1676
rect 6982 1670 6990 1672
rect 7006 1676 7014 1678
rect 7006 1672 7008 1676
rect 7012 1672 7014 1676
rect 7006 1670 7014 1672
rect 7030 1676 7038 1678
rect 7030 1672 7032 1676
rect 7036 1672 7038 1676
rect 7030 1670 7038 1672
rect 7054 1676 7062 1678
rect 7054 1672 7056 1676
rect 7060 1672 7062 1676
rect 7054 1670 7062 1672
rect 7078 1676 7086 1678
rect 7078 1672 7080 1676
rect 7084 1672 7086 1676
rect 7078 1670 7086 1672
rect 7102 1676 7110 1678
rect 7102 1672 7104 1676
rect 7108 1672 7110 1676
rect 7102 1670 7110 1672
rect 7126 1676 7134 1678
rect 7126 1672 7128 1676
rect 7132 1672 7134 1676
rect 7126 1670 7134 1672
rect 7150 1676 7158 1678
rect 7150 1672 7152 1676
rect 7156 1672 7158 1676
rect 7150 1670 7158 1672
rect 7174 1676 7182 1678
rect 7174 1672 7176 1676
rect 7180 1672 7182 1676
rect 7174 1670 7182 1672
rect 7198 1670 7200 1678
rect 2410 1664 2418 1666
rect 2410 1660 2412 1664
rect 2416 1660 2418 1664
rect 2410 1658 2418 1660
rect 2434 1664 2442 1666
rect 2434 1660 2436 1664
rect 2440 1660 2442 1664
rect 2434 1658 2442 1660
rect 2458 1664 2466 1666
rect 2458 1660 2460 1664
rect 2464 1660 2466 1664
rect 2458 1658 2466 1660
rect 2482 1664 2490 1666
rect 2482 1660 2484 1664
rect 2488 1660 2490 1664
rect 2482 1658 2490 1660
rect 2698 1664 2706 1666
rect 2698 1660 2700 1664
rect 2704 1660 2706 1664
rect 2698 1658 2706 1660
rect 2722 1664 2730 1666
rect 2722 1660 2724 1664
rect 2728 1660 2730 1664
rect 2722 1658 2730 1660
rect 2746 1664 2754 1666
rect 2746 1660 2748 1664
rect 2752 1660 2754 1664
rect 2746 1658 2754 1660
rect 2770 1664 2778 1666
rect 2770 1660 2772 1664
rect 2776 1660 2778 1664
rect 2770 1658 2778 1660
rect 2794 1664 2802 1666
rect 2794 1660 2796 1664
rect 2800 1660 2802 1664
rect 2794 1658 2802 1660
rect 2818 1664 2826 1666
rect 2818 1660 2820 1664
rect 2824 1660 2826 1664
rect 2818 1658 2826 1660
rect 2842 1664 2850 1666
rect 2842 1660 2844 1664
rect 2848 1660 2850 1664
rect 2842 1658 2850 1660
rect 2866 1664 2874 1666
rect 2866 1660 2868 1664
rect 2872 1660 2874 1664
rect 2866 1658 2874 1660
rect 2890 1664 2898 1666
rect 2890 1660 2892 1664
rect 2896 1660 2898 1664
rect 2890 1658 2898 1660
rect 2914 1664 2922 1666
rect 2914 1660 2916 1664
rect 2920 1660 2922 1664
rect 2914 1658 2922 1660
rect 2938 1664 2946 1666
rect 2938 1660 2940 1664
rect 2944 1660 2946 1664
rect 2938 1658 2946 1660
rect 2962 1664 2970 1666
rect 2962 1660 2964 1664
rect 2968 1660 2970 1664
rect 2962 1658 2970 1660
rect 2986 1664 2994 1666
rect 2986 1660 2988 1664
rect 2992 1660 2994 1664
rect 2986 1658 2994 1660
rect 3010 1664 3018 1666
rect 3010 1660 3012 1664
rect 3016 1660 3018 1664
rect 3010 1658 3018 1660
rect 3034 1664 3042 1666
rect 3034 1660 3036 1664
rect 3040 1660 3042 1664
rect 3034 1658 3042 1660
rect 3058 1664 3066 1666
rect 3058 1660 3060 1664
rect 3064 1660 3066 1664
rect 3058 1658 3066 1660
rect 3082 1664 3090 1666
rect 3082 1660 3084 1664
rect 3088 1660 3090 1664
rect 3082 1658 3090 1660
rect 3298 1664 3306 1666
rect 3298 1660 3300 1664
rect 3304 1660 3306 1664
rect 3298 1658 3306 1660
rect 3322 1664 3330 1666
rect 3322 1660 3324 1664
rect 3328 1660 3330 1664
rect 3322 1658 3330 1660
rect 3346 1664 3354 1666
rect 3346 1660 3348 1664
rect 3352 1660 3354 1664
rect 3346 1658 3354 1660
rect 3370 1664 3378 1666
rect 3370 1660 3372 1664
rect 3376 1660 3378 1664
rect 3370 1658 3378 1660
rect 3394 1664 3402 1666
rect 3394 1660 3396 1664
rect 3400 1660 3402 1664
rect 3394 1658 3402 1660
rect 3418 1664 3426 1666
rect 3418 1660 3420 1664
rect 3424 1660 3426 1664
rect 3418 1658 3426 1660
rect 3442 1664 3450 1666
rect 3442 1660 3444 1664
rect 3448 1660 3450 1664
rect 3442 1658 3450 1660
rect 3466 1664 3474 1666
rect 3466 1660 3468 1664
rect 3472 1660 3474 1664
rect 3466 1658 3474 1660
rect 3490 1664 3498 1666
rect 3490 1660 3492 1664
rect 3496 1660 3498 1664
rect 3490 1658 3498 1660
rect 3514 1664 3522 1666
rect 3514 1660 3516 1664
rect 3520 1660 3522 1664
rect 3514 1658 3522 1660
rect 3538 1664 3546 1666
rect 3538 1660 3540 1664
rect 3544 1660 3546 1664
rect 3538 1658 3546 1660
rect 3562 1664 3570 1666
rect 3562 1660 3564 1664
rect 3568 1660 3570 1664
rect 3562 1658 3570 1660
rect 3586 1664 3594 1666
rect 3586 1660 3588 1664
rect 3592 1660 3594 1664
rect 3586 1658 3594 1660
rect 3610 1664 3618 1666
rect 3610 1660 3612 1664
rect 3616 1660 3618 1664
rect 3610 1658 3618 1660
rect 3634 1664 3642 1666
rect 3634 1660 3636 1664
rect 3640 1660 3642 1664
rect 3634 1658 3642 1660
rect 3658 1664 3666 1666
rect 3658 1660 3660 1664
rect 3664 1660 3666 1664
rect 3658 1658 3666 1660
rect 3682 1664 3690 1666
rect 3682 1660 3684 1664
rect 3688 1660 3690 1664
rect 3682 1658 3690 1660
rect 3898 1664 3906 1666
rect 3898 1660 3900 1664
rect 3904 1660 3906 1664
rect 3898 1658 3906 1660
rect 3922 1664 3930 1666
rect 3922 1660 3924 1664
rect 3928 1660 3930 1664
rect 3922 1658 3930 1660
rect 3946 1664 3954 1666
rect 3946 1660 3948 1664
rect 3952 1660 3954 1664
rect 3946 1658 3954 1660
rect 3970 1664 3978 1666
rect 3970 1660 3972 1664
rect 3976 1660 3978 1664
rect 3970 1658 3978 1660
rect 3994 1664 4002 1666
rect 3994 1660 3996 1664
rect 4000 1660 4002 1664
rect 3994 1658 4002 1660
rect 4018 1664 4026 1666
rect 4018 1660 4020 1664
rect 4024 1660 4026 1664
rect 4018 1658 4026 1660
rect 4042 1664 4050 1666
rect 4042 1660 4044 1664
rect 4048 1660 4050 1664
rect 4042 1658 4050 1660
rect 4066 1664 4074 1666
rect 4066 1660 4068 1664
rect 4072 1660 4074 1664
rect 4066 1658 4074 1660
rect 4090 1664 4098 1666
rect 4090 1660 4092 1664
rect 4096 1660 4098 1664
rect 4090 1658 4098 1660
rect 4114 1664 4122 1666
rect 4114 1660 4116 1664
rect 4120 1660 4122 1664
rect 4114 1658 4122 1660
rect 4138 1664 4146 1666
rect 4138 1660 4140 1664
rect 4144 1660 4146 1664
rect 4138 1658 4146 1660
rect 4162 1664 4170 1666
rect 4162 1660 4164 1664
rect 4168 1660 4170 1664
rect 4162 1658 4170 1660
rect 4186 1664 4194 1666
rect 4186 1660 4188 1664
rect 4192 1660 4194 1664
rect 4186 1658 4194 1660
rect 4210 1664 4218 1666
rect 4210 1660 4212 1664
rect 4216 1660 4218 1664
rect 4210 1658 4218 1660
rect 4234 1664 4242 1666
rect 4234 1660 4236 1664
rect 4240 1660 4242 1664
rect 4234 1658 4242 1660
rect 4258 1664 4266 1666
rect 4258 1660 4260 1664
rect 4264 1660 4266 1664
rect 4258 1658 4266 1660
rect 4282 1664 4290 1666
rect 4282 1660 4284 1664
rect 4288 1660 4290 1664
rect 4282 1658 4290 1660
rect 4498 1664 4506 1666
rect 4498 1660 4500 1664
rect 4504 1660 4506 1664
rect 4498 1658 4506 1660
rect 4522 1664 4530 1666
rect 4522 1660 4524 1664
rect 4528 1660 4530 1664
rect 4522 1658 4530 1660
rect 4546 1664 4554 1666
rect 4546 1660 4548 1664
rect 4552 1660 4554 1664
rect 4546 1658 4554 1660
rect 4570 1664 4578 1666
rect 4570 1660 4572 1664
rect 4576 1660 4578 1664
rect 4570 1658 4578 1660
rect 4594 1664 4602 1666
rect 4594 1660 4596 1664
rect 4600 1660 4602 1664
rect 4594 1658 4602 1660
rect 4618 1664 4626 1666
rect 4618 1660 4620 1664
rect 4624 1660 4626 1664
rect 4618 1658 4626 1660
rect 4642 1664 4650 1666
rect 4642 1660 4644 1664
rect 4648 1660 4650 1664
rect 4642 1658 4650 1660
rect 4666 1664 4674 1666
rect 4666 1660 4668 1664
rect 4672 1660 4674 1664
rect 4666 1658 4674 1660
rect 4690 1664 4698 1666
rect 4690 1660 4692 1664
rect 4696 1660 4698 1664
rect 4690 1658 4698 1660
rect 4714 1664 4722 1666
rect 4714 1660 4716 1664
rect 4720 1660 4722 1664
rect 4714 1658 4722 1660
rect 4738 1664 4746 1666
rect 4738 1660 4740 1664
rect 4744 1660 4746 1664
rect 4738 1658 4746 1660
rect 4762 1664 4770 1666
rect 4762 1660 4764 1664
rect 4768 1660 4770 1664
rect 4762 1658 4770 1660
rect 4786 1664 4794 1666
rect 4786 1660 4788 1664
rect 4792 1660 4794 1664
rect 4786 1658 4794 1660
rect 5698 1664 5706 1666
rect 5698 1660 5700 1664
rect 5704 1660 5706 1664
rect 5698 1658 5706 1660
rect 5722 1664 5730 1666
rect 5722 1660 5724 1664
rect 5728 1660 5730 1664
rect 5722 1658 5730 1660
rect 5746 1664 5754 1666
rect 5746 1660 5748 1664
rect 5752 1660 5754 1664
rect 5746 1658 5754 1660
rect 5770 1664 5778 1666
rect 5770 1660 5772 1664
rect 5776 1660 5778 1664
rect 5770 1658 5778 1660
rect 5794 1664 5802 1666
rect 5794 1660 5796 1664
rect 5800 1660 5802 1664
rect 5794 1658 5802 1660
rect 5818 1664 5826 1666
rect 5818 1660 5820 1664
rect 5824 1660 5826 1664
rect 5818 1658 5826 1660
rect 5842 1664 5850 1666
rect 5842 1660 5844 1664
rect 5848 1660 5850 1664
rect 5842 1658 5850 1660
rect 5866 1664 5874 1666
rect 5866 1660 5868 1664
rect 5872 1660 5874 1664
rect 5866 1658 5874 1660
rect 5890 1664 5898 1666
rect 5890 1660 5892 1664
rect 5896 1660 5898 1664
rect 5890 1658 5898 1660
rect 5914 1664 5922 1666
rect 5914 1660 5916 1664
rect 5920 1660 5922 1664
rect 5914 1658 5922 1660
rect 5938 1664 5946 1666
rect 5938 1660 5940 1664
rect 5944 1660 5946 1664
rect 5938 1658 5946 1660
rect 5962 1664 5970 1666
rect 5962 1660 5964 1664
rect 5968 1660 5970 1664
rect 5962 1658 5970 1660
rect 5986 1664 5994 1666
rect 5986 1660 5988 1664
rect 5992 1660 5994 1664
rect 5986 1658 5994 1660
rect 6010 1664 6018 1666
rect 6010 1660 6012 1664
rect 6016 1660 6018 1664
rect 6010 1658 6018 1660
rect 6034 1664 6042 1666
rect 6034 1660 6036 1664
rect 6040 1660 6042 1664
rect 6034 1658 6042 1660
rect 6058 1664 6066 1666
rect 6058 1660 6060 1664
rect 6064 1660 6066 1664
rect 6058 1658 6066 1660
rect 6082 1664 6090 1666
rect 6082 1660 6084 1664
rect 6088 1660 6090 1664
rect 6082 1658 6090 1660
rect 6298 1664 6306 1666
rect 6298 1660 6300 1664
rect 6304 1660 6306 1664
rect 6298 1658 6306 1660
rect 6322 1664 6330 1666
rect 6322 1660 6324 1664
rect 6328 1660 6330 1664
rect 6322 1658 6330 1660
rect 6346 1664 6354 1666
rect 6346 1660 6348 1664
rect 6352 1660 6354 1664
rect 6346 1658 6354 1660
rect 6370 1664 6378 1666
rect 6370 1660 6372 1664
rect 6376 1660 6378 1664
rect 6370 1658 6378 1660
rect 6394 1664 6402 1666
rect 6394 1660 6396 1664
rect 6400 1660 6402 1664
rect 6394 1658 6402 1660
rect 6418 1664 6426 1666
rect 6418 1660 6420 1664
rect 6424 1660 6426 1664
rect 6418 1658 6426 1660
rect 6442 1664 6450 1666
rect 6442 1660 6444 1664
rect 6448 1660 6450 1664
rect 6442 1658 6450 1660
rect 6466 1664 6474 1666
rect 6466 1660 6468 1664
rect 6472 1660 6474 1664
rect 6466 1658 6474 1660
rect 6490 1664 6498 1666
rect 6490 1660 6492 1664
rect 6496 1660 6498 1664
rect 6490 1658 6498 1660
rect 6514 1664 6522 1666
rect 6514 1660 6516 1664
rect 6520 1660 6522 1664
rect 6514 1658 6522 1660
rect 6538 1664 6546 1666
rect 6538 1660 6540 1664
rect 6544 1660 6546 1664
rect 6538 1658 6546 1660
rect 6562 1664 6570 1666
rect 6562 1660 6564 1664
rect 6568 1660 6570 1664
rect 6562 1658 6570 1660
rect 6586 1664 6594 1666
rect 6586 1660 6588 1664
rect 6592 1660 6594 1664
rect 6586 1658 6594 1660
rect 6610 1664 6618 1666
rect 6610 1660 6612 1664
rect 6616 1660 6618 1664
rect 6610 1658 6618 1660
rect 6634 1664 6642 1666
rect 6634 1660 6636 1664
rect 6640 1660 6642 1664
rect 6634 1658 6642 1660
rect 6658 1664 6666 1666
rect 6658 1660 6660 1664
rect 6664 1660 6666 1664
rect 6658 1658 6666 1660
rect 6682 1664 6690 1666
rect 6682 1660 6684 1664
rect 6688 1660 6690 1664
rect 6682 1658 6690 1660
rect 6898 1664 6906 1666
rect 6898 1660 6900 1664
rect 6904 1660 6906 1664
rect 6898 1658 6906 1660
rect 6922 1664 6930 1666
rect 6922 1660 6924 1664
rect 6928 1660 6930 1664
rect 6922 1658 6930 1660
rect 6946 1664 6954 1666
rect 6946 1660 6948 1664
rect 6952 1660 6954 1664
rect 6946 1658 6954 1660
rect 6970 1664 6978 1666
rect 6970 1660 6972 1664
rect 6976 1660 6978 1664
rect 6970 1658 6978 1660
rect 6994 1664 7002 1666
rect 6994 1660 6996 1664
rect 7000 1660 7002 1664
rect 6994 1658 7002 1660
rect 7018 1664 7026 1666
rect 7018 1660 7020 1664
rect 7024 1660 7026 1664
rect 7018 1658 7026 1660
rect 7042 1664 7050 1666
rect 7042 1660 7044 1664
rect 7048 1660 7050 1664
rect 7042 1658 7050 1660
rect 7066 1664 7074 1666
rect 7066 1660 7068 1664
rect 7072 1660 7074 1664
rect 7066 1658 7074 1660
rect 7090 1664 7098 1666
rect 7090 1660 7092 1664
rect 7096 1660 7098 1664
rect 7090 1658 7098 1660
rect 7114 1664 7122 1666
rect 7114 1660 7116 1664
rect 7120 1660 7122 1664
rect 7114 1658 7122 1660
rect 7138 1664 7146 1666
rect 7138 1660 7140 1664
rect 7144 1660 7146 1664
rect 7138 1658 7146 1660
rect 7162 1664 7170 1666
rect 7162 1660 7164 1664
rect 7168 1660 7170 1664
rect 7162 1658 7170 1660
rect 7186 1664 7194 1666
rect 7186 1660 7188 1664
rect 7192 1660 7194 1664
rect 7186 1658 7194 1660
rect 2400 1652 2406 1654
rect 2404 1648 2406 1652
rect 2400 1646 2406 1648
rect 2422 1652 2430 1654
rect 2422 1648 2424 1652
rect 2428 1648 2430 1652
rect 2422 1646 2430 1648
rect 2446 1652 2454 1654
rect 2446 1648 2448 1652
rect 2452 1648 2454 1652
rect 2446 1646 2454 1648
rect 2470 1652 2478 1654
rect 2470 1648 2472 1652
rect 2476 1648 2478 1652
rect 2470 1646 2478 1648
rect 2494 1652 2502 1654
rect 2494 1648 2496 1652
rect 2500 1648 2502 1652
rect 2494 1646 2502 1648
rect 2710 1652 2718 1654
rect 2710 1648 2712 1652
rect 2716 1648 2718 1652
rect 2710 1646 2718 1648
rect 2734 1652 2742 1654
rect 2734 1648 2736 1652
rect 2740 1648 2742 1652
rect 2734 1646 2742 1648
rect 2758 1652 2766 1654
rect 2758 1648 2760 1652
rect 2764 1648 2766 1652
rect 2758 1646 2766 1648
rect 2782 1652 2790 1654
rect 2782 1648 2784 1652
rect 2788 1648 2790 1652
rect 2782 1646 2790 1648
rect 2806 1652 2814 1654
rect 2806 1648 2808 1652
rect 2812 1648 2814 1652
rect 2806 1646 2814 1648
rect 2830 1652 2838 1654
rect 2830 1648 2832 1652
rect 2836 1648 2838 1652
rect 2830 1646 2838 1648
rect 2854 1652 2862 1654
rect 2854 1648 2856 1652
rect 2860 1648 2862 1652
rect 2854 1646 2862 1648
rect 2878 1652 2886 1654
rect 2878 1648 2880 1652
rect 2884 1648 2886 1652
rect 2878 1646 2886 1648
rect 2902 1652 2910 1654
rect 2902 1648 2904 1652
rect 2908 1648 2910 1652
rect 2902 1646 2910 1648
rect 2926 1652 2934 1654
rect 2926 1648 2928 1652
rect 2932 1648 2934 1652
rect 2926 1646 2934 1648
rect 2950 1652 2958 1654
rect 2950 1648 2952 1652
rect 2956 1648 2958 1652
rect 2950 1646 2958 1648
rect 2974 1652 2982 1654
rect 2974 1648 2976 1652
rect 2980 1648 2982 1652
rect 2974 1646 2982 1648
rect 2998 1652 3006 1654
rect 2998 1648 3000 1652
rect 3004 1648 3006 1652
rect 2998 1646 3006 1648
rect 3022 1652 3030 1654
rect 3022 1648 3024 1652
rect 3028 1648 3030 1652
rect 3022 1646 3030 1648
rect 3046 1652 3054 1654
rect 3046 1648 3048 1652
rect 3052 1648 3054 1652
rect 3046 1646 3054 1648
rect 3070 1652 3078 1654
rect 3070 1648 3072 1652
rect 3076 1648 3078 1652
rect 3070 1646 3078 1648
rect 3094 1652 3102 1654
rect 3094 1648 3096 1652
rect 3100 1648 3102 1652
rect 3094 1646 3102 1648
rect 3310 1652 3318 1654
rect 3310 1648 3312 1652
rect 3316 1648 3318 1652
rect 3310 1646 3318 1648
rect 3334 1652 3342 1654
rect 3334 1648 3336 1652
rect 3340 1648 3342 1652
rect 3334 1646 3342 1648
rect 3358 1652 3366 1654
rect 3358 1648 3360 1652
rect 3364 1648 3366 1652
rect 3358 1646 3366 1648
rect 3382 1652 3390 1654
rect 3382 1648 3384 1652
rect 3388 1648 3390 1652
rect 3382 1646 3390 1648
rect 3406 1652 3414 1654
rect 3406 1648 3408 1652
rect 3412 1648 3414 1652
rect 3406 1646 3414 1648
rect 3430 1652 3438 1654
rect 3430 1648 3432 1652
rect 3436 1648 3438 1652
rect 3430 1646 3438 1648
rect 3454 1652 3462 1654
rect 3454 1648 3456 1652
rect 3460 1648 3462 1652
rect 3454 1646 3462 1648
rect 3478 1652 3486 1654
rect 3478 1648 3480 1652
rect 3484 1648 3486 1652
rect 3478 1646 3486 1648
rect 3502 1652 3510 1654
rect 3502 1648 3504 1652
rect 3508 1648 3510 1652
rect 3502 1646 3510 1648
rect 3526 1652 3534 1654
rect 3526 1648 3528 1652
rect 3532 1648 3534 1652
rect 3526 1646 3534 1648
rect 3550 1652 3558 1654
rect 3550 1648 3552 1652
rect 3556 1648 3558 1652
rect 3550 1646 3558 1648
rect 3574 1652 3582 1654
rect 3574 1648 3576 1652
rect 3580 1648 3582 1652
rect 3574 1646 3582 1648
rect 3598 1652 3606 1654
rect 3598 1648 3600 1652
rect 3604 1648 3606 1652
rect 3598 1646 3606 1648
rect 3622 1652 3630 1654
rect 3622 1648 3624 1652
rect 3628 1648 3630 1652
rect 3622 1646 3630 1648
rect 3646 1652 3654 1654
rect 3646 1648 3648 1652
rect 3652 1648 3654 1652
rect 3646 1646 3654 1648
rect 3670 1652 3678 1654
rect 3670 1648 3672 1652
rect 3676 1648 3678 1652
rect 3670 1646 3678 1648
rect 3694 1652 3702 1654
rect 3694 1648 3696 1652
rect 3700 1648 3702 1652
rect 3694 1646 3702 1648
rect 3910 1652 3918 1654
rect 3910 1648 3912 1652
rect 3916 1648 3918 1652
rect 3910 1646 3918 1648
rect 3934 1652 3942 1654
rect 3934 1648 3936 1652
rect 3940 1648 3942 1652
rect 3934 1646 3942 1648
rect 3958 1652 3966 1654
rect 3958 1648 3960 1652
rect 3964 1648 3966 1652
rect 3958 1646 3966 1648
rect 3982 1652 3990 1654
rect 3982 1648 3984 1652
rect 3988 1648 3990 1652
rect 3982 1646 3990 1648
rect 4006 1652 4014 1654
rect 4006 1648 4008 1652
rect 4012 1648 4014 1652
rect 4006 1646 4014 1648
rect 4030 1652 4038 1654
rect 4030 1648 4032 1652
rect 4036 1648 4038 1652
rect 4030 1646 4038 1648
rect 4054 1652 4062 1654
rect 4054 1648 4056 1652
rect 4060 1648 4062 1652
rect 4054 1646 4062 1648
rect 4078 1652 4086 1654
rect 4078 1648 4080 1652
rect 4084 1648 4086 1652
rect 4078 1646 4086 1648
rect 4102 1652 4110 1654
rect 4102 1648 4104 1652
rect 4108 1648 4110 1652
rect 4102 1646 4110 1648
rect 4126 1652 4134 1654
rect 4126 1648 4128 1652
rect 4132 1648 4134 1652
rect 4126 1646 4134 1648
rect 4150 1652 4158 1654
rect 4150 1648 4152 1652
rect 4156 1648 4158 1652
rect 4150 1646 4158 1648
rect 4174 1652 4182 1654
rect 4174 1648 4176 1652
rect 4180 1648 4182 1652
rect 4174 1646 4182 1648
rect 4198 1652 4206 1654
rect 4198 1648 4200 1652
rect 4204 1648 4206 1652
rect 4198 1646 4206 1648
rect 4222 1652 4230 1654
rect 4222 1648 4224 1652
rect 4228 1648 4230 1652
rect 4222 1646 4230 1648
rect 4246 1652 4254 1654
rect 4246 1648 4248 1652
rect 4252 1648 4254 1652
rect 4246 1646 4254 1648
rect 4270 1652 4278 1654
rect 4270 1648 4272 1652
rect 4276 1648 4278 1652
rect 4270 1646 4278 1648
rect 4294 1652 4302 1654
rect 4294 1648 4296 1652
rect 4300 1648 4302 1652
rect 4294 1646 4302 1648
rect 4510 1652 4518 1654
rect 4510 1648 4512 1652
rect 4516 1648 4518 1652
rect 4510 1646 4518 1648
rect 4534 1652 4542 1654
rect 4534 1648 4536 1652
rect 4540 1648 4542 1652
rect 4534 1646 4542 1648
rect 4558 1652 4566 1654
rect 4558 1648 4560 1652
rect 4564 1648 4566 1652
rect 4558 1646 4566 1648
rect 4582 1652 4590 1654
rect 4582 1648 4584 1652
rect 4588 1648 4590 1652
rect 4582 1646 4590 1648
rect 4606 1652 4614 1654
rect 4606 1648 4608 1652
rect 4612 1648 4614 1652
rect 4606 1646 4614 1648
rect 4630 1652 4638 1654
rect 4630 1648 4632 1652
rect 4636 1648 4638 1652
rect 4630 1646 4638 1648
rect 4654 1652 4662 1654
rect 4654 1648 4656 1652
rect 4660 1648 4662 1652
rect 4654 1646 4662 1648
rect 4678 1652 4686 1654
rect 4678 1648 4680 1652
rect 4684 1648 4686 1652
rect 4678 1646 4686 1648
rect 4702 1652 4710 1654
rect 4702 1648 4704 1652
rect 4708 1648 4710 1652
rect 4702 1646 4710 1648
rect 4726 1652 4734 1654
rect 4726 1648 4728 1652
rect 4732 1648 4734 1652
rect 4726 1646 4734 1648
rect 4750 1652 4758 1654
rect 4750 1648 4752 1652
rect 4756 1648 4758 1652
rect 4750 1646 4758 1648
rect 4774 1652 4782 1654
rect 4774 1648 4776 1652
rect 4780 1648 4782 1652
rect 4774 1646 4782 1648
rect 4798 1646 4800 1654
rect 5710 1652 5718 1654
rect 5710 1648 5712 1652
rect 5716 1648 5718 1652
rect 5710 1646 5718 1648
rect 5734 1652 5742 1654
rect 5734 1648 5736 1652
rect 5740 1648 5742 1652
rect 5734 1646 5742 1648
rect 5758 1652 5766 1654
rect 5758 1648 5760 1652
rect 5764 1648 5766 1652
rect 5758 1646 5766 1648
rect 5782 1652 5790 1654
rect 5782 1648 5784 1652
rect 5788 1648 5790 1652
rect 5782 1646 5790 1648
rect 5806 1652 5814 1654
rect 5806 1648 5808 1652
rect 5812 1648 5814 1652
rect 5806 1646 5814 1648
rect 5830 1652 5838 1654
rect 5830 1648 5832 1652
rect 5836 1648 5838 1652
rect 5830 1646 5838 1648
rect 5854 1652 5862 1654
rect 5854 1648 5856 1652
rect 5860 1648 5862 1652
rect 5854 1646 5862 1648
rect 5878 1652 5886 1654
rect 5878 1648 5880 1652
rect 5884 1648 5886 1652
rect 5878 1646 5886 1648
rect 5902 1652 5910 1654
rect 5902 1648 5904 1652
rect 5908 1648 5910 1652
rect 5902 1646 5910 1648
rect 5926 1652 5934 1654
rect 5926 1648 5928 1652
rect 5932 1648 5934 1652
rect 5926 1646 5934 1648
rect 5950 1652 5958 1654
rect 5950 1648 5952 1652
rect 5956 1648 5958 1652
rect 5950 1646 5958 1648
rect 5974 1652 5982 1654
rect 5974 1648 5976 1652
rect 5980 1648 5982 1652
rect 5974 1646 5982 1648
rect 5998 1652 6006 1654
rect 5998 1648 6000 1652
rect 6004 1648 6006 1652
rect 5998 1646 6006 1648
rect 6022 1652 6030 1654
rect 6022 1648 6024 1652
rect 6028 1648 6030 1652
rect 6022 1646 6030 1648
rect 6046 1652 6054 1654
rect 6046 1648 6048 1652
rect 6052 1648 6054 1652
rect 6046 1646 6054 1648
rect 6070 1652 6078 1654
rect 6070 1648 6072 1652
rect 6076 1648 6078 1652
rect 6070 1646 6078 1648
rect 6094 1652 6102 1654
rect 6094 1648 6096 1652
rect 6100 1648 6102 1652
rect 6094 1646 6102 1648
rect 6310 1652 6318 1654
rect 6310 1648 6312 1652
rect 6316 1648 6318 1652
rect 6310 1646 6318 1648
rect 6334 1652 6342 1654
rect 6334 1648 6336 1652
rect 6340 1648 6342 1652
rect 6334 1646 6342 1648
rect 6358 1652 6366 1654
rect 6358 1648 6360 1652
rect 6364 1648 6366 1652
rect 6358 1646 6366 1648
rect 6382 1652 6390 1654
rect 6382 1648 6384 1652
rect 6388 1648 6390 1652
rect 6382 1646 6390 1648
rect 6406 1652 6414 1654
rect 6406 1648 6408 1652
rect 6412 1648 6414 1652
rect 6406 1646 6414 1648
rect 6430 1652 6438 1654
rect 6430 1648 6432 1652
rect 6436 1648 6438 1652
rect 6430 1646 6438 1648
rect 6454 1652 6462 1654
rect 6454 1648 6456 1652
rect 6460 1648 6462 1652
rect 6454 1646 6462 1648
rect 6478 1652 6486 1654
rect 6478 1648 6480 1652
rect 6484 1648 6486 1652
rect 6478 1646 6486 1648
rect 6502 1652 6510 1654
rect 6502 1648 6504 1652
rect 6508 1648 6510 1652
rect 6502 1646 6510 1648
rect 6526 1652 6534 1654
rect 6526 1648 6528 1652
rect 6532 1648 6534 1652
rect 6526 1646 6534 1648
rect 6550 1652 6558 1654
rect 6550 1648 6552 1652
rect 6556 1648 6558 1652
rect 6550 1646 6558 1648
rect 6574 1652 6582 1654
rect 6574 1648 6576 1652
rect 6580 1648 6582 1652
rect 6574 1646 6582 1648
rect 6598 1652 6606 1654
rect 6598 1648 6600 1652
rect 6604 1648 6606 1652
rect 6598 1646 6606 1648
rect 6622 1652 6630 1654
rect 6622 1648 6624 1652
rect 6628 1648 6630 1652
rect 6622 1646 6630 1648
rect 6646 1652 6654 1654
rect 6646 1648 6648 1652
rect 6652 1648 6654 1652
rect 6646 1646 6654 1648
rect 6670 1652 6678 1654
rect 6670 1648 6672 1652
rect 6676 1648 6678 1652
rect 6670 1646 6678 1648
rect 6694 1652 6702 1654
rect 6694 1648 6696 1652
rect 6700 1648 6702 1652
rect 6694 1646 6702 1648
rect 6910 1652 6918 1654
rect 6910 1648 6912 1652
rect 6916 1648 6918 1652
rect 6910 1646 6918 1648
rect 6934 1652 6942 1654
rect 6934 1648 6936 1652
rect 6940 1648 6942 1652
rect 6934 1646 6942 1648
rect 6958 1652 6966 1654
rect 6958 1648 6960 1652
rect 6964 1648 6966 1652
rect 6958 1646 6966 1648
rect 6982 1652 6990 1654
rect 6982 1648 6984 1652
rect 6988 1648 6990 1652
rect 6982 1646 6990 1648
rect 7006 1652 7014 1654
rect 7006 1648 7008 1652
rect 7012 1648 7014 1652
rect 7006 1646 7014 1648
rect 7030 1652 7038 1654
rect 7030 1648 7032 1652
rect 7036 1648 7038 1652
rect 7030 1646 7038 1648
rect 7054 1652 7062 1654
rect 7054 1648 7056 1652
rect 7060 1648 7062 1652
rect 7054 1646 7062 1648
rect 7078 1652 7086 1654
rect 7078 1648 7080 1652
rect 7084 1648 7086 1652
rect 7078 1646 7086 1648
rect 7102 1652 7110 1654
rect 7102 1648 7104 1652
rect 7108 1648 7110 1652
rect 7102 1646 7110 1648
rect 7126 1652 7134 1654
rect 7126 1648 7128 1652
rect 7132 1648 7134 1652
rect 7126 1646 7134 1648
rect 7150 1652 7158 1654
rect 7150 1648 7152 1652
rect 7156 1648 7158 1652
rect 7150 1646 7158 1648
rect 7174 1652 7182 1654
rect 7174 1648 7176 1652
rect 7180 1648 7182 1652
rect 7174 1646 7182 1648
rect 7198 1646 7200 1654
rect 2410 1640 2418 1642
rect 2410 1636 2412 1640
rect 2416 1636 2418 1640
rect 2410 1634 2418 1636
rect 2434 1640 2442 1642
rect 2434 1636 2436 1640
rect 2440 1636 2442 1640
rect 2434 1634 2442 1636
rect 2458 1640 2466 1642
rect 2458 1636 2460 1640
rect 2464 1636 2466 1640
rect 2458 1634 2466 1636
rect 2482 1640 2490 1642
rect 2482 1636 2484 1640
rect 2488 1636 2490 1640
rect 2482 1634 2490 1636
rect 2698 1640 2706 1642
rect 2698 1636 2700 1640
rect 2704 1636 2706 1640
rect 2698 1634 2706 1636
rect 2722 1640 2730 1642
rect 2722 1636 2724 1640
rect 2728 1636 2730 1640
rect 2722 1634 2730 1636
rect 2746 1640 2754 1642
rect 2746 1636 2748 1640
rect 2752 1636 2754 1640
rect 2746 1634 2754 1636
rect 2770 1640 2778 1642
rect 2770 1636 2772 1640
rect 2776 1636 2778 1640
rect 2770 1634 2778 1636
rect 2794 1640 2802 1642
rect 2794 1636 2796 1640
rect 2800 1636 2802 1640
rect 2794 1634 2802 1636
rect 2818 1640 2826 1642
rect 2818 1636 2820 1640
rect 2824 1636 2826 1640
rect 2818 1634 2826 1636
rect 2842 1640 2850 1642
rect 2842 1636 2844 1640
rect 2848 1636 2850 1640
rect 2842 1634 2850 1636
rect 2866 1640 2874 1642
rect 2866 1636 2868 1640
rect 2872 1636 2874 1640
rect 2866 1634 2874 1636
rect 2890 1640 2898 1642
rect 2890 1636 2892 1640
rect 2896 1636 2898 1640
rect 2890 1634 2898 1636
rect 2914 1640 2922 1642
rect 2914 1636 2916 1640
rect 2920 1636 2922 1640
rect 2914 1634 2922 1636
rect 2938 1640 2946 1642
rect 2938 1636 2940 1640
rect 2944 1636 2946 1640
rect 2938 1634 2946 1636
rect 2962 1640 2970 1642
rect 2962 1636 2964 1640
rect 2968 1636 2970 1640
rect 2962 1634 2970 1636
rect 2986 1640 2994 1642
rect 2986 1636 2988 1640
rect 2992 1636 2994 1640
rect 2986 1634 2994 1636
rect 3010 1640 3018 1642
rect 3010 1636 3012 1640
rect 3016 1636 3018 1640
rect 3010 1634 3018 1636
rect 3034 1640 3042 1642
rect 3034 1636 3036 1640
rect 3040 1636 3042 1640
rect 3034 1634 3042 1636
rect 3058 1640 3066 1642
rect 3058 1636 3060 1640
rect 3064 1636 3066 1640
rect 3058 1634 3066 1636
rect 3082 1640 3090 1642
rect 3082 1636 3084 1640
rect 3088 1636 3090 1640
rect 3082 1634 3090 1636
rect 3298 1640 3306 1642
rect 3298 1636 3300 1640
rect 3304 1636 3306 1640
rect 3298 1634 3306 1636
rect 3322 1640 3330 1642
rect 3322 1636 3324 1640
rect 3328 1636 3330 1640
rect 3322 1634 3330 1636
rect 3346 1640 3354 1642
rect 3346 1636 3348 1640
rect 3352 1636 3354 1640
rect 3346 1634 3354 1636
rect 3370 1640 3378 1642
rect 3370 1636 3372 1640
rect 3376 1636 3378 1640
rect 3370 1634 3378 1636
rect 3394 1640 3402 1642
rect 3394 1636 3396 1640
rect 3400 1636 3402 1640
rect 3394 1634 3402 1636
rect 3418 1640 3426 1642
rect 3418 1636 3420 1640
rect 3424 1636 3426 1640
rect 3418 1634 3426 1636
rect 3442 1640 3450 1642
rect 3442 1636 3444 1640
rect 3448 1636 3450 1640
rect 3442 1634 3450 1636
rect 3466 1640 3474 1642
rect 3466 1636 3468 1640
rect 3472 1636 3474 1640
rect 3466 1634 3474 1636
rect 3490 1640 3498 1642
rect 3490 1636 3492 1640
rect 3496 1636 3498 1640
rect 3490 1634 3498 1636
rect 3514 1640 3522 1642
rect 3514 1636 3516 1640
rect 3520 1636 3522 1640
rect 3514 1634 3522 1636
rect 3538 1640 3546 1642
rect 3538 1636 3540 1640
rect 3544 1636 3546 1640
rect 3538 1634 3546 1636
rect 3562 1640 3570 1642
rect 3562 1636 3564 1640
rect 3568 1636 3570 1640
rect 3562 1634 3570 1636
rect 3586 1640 3594 1642
rect 3586 1636 3588 1640
rect 3592 1636 3594 1640
rect 3586 1634 3594 1636
rect 3610 1640 3618 1642
rect 3610 1636 3612 1640
rect 3616 1636 3618 1640
rect 3610 1634 3618 1636
rect 3634 1640 3642 1642
rect 3634 1636 3636 1640
rect 3640 1636 3642 1640
rect 3634 1634 3642 1636
rect 3658 1640 3666 1642
rect 3658 1636 3660 1640
rect 3664 1636 3666 1640
rect 3658 1634 3666 1636
rect 3682 1640 3690 1642
rect 3682 1636 3684 1640
rect 3688 1636 3690 1640
rect 3682 1634 3690 1636
rect 3898 1640 3906 1642
rect 3898 1636 3900 1640
rect 3904 1636 3906 1640
rect 3898 1634 3906 1636
rect 3922 1640 3930 1642
rect 3922 1636 3924 1640
rect 3928 1636 3930 1640
rect 3922 1634 3930 1636
rect 3946 1640 3954 1642
rect 3946 1636 3948 1640
rect 3952 1636 3954 1640
rect 3946 1634 3954 1636
rect 3970 1640 3978 1642
rect 3970 1636 3972 1640
rect 3976 1636 3978 1640
rect 3970 1634 3978 1636
rect 3994 1640 4002 1642
rect 3994 1636 3996 1640
rect 4000 1636 4002 1640
rect 3994 1634 4002 1636
rect 4018 1640 4026 1642
rect 4018 1636 4020 1640
rect 4024 1636 4026 1640
rect 4018 1634 4026 1636
rect 4042 1640 4050 1642
rect 4042 1636 4044 1640
rect 4048 1636 4050 1640
rect 4042 1634 4050 1636
rect 4066 1640 4074 1642
rect 4066 1636 4068 1640
rect 4072 1636 4074 1640
rect 4066 1634 4074 1636
rect 4090 1640 4098 1642
rect 4090 1636 4092 1640
rect 4096 1636 4098 1640
rect 4090 1634 4098 1636
rect 4114 1640 4122 1642
rect 4114 1636 4116 1640
rect 4120 1636 4122 1640
rect 4114 1634 4122 1636
rect 4138 1640 4146 1642
rect 4138 1636 4140 1640
rect 4144 1636 4146 1640
rect 4138 1634 4146 1636
rect 4162 1640 4170 1642
rect 4162 1636 4164 1640
rect 4168 1636 4170 1640
rect 4162 1634 4170 1636
rect 4186 1640 4194 1642
rect 4186 1636 4188 1640
rect 4192 1636 4194 1640
rect 4186 1634 4194 1636
rect 4210 1640 4218 1642
rect 4210 1636 4212 1640
rect 4216 1636 4218 1640
rect 4210 1634 4218 1636
rect 4234 1640 4242 1642
rect 4234 1636 4236 1640
rect 4240 1636 4242 1640
rect 4234 1634 4242 1636
rect 4258 1640 4266 1642
rect 4258 1636 4260 1640
rect 4264 1636 4266 1640
rect 4258 1634 4266 1636
rect 4282 1640 4290 1642
rect 4282 1636 4284 1640
rect 4288 1636 4290 1640
rect 4282 1634 4290 1636
rect 4498 1640 4506 1642
rect 4498 1636 4500 1640
rect 4504 1636 4506 1640
rect 4498 1634 4506 1636
rect 4522 1640 4530 1642
rect 4522 1636 4524 1640
rect 4528 1636 4530 1640
rect 4522 1634 4530 1636
rect 4546 1640 4554 1642
rect 4546 1636 4548 1640
rect 4552 1636 4554 1640
rect 4546 1634 4554 1636
rect 4570 1640 4578 1642
rect 4570 1636 4572 1640
rect 4576 1636 4578 1640
rect 4570 1634 4578 1636
rect 4594 1640 4602 1642
rect 4594 1636 4596 1640
rect 4600 1636 4602 1640
rect 4594 1634 4602 1636
rect 4618 1640 4626 1642
rect 4618 1636 4620 1640
rect 4624 1636 4626 1640
rect 4618 1634 4626 1636
rect 4642 1640 4650 1642
rect 4642 1636 4644 1640
rect 4648 1636 4650 1640
rect 4642 1634 4650 1636
rect 4666 1640 4674 1642
rect 4666 1636 4668 1640
rect 4672 1636 4674 1640
rect 4666 1634 4674 1636
rect 4690 1640 4698 1642
rect 4690 1636 4692 1640
rect 4696 1636 4698 1640
rect 4690 1634 4698 1636
rect 4714 1640 4722 1642
rect 4714 1636 4716 1640
rect 4720 1636 4722 1640
rect 4714 1634 4722 1636
rect 4738 1640 4746 1642
rect 4738 1636 4740 1640
rect 4744 1636 4746 1640
rect 4738 1634 4746 1636
rect 4762 1640 4770 1642
rect 4762 1636 4764 1640
rect 4768 1636 4770 1640
rect 4762 1634 4770 1636
rect 4786 1640 4794 1642
rect 4786 1636 4788 1640
rect 4792 1636 4794 1640
rect 4786 1634 4794 1636
rect 5698 1640 5706 1642
rect 5698 1636 5700 1640
rect 5704 1636 5706 1640
rect 5698 1634 5706 1636
rect 5722 1640 5730 1642
rect 5722 1636 5724 1640
rect 5728 1636 5730 1640
rect 5722 1634 5730 1636
rect 5746 1640 5754 1642
rect 5746 1636 5748 1640
rect 5752 1636 5754 1640
rect 5746 1634 5754 1636
rect 5770 1640 5778 1642
rect 5770 1636 5772 1640
rect 5776 1636 5778 1640
rect 5770 1634 5778 1636
rect 5794 1640 5802 1642
rect 5794 1636 5796 1640
rect 5800 1636 5802 1640
rect 5794 1634 5802 1636
rect 5818 1640 5826 1642
rect 5818 1636 5820 1640
rect 5824 1636 5826 1640
rect 5818 1634 5826 1636
rect 5842 1640 5850 1642
rect 5842 1636 5844 1640
rect 5848 1636 5850 1640
rect 5842 1634 5850 1636
rect 5866 1640 5874 1642
rect 5866 1636 5868 1640
rect 5872 1636 5874 1640
rect 5866 1634 5874 1636
rect 5890 1640 5898 1642
rect 5890 1636 5892 1640
rect 5896 1636 5898 1640
rect 5890 1634 5898 1636
rect 5914 1640 5922 1642
rect 5914 1636 5916 1640
rect 5920 1636 5922 1640
rect 5914 1634 5922 1636
rect 5938 1640 5946 1642
rect 5938 1636 5940 1640
rect 5944 1636 5946 1640
rect 5938 1634 5946 1636
rect 5962 1640 5970 1642
rect 5962 1636 5964 1640
rect 5968 1636 5970 1640
rect 5962 1634 5970 1636
rect 5986 1640 5994 1642
rect 5986 1636 5988 1640
rect 5992 1636 5994 1640
rect 5986 1634 5994 1636
rect 6010 1640 6018 1642
rect 6010 1636 6012 1640
rect 6016 1636 6018 1640
rect 6010 1634 6018 1636
rect 6034 1640 6042 1642
rect 6034 1636 6036 1640
rect 6040 1636 6042 1640
rect 6034 1634 6042 1636
rect 6058 1640 6066 1642
rect 6058 1636 6060 1640
rect 6064 1636 6066 1640
rect 6058 1634 6066 1636
rect 6082 1640 6090 1642
rect 6082 1636 6084 1640
rect 6088 1636 6090 1640
rect 6082 1634 6090 1636
rect 6298 1640 6306 1642
rect 6298 1636 6300 1640
rect 6304 1636 6306 1640
rect 6298 1634 6306 1636
rect 6322 1640 6330 1642
rect 6322 1636 6324 1640
rect 6328 1636 6330 1640
rect 6322 1634 6330 1636
rect 6346 1640 6354 1642
rect 6346 1636 6348 1640
rect 6352 1636 6354 1640
rect 6346 1634 6354 1636
rect 6370 1640 6378 1642
rect 6370 1636 6372 1640
rect 6376 1636 6378 1640
rect 6370 1634 6378 1636
rect 6394 1640 6402 1642
rect 6394 1636 6396 1640
rect 6400 1636 6402 1640
rect 6394 1634 6402 1636
rect 6418 1640 6426 1642
rect 6418 1636 6420 1640
rect 6424 1636 6426 1640
rect 6418 1634 6426 1636
rect 6442 1640 6450 1642
rect 6442 1636 6444 1640
rect 6448 1636 6450 1640
rect 6442 1634 6450 1636
rect 6466 1640 6474 1642
rect 6466 1636 6468 1640
rect 6472 1636 6474 1640
rect 6466 1634 6474 1636
rect 6490 1640 6498 1642
rect 6490 1636 6492 1640
rect 6496 1636 6498 1640
rect 6490 1634 6498 1636
rect 6514 1640 6522 1642
rect 6514 1636 6516 1640
rect 6520 1636 6522 1640
rect 6514 1634 6522 1636
rect 6538 1640 6546 1642
rect 6538 1636 6540 1640
rect 6544 1636 6546 1640
rect 6538 1634 6546 1636
rect 6562 1640 6570 1642
rect 6562 1636 6564 1640
rect 6568 1636 6570 1640
rect 6562 1634 6570 1636
rect 6586 1640 6594 1642
rect 6586 1636 6588 1640
rect 6592 1636 6594 1640
rect 6586 1634 6594 1636
rect 6610 1640 6618 1642
rect 6610 1636 6612 1640
rect 6616 1636 6618 1640
rect 6610 1634 6618 1636
rect 6634 1640 6642 1642
rect 6634 1636 6636 1640
rect 6640 1636 6642 1640
rect 6634 1634 6642 1636
rect 6658 1640 6666 1642
rect 6658 1636 6660 1640
rect 6664 1636 6666 1640
rect 6658 1634 6666 1636
rect 6682 1640 6690 1642
rect 6682 1636 6684 1640
rect 6688 1636 6690 1640
rect 6682 1634 6690 1636
rect 6898 1640 6906 1642
rect 6898 1636 6900 1640
rect 6904 1636 6906 1640
rect 6898 1634 6906 1636
rect 6922 1640 6930 1642
rect 6922 1636 6924 1640
rect 6928 1636 6930 1640
rect 6922 1634 6930 1636
rect 6946 1640 6954 1642
rect 6946 1636 6948 1640
rect 6952 1636 6954 1640
rect 6946 1634 6954 1636
rect 6970 1640 6978 1642
rect 6970 1636 6972 1640
rect 6976 1636 6978 1640
rect 6970 1634 6978 1636
rect 6994 1640 7002 1642
rect 6994 1636 6996 1640
rect 7000 1636 7002 1640
rect 6994 1634 7002 1636
rect 7018 1640 7026 1642
rect 7018 1636 7020 1640
rect 7024 1636 7026 1640
rect 7018 1634 7026 1636
rect 7042 1640 7050 1642
rect 7042 1636 7044 1640
rect 7048 1636 7050 1640
rect 7042 1634 7050 1636
rect 7066 1640 7074 1642
rect 7066 1636 7068 1640
rect 7072 1636 7074 1640
rect 7066 1634 7074 1636
rect 7090 1640 7098 1642
rect 7090 1636 7092 1640
rect 7096 1636 7098 1640
rect 7090 1634 7098 1636
rect 7114 1640 7122 1642
rect 7114 1636 7116 1640
rect 7120 1636 7122 1640
rect 7114 1634 7122 1636
rect 7138 1640 7146 1642
rect 7138 1636 7140 1640
rect 7144 1636 7146 1640
rect 7138 1634 7146 1636
rect 7162 1640 7170 1642
rect 7162 1636 7164 1640
rect 7168 1636 7170 1640
rect 7162 1634 7170 1636
rect 7186 1640 7194 1642
rect 7186 1636 7188 1640
rect 7192 1636 7194 1640
rect 7186 1634 7194 1636
rect 2400 1628 2406 1630
rect 2404 1624 2406 1628
rect 2400 1622 2406 1624
rect 2422 1628 2430 1630
rect 2422 1624 2424 1628
rect 2428 1624 2430 1628
rect 2422 1622 2430 1624
rect 2446 1628 2454 1630
rect 2446 1624 2448 1628
rect 2452 1624 2454 1628
rect 2446 1622 2454 1624
rect 2470 1628 2478 1630
rect 2470 1624 2472 1628
rect 2476 1624 2478 1628
rect 2470 1622 2478 1624
rect 2494 1628 2502 1630
rect 2494 1624 2496 1628
rect 2500 1624 2502 1628
rect 2494 1622 2502 1624
rect 2710 1628 2718 1630
rect 2710 1624 2712 1628
rect 2716 1624 2718 1628
rect 2710 1622 2718 1624
rect 2734 1628 2742 1630
rect 2734 1624 2736 1628
rect 2740 1624 2742 1628
rect 2734 1622 2742 1624
rect 2758 1628 2766 1630
rect 2758 1624 2760 1628
rect 2764 1624 2766 1628
rect 2758 1622 2766 1624
rect 2782 1628 2790 1630
rect 2782 1624 2784 1628
rect 2788 1624 2790 1628
rect 2782 1622 2790 1624
rect 2806 1628 2814 1630
rect 2806 1624 2808 1628
rect 2812 1624 2814 1628
rect 2806 1622 2814 1624
rect 2830 1628 2838 1630
rect 2830 1624 2832 1628
rect 2836 1624 2838 1628
rect 2830 1622 2838 1624
rect 2854 1628 2862 1630
rect 2854 1624 2856 1628
rect 2860 1624 2862 1628
rect 2854 1622 2862 1624
rect 2878 1628 2886 1630
rect 2878 1624 2880 1628
rect 2884 1624 2886 1628
rect 2878 1622 2886 1624
rect 2902 1628 2910 1630
rect 2902 1624 2904 1628
rect 2908 1624 2910 1628
rect 2902 1622 2910 1624
rect 2926 1628 2934 1630
rect 2926 1624 2928 1628
rect 2932 1624 2934 1628
rect 2926 1622 2934 1624
rect 2950 1628 2958 1630
rect 2950 1624 2952 1628
rect 2956 1624 2958 1628
rect 2950 1622 2958 1624
rect 2974 1628 2982 1630
rect 2974 1624 2976 1628
rect 2980 1624 2982 1628
rect 2974 1622 2982 1624
rect 2998 1628 3006 1630
rect 2998 1624 3000 1628
rect 3004 1624 3006 1628
rect 2998 1622 3006 1624
rect 3022 1628 3030 1630
rect 3022 1624 3024 1628
rect 3028 1624 3030 1628
rect 3022 1622 3030 1624
rect 3046 1628 3054 1630
rect 3046 1624 3048 1628
rect 3052 1624 3054 1628
rect 3046 1622 3054 1624
rect 3070 1628 3078 1630
rect 3070 1624 3072 1628
rect 3076 1624 3078 1628
rect 3070 1622 3078 1624
rect 3094 1628 3102 1630
rect 3094 1624 3096 1628
rect 3100 1624 3102 1628
rect 3094 1622 3102 1624
rect 3310 1628 3318 1630
rect 3310 1624 3312 1628
rect 3316 1624 3318 1628
rect 3310 1622 3318 1624
rect 3334 1628 3342 1630
rect 3334 1624 3336 1628
rect 3340 1624 3342 1628
rect 3334 1622 3342 1624
rect 3358 1628 3366 1630
rect 3358 1624 3360 1628
rect 3364 1624 3366 1628
rect 3358 1622 3366 1624
rect 3382 1628 3390 1630
rect 3382 1624 3384 1628
rect 3388 1624 3390 1628
rect 3382 1622 3390 1624
rect 3406 1628 3414 1630
rect 3406 1624 3408 1628
rect 3412 1624 3414 1628
rect 3406 1622 3414 1624
rect 3430 1628 3438 1630
rect 3430 1624 3432 1628
rect 3436 1624 3438 1628
rect 3430 1622 3438 1624
rect 3454 1628 3462 1630
rect 3454 1624 3456 1628
rect 3460 1624 3462 1628
rect 3454 1622 3462 1624
rect 3478 1628 3486 1630
rect 3478 1624 3480 1628
rect 3484 1624 3486 1628
rect 3478 1622 3486 1624
rect 3502 1628 3510 1630
rect 3502 1624 3504 1628
rect 3508 1624 3510 1628
rect 3502 1622 3510 1624
rect 3526 1628 3534 1630
rect 3526 1624 3528 1628
rect 3532 1624 3534 1628
rect 3526 1622 3534 1624
rect 3550 1628 3558 1630
rect 3550 1624 3552 1628
rect 3556 1624 3558 1628
rect 3550 1622 3558 1624
rect 3574 1628 3582 1630
rect 3574 1624 3576 1628
rect 3580 1624 3582 1628
rect 3574 1622 3582 1624
rect 3598 1628 3606 1630
rect 3598 1624 3600 1628
rect 3604 1624 3606 1628
rect 3598 1622 3606 1624
rect 3622 1628 3630 1630
rect 3622 1624 3624 1628
rect 3628 1624 3630 1628
rect 3622 1622 3630 1624
rect 3646 1628 3654 1630
rect 3646 1624 3648 1628
rect 3652 1624 3654 1628
rect 3646 1622 3654 1624
rect 3670 1628 3678 1630
rect 3670 1624 3672 1628
rect 3676 1624 3678 1628
rect 3670 1622 3678 1624
rect 3694 1628 3702 1630
rect 3694 1624 3696 1628
rect 3700 1624 3702 1628
rect 3694 1622 3702 1624
rect 3910 1628 3918 1630
rect 3910 1624 3912 1628
rect 3916 1624 3918 1628
rect 3910 1622 3918 1624
rect 3934 1628 3942 1630
rect 3934 1624 3936 1628
rect 3940 1624 3942 1628
rect 3934 1622 3942 1624
rect 3958 1628 3966 1630
rect 3958 1624 3960 1628
rect 3964 1624 3966 1628
rect 3958 1622 3966 1624
rect 3982 1628 3990 1630
rect 3982 1624 3984 1628
rect 3988 1624 3990 1628
rect 3982 1622 3990 1624
rect 4006 1628 4014 1630
rect 4006 1624 4008 1628
rect 4012 1624 4014 1628
rect 4006 1622 4014 1624
rect 4030 1628 4038 1630
rect 4030 1624 4032 1628
rect 4036 1624 4038 1628
rect 4030 1622 4038 1624
rect 4054 1628 4062 1630
rect 4054 1624 4056 1628
rect 4060 1624 4062 1628
rect 4054 1622 4062 1624
rect 4078 1628 4086 1630
rect 4078 1624 4080 1628
rect 4084 1624 4086 1628
rect 4078 1622 4086 1624
rect 4102 1628 4110 1630
rect 4102 1624 4104 1628
rect 4108 1624 4110 1628
rect 4102 1622 4110 1624
rect 4126 1628 4134 1630
rect 4126 1624 4128 1628
rect 4132 1624 4134 1628
rect 4126 1622 4134 1624
rect 4150 1628 4158 1630
rect 4150 1624 4152 1628
rect 4156 1624 4158 1628
rect 4150 1622 4158 1624
rect 4174 1628 4182 1630
rect 4174 1624 4176 1628
rect 4180 1624 4182 1628
rect 4174 1622 4182 1624
rect 4198 1628 4206 1630
rect 4198 1624 4200 1628
rect 4204 1624 4206 1628
rect 4198 1622 4206 1624
rect 4222 1628 4230 1630
rect 4222 1624 4224 1628
rect 4228 1624 4230 1628
rect 4222 1622 4230 1624
rect 4246 1628 4254 1630
rect 4246 1624 4248 1628
rect 4252 1624 4254 1628
rect 4246 1622 4254 1624
rect 4270 1628 4278 1630
rect 4270 1624 4272 1628
rect 4276 1624 4278 1628
rect 4270 1622 4278 1624
rect 4294 1628 4302 1630
rect 4294 1624 4296 1628
rect 4300 1624 4302 1628
rect 4294 1622 4302 1624
rect 4510 1628 4518 1630
rect 4510 1624 4512 1628
rect 4516 1624 4518 1628
rect 4510 1622 4518 1624
rect 4534 1628 4542 1630
rect 4534 1624 4536 1628
rect 4540 1624 4542 1628
rect 4534 1622 4542 1624
rect 4558 1628 4566 1630
rect 4558 1624 4560 1628
rect 4564 1624 4566 1628
rect 4558 1622 4566 1624
rect 4582 1628 4590 1630
rect 4582 1624 4584 1628
rect 4588 1624 4590 1628
rect 4582 1622 4590 1624
rect 4606 1628 4614 1630
rect 4606 1624 4608 1628
rect 4612 1624 4614 1628
rect 4606 1622 4614 1624
rect 4630 1628 4638 1630
rect 4630 1624 4632 1628
rect 4636 1624 4638 1628
rect 4630 1622 4638 1624
rect 4654 1628 4662 1630
rect 4654 1624 4656 1628
rect 4660 1624 4662 1628
rect 4654 1622 4662 1624
rect 4678 1628 4686 1630
rect 4678 1624 4680 1628
rect 4684 1624 4686 1628
rect 4678 1622 4686 1624
rect 4702 1628 4710 1630
rect 4702 1624 4704 1628
rect 4708 1624 4710 1628
rect 4702 1622 4710 1624
rect 4726 1628 4734 1630
rect 4726 1624 4728 1628
rect 4732 1624 4734 1628
rect 4726 1622 4734 1624
rect 4750 1628 4758 1630
rect 4750 1624 4752 1628
rect 4756 1624 4758 1628
rect 4750 1622 4758 1624
rect 4774 1628 4782 1630
rect 4774 1624 4776 1628
rect 4780 1624 4782 1628
rect 4774 1622 4782 1624
rect 4798 1622 4800 1630
rect 5710 1628 5718 1630
rect 5710 1624 5712 1628
rect 5716 1624 5718 1628
rect 5710 1622 5718 1624
rect 5734 1628 5742 1630
rect 5734 1624 5736 1628
rect 5740 1624 5742 1628
rect 5734 1622 5742 1624
rect 5758 1628 5766 1630
rect 5758 1624 5760 1628
rect 5764 1624 5766 1628
rect 5758 1622 5766 1624
rect 5782 1628 5790 1630
rect 5782 1624 5784 1628
rect 5788 1624 5790 1628
rect 5782 1622 5790 1624
rect 5806 1628 5814 1630
rect 5806 1624 5808 1628
rect 5812 1624 5814 1628
rect 5806 1622 5814 1624
rect 5830 1628 5838 1630
rect 5830 1624 5832 1628
rect 5836 1624 5838 1628
rect 5830 1622 5838 1624
rect 5854 1628 5862 1630
rect 5854 1624 5856 1628
rect 5860 1624 5862 1628
rect 5854 1622 5862 1624
rect 5878 1628 5886 1630
rect 5878 1624 5880 1628
rect 5884 1624 5886 1628
rect 5878 1622 5886 1624
rect 5902 1628 5910 1630
rect 5902 1624 5904 1628
rect 5908 1624 5910 1628
rect 5902 1622 5910 1624
rect 5926 1628 5934 1630
rect 5926 1624 5928 1628
rect 5932 1624 5934 1628
rect 5926 1622 5934 1624
rect 5950 1628 5958 1630
rect 5950 1624 5952 1628
rect 5956 1624 5958 1628
rect 5950 1622 5958 1624
rect 5974 1628 5982 1630
rect 5974 1624 5976 1628
rect 5980 1624 5982 1628
rect 5974 1622 5982 1624
rect 5998 1628 6006 1630
rect 5998 1624 6000 1628
rect 6004 1624 6006 1628
rect 5998 1622 6006 1624
rect 6022 1628 6030 1630
rect 6022 1624 6024 1628
rect 6028 1624 6030 1628
rect 6022 1622 6030 1624
rect 6046 1628 6054 1630
rect 6046 1624 6048 1628
rect 6052 1624 6054 1628
rect 6046 1622 6054 1624
rect 6070 1628 6078 1630
rect 6070 1624 6072 1628
rect 6076 1624 6078 1628
rect 6070 1622 6078 1624
rect 6094 1628 6102 1630
rect 6094 1624 6096 1628
rect 6100 1624 6102 1628
rect 6094 1622 6102 1624
rect 6310 1628 6318 1630
rect 6310 1624 6312 1628
rect 6316 1624 6318 1628
rect 6310 1622 6318 1624
rect 6334 1628 6342 1630
rect 6334 1624 6336 1628
rect 6340 1624 6342 1628
rect 6334 1622 6342 1624
rect 6358 1628 6366 1630
rect 6358 1624 6360 1628
rect 6364 1624 6366 1628
rect 6358 1622 6366 1624
rect 6382 1628 6390 1630
rect 6382 1624 6384 1628
rect 6388 1624 6390 1628
rect 6382 1622 6390 1624
rect 6406 1628 6414 1630
rect 6406 1624 6408 1628
rect 6412 1624 6414 1628
rect 6406 1622 6414 1624
rect 6430 1628 6438 1630
rect 6430 1624 6432 1628
rect 6436 1624 6438 1628
rect 6430 1622 6438 1624
rect 6454 1628 6462 1630
rect 6454 1624 6456 1628
rect 6460 1624 6462 1628
rect 6454 1622 6462 1624
rect 6478 1628 6486 1630
rect 6478 1624 6480 1628
rect 6484 1624 6486 1628
rect 6478 1622 6486 1624
rect 6502 1628 6510 1630
rect 6502 1624 6504 1628
rect 6508 1624 6510 1628
rect 6502 1622 6510 1624
rect 6526 1628 6534 1630
rect 6526 1624 6528 1628
rect 6532 1624 6534 1628
rect 6526 1622 6534 1624
rect 6550 1628 6558 1630
rect 6550 1624 6552 1628
rect 6556 1624 6558 1628
rect 6550 1622 6558 1624
rect 6574 1628 6582 1630
rect 6574 1624 6576 1628
rect 6580 1624 6582 1628
rect 6574 1622 6582 1624
rect 6598 1628 6606 1630
rect 6598 1624 6600 1628
rect 6604 1624 6606 1628
rect 6598 1622 6606 1624
rect 6622 1628 6630 1630
rect 6622 1624 6624 1628
rect 6628 1624 6630 1628
rect 6622 1622 6630 1624
rect 6646 1628 6654 1630
rect 6646 1624 6648 1628
rect 6652 1624 6654 1628
rect 6646 1622 6654 1624
rect 6670 1628 6678 1630
rect 6670 1624 6672 1628
rect 6676 1624 6678 1628
rect 6670 1622 6678 1624
rect 6694 1628 6702 1630
rect 6694 1624 6696 1628
rect 6700 1624 6702 1628
rect 6694 1622 6702 1624
rect 6910 1628 6918 1630
rect 6910 1624 6912 1628
rect 6916 1624 6918 1628
rect 6910 1622 6918 1624
rect 6934 1628 6942 1630
rect 6934 1624 6936 1628
rect 6940 1624 6942 1628
rect 6934 1622 6942 1624
rect 6958 1628 6966 1630
rect 6958 1624 6960 1628
rect 6964 1624 6966 1628
rect 6958 1622 6966 1624
rect 6982 1628 6990 1630
rect 6982 1624 6984 1628
rect 6988 1624 6990 1628
rect 6982 1622 6990 1624
rect 7006 1628 7014 1630
rect 7006 1624 7008 1628
rect 7012 1624 7014 1628
rect 7006 1622 7014 1624
rect 7030 1628 7038 1630
rect 7030 1624 7032 1628
rect 7036 1624 7038 1628
rect 7030 1622 7038 1624
rect 7054 1628 7062 1630
rect 7054 1624 7056 1628
rect 7060 1624 7062 1628
rect 7054 1622 7062 1624
rect 7078 1628 7086 1630
rect 7078 1624 7080 1628
rect 7084 1624 7086 1628
rect 7078 1622 7086 1624
rect 7102 1628 7110 1630
rect 7102 1624 7104 1628
rect 7108 1624 7110 1628
rect 7102 1622 7110 1624
rect 7126 1628 7134 1630
rect 7126 1624 7128 1628
rect 7132 1624 7134 1628
rect 7126 1622 7134 1624
rect 7150 1628 7158 1630
rect 7150 1624 7152 1628
rect 7156 1624 7158 1628
rect 7150 1622 7158 1624
rect 7174 1628 7182 1630
rect 7174 1624 7176 1628
rect 7180 1624 7182 1628
rect 7174 1622 7182 1624
rect 7198 1622 7200 1630
rect 2410 1616 2418 1618
rect 2410 1612 2412 1616
rect 2416 1612 2418 1616
rect 2410 1610 2418 1612
rect 2434 1616 2442 1618
rect 2434 1612 2436 1616
rect 2440 1612 2442 1616
rect 2434 1610 2442 1612
rect 2458 1616 2466 1618
rect 2458 1612 2460 1616
rect 2464 1612 2466 1616
rect 2458 1610 2466 1612
rect 2482 1616 2490 1618
rect 2482 1612 2484 1616
rect 2488 1612 2490 1616
rect 2482 1610 2490 1612
rect 2698 1616 2706 1618
rect 2698 1612 2700 1616
rect 2704 1612 2706 1616
rect 2698 1610 2706 1612
rect 2722 1616 2730 1618
rect 2722 1612 2724 1616
rect 2728 1612 2730 1616
rect 2722 1610 2730 1612
rect 2746 1616 2754 1618
rect 2746 1612 2748 1616
rect 2752 1612 2754 1616
rect 2746 1610 2754 1612
rect 2770 1616 2778 1618
rect 2770 1612 2772 1616
rect 2776 1612 2778 1616
rect 2770 1610 2778 1612
rect 2794 1616 2802 1618
rect 2794 1612 2796 1616
rect 2800 1612 2802 1616
rect 2794 1610 2802 1612
rect 2818 1616 2826 1618
rect 2818 1612 2820 1616
rect 2824 1612 2826 1616
rect 2818 1610 2826 1612
rect 2842 1616 2850 1618
rect 2842 1612 2844 1616
rect 2848 1612 2850 1616
rect 2842 1610 2850 1612
rect 2866 1616 2874 1618
rect 2866 1612 2868 1616
rect 2872 1612 2874 1616
rect 2866 1610 2874 1612
rect 2890 1616 2898 1618
rect 2890 1612 2892 1616
rect 2896 1612 2898 1616
rect 2890 1610 2898 1612
rect 2914 1616 2922 1618
rect 2914 1612 2916 1616
rect 2920 1612 2922 1616
rect 2914 1610 2922 1612
rect 2938 1616 2946 1618
rect 2938 1612 2940 1616
rect 2944 1612 2946 1616
rect 2938 1610 2946 1612
rect 2962 1616 2970 1618
rect 2962 1612 2964 1616
rect 2968 1612 2970 1616
rect 2962 1610 2970 1612
rect 2986 1616 2994 1618
rect 2986 1612 2988 1616
rect 2992 1612 2994 1616
rect 2986 1610 2994 1612
rect 3010 1616 3018 1618
rect 3010 1612 3012 1616
rect 3016 1612 3018 1616
rect 3010 1610 3018 1612
rect 3034 1616 3042 1618
rect 3034 1612 3036 1616
rect 3040 1612 3042 1616
rect 3034 1610 3042 1612
rect 3058 1616 3066 1618
rect 3058 1612 3060 1616
rect 3064 1612 3066 1616
rect 3058 1610 3066 1612
rect 3082 1616 3090 1618
rect 3082 1612 3084 1616
rect 3088 1612 3090 1616
rect 3082 1610 3090 1612
rect 3298 1616 3306 1618
rect 3298 1612 3300 1616
rect 3304 1612 3306 1616
rect 3298 1610 3306 1612
rect 3322 1616 3330 1618
rect 3322 1612 3324 1616
rect 3328 1612 3330 1616
rect 3322 1610 3330 1612
rect 3346 1616 3354 1618
rect 3346 1612 3348 1616
rect 3352 1612 3354 1616
rect 3346 1610 3354 1612
rect 3370 1616 3378 1618
rect 3370 1612 3372 1616
rect 3376 1612 3378 1616
rect 3370 1610 3378 1612
rect 3394 1616 3402 1618
rect 3394 1612 3396 1616
rect 3400 1612 3402 1616
rect 3394 1610 3402 1612
rect 3418 1616 3426 1618
rect 3418 1612 3420 1616
rect 3424 1612 3426 1616
rect 3418 1610 3426 1612
rect 3442 1616 3450 1618
rect 3442 1612 3444 1616
rect 3448 1612 3450 1616
rect 3442 1610 3450 1612
rect 3466 1616 3474 1618
rect 3466 1612 3468 1616
rect 3472 1612 3474 1616
rect 3466 1610 3474 1612
rect 3490 1616 3498 1618
rect 3490 1612 3492 1616
rect 3496 1612 3498 1616
rect 3490 1610 3498 1612
rect 3514 1616 3522 1618
rect 3514 1612 3516 1616
rect 3520 1612 3522 1616
rect 3514 1610 3522 1612
rect 3538 1616 3546 1618
rect 3538 1612 3540 1616
rect 3544 1612 3546 1616
rect 3538 1610 3546 1612
rect 3562 1616 3570 1618
rect 3562 1612 3564 1616
rect 3568 1612 3570 1616
rect 3562 1610 3570 1612
rect 3586 1616 3594 1618
rect 3586 1612 3588 1616
rect 3592 1612 3594 1616
rect 3586 1610 3594 1612
rect 3610 1616 3618 1618
rect 3610 1612 3612 1616
rect 3616 1612 3618 1616
rect 3610 1610 3618 1612
rect 3634 1616 3642 1618
rect 3634 1612 3636 1616
rect 3640 1612 3642 1616
rect 3634 1610 3642 1612
rect 3658 1616 3666 1618
rect 3658 1612 3660 1616
rect 3664 1612 3666 1616
rect 3658 1610 3666 1612
rect 3682 1616 3690 1618
rect 3682 1612 3684 1616
rect 3688 1612 3690 1616
rect 3682 1610 3690 1612
rect 3898 1616 3906 1618
rect 3898 1612 3900 1616
rect 3904 1612 3906 1616
rect 3898 1610 3906 1612
rect 3922 1616 3930 1618
rect 3922 1612 3924 1616
rect 3928 1612 3930 1616
rect 3922 1610 3930 1612
rect 3946 1616 3954 1618
rect 3946 1612 3948 1616
rect 3952 1612 3954 1616
rect 3946 1610 3954 1612
rect 3970 1616 3978 1618
rect 3970 1612 3972 1616
rect 3976 1612 3978 1616
rect 3970 1610 3978 1612
rect 3994 1616 4002 1618
rect 3994 1612 3996 1616
rect 4000 1612 4002 1616
rect 3994 1610 4002 1612
rect 4018 1616 4026 1618
rect 4018 1612 4020 1616
rect 4024 1612 4026 1616
rect 4018 1610 4026 1612
rect 4042 1616 4050 1618
rect 4042 1612 4044 1616
rect 4048 1612 4050 1616
rect 4042 1610 4050 1612
rect 4066 1616 4074 1618
rect 4066 1612 4068 1616
rect 4072 1612 4074 1616
rect 4066 1610 4074 1612
rect 4090 1616 4098 1618
rect 4090 1612 4092 1616
rect 4096 1612 4098 1616
rect 4090 1610 4098 1612
rect 4114 1616 4122 1618
rect 4114 1612 4116 1616
rect 4120 1612 4122 1616
rect 4114 1610 4122 1612
rect 4138 1616 4146 1618
rect 4138 1612 4140 1616
rect 4144 1612 4146 1616
rect 4138 1610 4146 1612
rect 4162 1616 4170 1618
rect 4162 1612 4164 1616
rect 4168 1612 4170 1616
rect 4162 1610 4170 1612
rect 4186 1616 4194 1618
rect 4186 1612 4188 1616
rect 4192 1612 4194 1616
rect 4186 1610 4194 1612
rect 4210 1616 4218 1618
rect 4210 1612 4212 1616
rect 4216 1612 4218 1616
rect 4210 1610 4218 1612
rect 4234 1616 4242 1618
rect 4234 1612 4236 1616
rect 4240 1612 4242 1616
rect 4234 1610 4242 1612
rect 4258 1616 4266 1618
rect 4258 1612 4260 1616
rect 4264 1612 4266 1616
rect 4258 1610 4266 1612
rect 4282 1616 4290 1618
rect 4282 1612 4284 1616
rect 4288 1612 4290 1616
rect 4282 1610 4290 1612
rect 4498 1616 4506 1618
rect 4498 1612 4500 1616
rect 4504 1612 4506 1616
rect 4498 1610 4506 1612
rect 4522 1616 4530 1618
rect 4522 1612 4524 1616
rect 4528 1612 4530 1616
rect 4522 1610 4530 1612
rect 4546 1616 4554 1618
rect 4546 1612 4548 1616
rect 4552 1612 4554 1616
rect 4546 1610 4554 1612
rect 4570 1616 4578 1618
rect 4570 1612 4572 1616
rect 4576 1612 4578 1616
rect 4570 1610 4578 1612
rect 4594 1616 4602 1618
rect 4594 1612 4596 1616
rect 4600 1612 4602 1616
rect 4594 1610 4602 1612
rect 4618 1616 4626 1618
rect 4618 1612 4620 1616
rect 4624 1612 4626 1616
rect 4618 1610 4626 1612
rect 4642 1616 4650 1618
rect 4642 1612 4644 1616
rect 4648 1612 4650 1616
rect 4642 1610 4650 1612
rect 4666 1616 4674 1618
rect 4666 1612 4668 1616
rect 4672 1612 4674 1616
rect 4666 1610 4674 1612
rect 4690 1616 4698 1618
rect 4690 1612 4692 1616
rect 4696 1612 4698 1616
rect 4690 1610 4698 1612
rect 4714 1616 4722 1618
rect 4714 1612 4716 1616
rect 4720 1612 4722 1616
rect 4714 1610 4722 1612
rect 4738 1616 4746 1618
rect 4738 1612 4740 1616
rect 4744 1612 4746 1616
rect 4738 1610 4746 1612
rect 4762 1616 4770 1618
rect 4762 1612 4764 1616
rect 4768 1612 4770 1616
rect 4762 1610 4770 1612
rect 4786 1616 4794 1618
rect 4786 1612 4788 1616
rect 4792 1612 4794 1616
rect 4786 1610 4794 1612
rect 5698 1616 5706 1618
rect 5698 1612 5700 1616
rect 5704 1612 5706 1616
rect 5698 1610 5706 1612
rect 5722 1616 5730 1618
rect 5722 1612 5724 1616
rect 5728 1612 5730 1616
rect 5722 1610 5730 1612
rect 5746 1616 5754 1618
rect 5746 1612 5748 1616
rect 5752 1612 5754 1616
rect 5746 1610 5754 1612
rect 5770 1616 5778 1618
rect 5770 1612 5772 1616
rect 5776 1612 5778 1616
rect 5770 1610 5778 1612
rect 5794 1616 5802 1618
rect 5794 1612 5796 1616
rect 5800 1612 5802 1616
rect 5794 1610 5802 1612
rect 5818 1616 5826 1618
rect 5818 1612 5820 1616
rect 5824 1612 5826 1616
rect 5818 1610 5826 1612
rect 5842 1616 5850 1618
rect 5842 1612 5844 1616
rect 5848 1612 5850 1616
rect 5842 1610 5850 1612
rect 5866 1616 5874 1618
rect 5866 1612 5868 1616
rect 5872 1612 5874 1616
rect 5866 1610 5874 1612
rect 5890 1616 5898 1618
rect 5890 1612 5892 1616
rect 5896 1612 5898 1616
rect 5890 1610 5898 1612
rect 5914 1616 5922 1618
rect 5914 1612 5916 1616
rect 5920 1612 5922 1616
rect 5914 1610 5922 1612
rect 5938 1616 5946 1618
rect 5938 1612 5940 1616
rect 5944 1612 5946 1616
rect 5938 1610 5946 1612
rect 5962 1616 5970 1618
rect 5962 1612 5964 1616
rect 5968 1612 5970 1616
rect 5962 1610 5970 1612
rect 5986 1616 5994 1618
rect 5986 1612 5988 1616
rect 5992 1612 5994 1616
rect 5986 1610 5994 1612
rect 6010 1616 6018 1618
rect 6010 1612 6012 1616
rect 6016 1612 6018 1616
rect 6010 1610 6018 1612
rect 6034 1616 6042 1618
rect 6034 1612 6036 1616
rect 6040 1612 6042 1616
rect 6034 1610 6042 1612
rect 6058 1616 6066 1618
rect 6058 1612 6060 1616
rect 6064 1612 6066 1616
rect 6058 1610 6066 1612
rect 6082 1616 6090 1618
rect 6082 1612 6084 1616
rect 6088 1612 6090 1616
rect 6082 1610 6090 1612
rect 6298 1616 6306 1618
rect 6298 1612 6300 1616
rect 6304 1612 6306 1616
rect 6298 1610 6306 1612
rect 6322 1616 6330 1618
rect 6322 1612 6324 1616
rect 6328 1612 6330 1616
rect 6322 1610 6330 1612
rect 6346 1616 6354 1618
rect 6346 1612 6348 1616
rect 6352 1612 6354 1616
rect 6346 1610 6354 1612
rect 6370 1616 6378 1618
rect 6370 1612 6372 1616
rect 6376 1612 6378 1616
rect 6370 1610 6378 1612
rect 6394 1616 6402 1618
rect 6394 1612 6396 1616
rect 6400 1612 6402 1616
rect 6394 1610 6402 1612
rect 6418 1616 6426 1618
rect 6418 1612 6420 1616
rect 6424 1612 6426 1616
rect 6418 1610 6426 1612
rect 6442 1616 6450 1618
rect 6442 1612 6444 1616
rect 6448 1612 6450 1616
rect 6442 1610 6450 1612
rect 6466 1616 6474 1618
rect 6466 1612 6468 1616
rect 6472 1612 6474 1616
rect 6466 1610 6474 1612
rect 6490 1616 6498 1618
rect 6490 1612 6492 1616
rect 6496 1612 6498 1616
rect 6490 1610 6498 1612
rect 6514 1616 6522 1618
rect 6514 1612 6516 1616
rect 6520 1612 6522 1616
rect 6514 1610 6522 1612
rect 6538 1616 6546 1618
rect 6538 1612 6540 1616
rect 6544 1612 6546 1616
rect 6538 1610 6546 1612
rect 6562 1616 6570 1618
rect 6562 1612 6564 1616
rect 6568 1612 6570 1616
rect 6562 1610 6570 1612
rect 6586 1616 6594 1618
rect 6586 1612 6588 1616
rect 6592 1612 6594 1616
rect 6586 1610 6594 1612
rect 6610 1616 6618 1618
rect 6610 1612 6612 1616
rect 6616 1612 6618 1616
rect 6610 1610 6618 1612
rect 6634 1616 6642 1618
rect 6634 1612 6636 1616
rect 6640 1612 6642 1616
rect 6634 1610 6642 1612
rect 6658 1616 6666 1618
rect 6658 1612 6660 1616
rect 6664 1612 6666 1616
rect 6658 1610 6666 1612
rect 6682 1616 6690 1618
rect 6682 1612 6684 1616
rect 6688 1612 6690 1616
rect 6682 1610 6690 1612
rect 6898 1616 6906 1618
rect 6898 1612 6900 1616
rect 6904 1612 6906 1616
rect 6898 1610 6906 1612
rect 6922 1616 6930 1618
rect 6922 1612 6924 1616
rect 6928 1612 6930 1616
rect 6922 1610 6930 1612
rect 6946 1616 6954 1618
rect 6946 1612 6948 1616
rect 6952 1612 6954 1616
rect 6946 1610 6954 1612
rect 6970 1616 6978 1618
rect 6970 1612 6972 1616
rect 6976 1612 6978 1616
rect 6970 1610 6978 1612
rect 6994 1616 7002 1618
rect 6994 1612 6996 1616
rect 7000 1612 7002 1616
rect 6994 1610 7002 1612
rect 7018 1616 7026 1618
rect 7018 1612 7020 1616
rect 7024 1612 7026 1616
rect 7018 1610 7026 1612
rect 7042 1616 7050 1618
rect 7042 1612 7044 1616
rect 7048 1612 7050 1616
rect 7042 1610 7050 1612
rect 7066 1616 7074 1618
rect 7066 1612 7068 1616
rect 7072 1612 7074 1616
rect 7066 1610 7074 1612
rect 7090 1616 7098 1618
rect 7090 1612 7092 1616
rect 7096 1612 7098 1616
rect 7090 1610 7098 1612
rect 7114 1616 7122 1618
rect 7114 1612 7116 1616
rect 7120 1612 7122 1616
rect 7114 1610 7122 1612
rect 7138 1616 7146 1618
rect 7138 1612 7140 1616
rect 7144 1612 7146 1616
rect 7138 1610 7146 1612
rect 7162 1616 7170 1618
rect 7162 1612 7164 1616
rect 7168 1612 7170 1616
rect 7162 1610 7170 1612
rect 7186 1616 7194 1618
rect 7186 1612 7188 1616
rect 7192 1612 7194 1616
rect 7186 1610 7194 1612
rect 2400 1604 2406 1606
rect 2404 1600 2406 1604
rect 2110 1598 2118 1600
rect 2134 1598 2142 1600
rect 2158 1598 2166 1600
rect 2182 1598 2190 1600
rect 2206 1598 2214 1600
rect 2230 1598 2238 1600
rect 2254 1598 2262 1600
rect 2278 1598 2286 1600
rect 2302 1598 2310 1600
rect 2326 1598 2334 1600
rect 2350 1598 2358 1600
rect 2374 1598 2382 1600
rect 2398 1598 2406 1600
rect 2422 1604 2430 1606
rect 2422 1600 2424 1604
rect 2428 1600 2430 1604
rect 2422 1598 2430 1600
rect 2446 1604 2454 1606
rect 2446 1600 2448 1604
rect 2452 1600 2454 1604
rect 2446 1598 2454 1600
rect 2470 1604 2478 1606
rect 2470 1600 2472 1604
rect 2476 1600 2478 1604
rect 2470 1598 2478 1600
rect 2494 1604 2502 1606
rect 2494 1600 2496 1604
rect 2500 1600 2502 1604
rect 2494 1598 2502 1600
rect 2710 1604 2718 1606
rect 2710 1600 2712 1604
rect 2716 1600 2718 1604
rect 2710 1598 2718 1600
rect 2734 1604 2742 1606
rect 2734 1600 2736 1604
rect 2740 1600 2742 1604
rect 2734 1598 2742 1600
rect 2758 1604 2766 1606
rect 2758 1600 2760 1604
rect 2764 1600 2766 1604
rect 2758 1598 2766 1600
rect 2782 1604 2790 1606
rect 2782 1600 2784 1604
rect 2788 1600 2790 1604
rect 2782 1598 2790 1600
rect 2806 1604 2814 1606
rect 2806 1600 2808 1604
rect 2812 1600 2814 1604
rect 2806 1598 2814 1600
rect 2830 1604 2838 1606
rect 2830 1600 2832 1604
rect 2836 1600 2838 1604
rect 2830 1598 2838 1600
rect 2854 1604 2862 1606
rect 2854 1600 2856 1604
rect 2860 1600 2862 1604
rect 2854 1598 2862 1600
rect 2878 1604 2886 1606
rect 2878 1600 2880 1604
rect 2884 1600 2886 1604
rect 2878 1598 2886 1600
rect 2902 1604 2910 1606
rect 2902 1600 2904 1604
rect 2908 1600 2910 1604
rect 2902 1598 2910 1600
rect 2926 1604 2934 1606
rect 2926 1600 2928 1604
rect 2932 1600 2934 1604
rect 2926 1598 2934 1600
rect 2950 1604 2958 1606
rect 2950 1600 2952 1604
rect 2956 1600 2958 1604
rect 2950 1598 2958 1600
rect 2974 1604 2982 1606
rect 2974 1600 2976 1604
rect 2980 1600 2982 1604
rect 2974 1598 2982 1600
rect 2998 1604 3006 1606
rect 2998 1600 3000 1604
rect 3004 1600 3006 1604
rect 2998 1598 3006 1600
rect 3022 1604 3030 1606
rect 3022 1600 3024 1604
rect 3028 1600 3030 1604
rect 3022 1598 3030 1600
rect 3046 1604 3054 1606
rect 3046 1600 3048 1604
rect 3052 1600 3054 1604
rect 3046 1598 3054 1600
rect 3070 1604 3078 1606
rect 3070 1600 3072 1604
rect 3076 1600 3078 1604
rect 3070 1598 3078 1600
rect 3094 1604 3102 1606
rect 3094 1600 3096 1604
rect 3100 1600 3102 1604
rect 3094 1598 3102 1600
rect 3310 1604 3318 1606
rect 3310 1600 3312 1604
rect 3316 1600 3318 1604
rect 3310 1598 3318 1600
rect 3334 1604 3342 1606
rect 3334 1600 3336 1604
rect 3340 1600 3342 1604
rect 3334 1598 3342 1600
rect 3358 1604 3366 1606
rect 3358 1600 3360 1604
rect 3364 1600 3366 1604
rect 3358 1598 3366 1600
rect 3382 1604 3390 1606
rect 3382 1600 3384 1604
rect 3388 1600 3390 1604
rect 3382 1598 3390 1600
rect 3406 1604 3414 1606
rect 3406 1600 3408 1604
rect 3412 1600 3414 1604
rect 3406 1598 3414 1600
rect 3430 1604 3438 1606
rect 3430 1600 3432 1604
rect 3436 1600 3438 1604
rect 3430 1598 3438 1600
rect 3454 1604 3462 1606
rect 3454 1600 3456 1604
rect 3460 1600 3462 1604
rect 3454 1598 3462 1600
rect 3478 1604 3486 1606
rect 3478 1600 3480 1604
rect 3484 1600 3486 1604
rect 3478 1598 3486 1600
rect 3502 1604 3510 1606
rect 3502 1600 3504 1604
rect 3508 1600 3510 1604
rect 3502 1598 3510 1600
rect 3526 1604 3534 1606
rect 3526 1600 3528 1604
rect 3532 1600 3534 1604
rect 3526 1598 3534 1600
rect 3550 1604 3558 1606
rect 3550 1600 3552 1604
rect 3556 1600 3558 1604
rect 3550 1598 3558 1600
rect 3574 1604 3582 1606
rect 3574 1600 3576 1604
rect 3580 1600 3582 1604
rect 3574 1598 3582 1600
rect 3598 1604 3606 1606
rect 3598 1600 3600 1604
rect 3604 1600 3606 1604
rect 3598 1598 3606 1600
rect 3622 1604 3630 1606
rect 3622 1600 3624 1604
rect 3628 1600 3630 1604
rect 3622 1598 3630 1600
rect 3646 1604 3654 1606
rect 3646 1600 3648 1604
rect 3652 1600 3654 1604
rect 3646 1598 3654 1600
rect 3670 1604 3678 1606
rect 3670 1600 3672 1604
rect 3676 1600 3678 1604
rect 3670 1598 3678 1600
rect 3694 1604 3702 1606
rect 3694 1600 3696 1604
rect 3700 1600 3702 1604
rect 3694 1598 3702 1600
rect 3910 1604 3918 1606
rect 3910 1600 3912 1604
rect 3916 1600 3918 1604
rect 3910 1598 3918 1600
rect 3934 1604 3942 1606
rect 3934 1600 3936 1604
rect 3940 1600 3942 1604
rect 3934 1598 3942 1600
rect 3958 1604 3966 1606
rect 3958 1600 3960 1604
rect 3964 1600 3966 1604
rect 3958 1598 3966 1600
rect 3982 1604 3990 1606
rect 3982 1600 3984 1604
rect 3988 1600 3990 1604
rect 3982 1598 3990 1600
rect 4006 1604 4014 1606
rect 4006 1600 4008 1604
rect 4012 1600 4014 1604
rect 4006 1598 4014 1600
rect 4030 1604 4038 1606
rect 4030 1600 4032 1604
rect 4036 1600 4038 1604
rect 4030 1598 4038 1600
rect 4054 1604 4062 1606
rect 4054 1600 4056 1604
rect 4060 1600 4062 1604
rect 4054 1598 4062 1600
rect 4078 1604 4086 1606
rect 4078 1600 4080 1604
rect 4084 1600 4086 1604
rect 4078 1598 4086 1600
rect 4102 1604 4110 1606
rect 4102 1600 4104 1604
rect 4108 1600 4110 1604
rect 4102 1598 4110 1600
rect 4126 1604 4134 1606
rect 4126 1600 4128 1604
rect 4132 1600 4134 1604
rect 4126 1598 4134 1600
rect 4150 1604 4158 1606
rect 4150 1600 4152 1604
rect 4156 1600 4158 1604
rect 4150 1598 4158 1600
rect 4174 1604 4182 1606
rect 4174 1600 4176 1604
rect 4180 1600 4182 1604
rect 4174 1598 4182 1600
rect 4198 1604 4206 1606
rect 4198 1600 4200 1604
rect 4204 1600 4206 1604
rect 4198 1598 4206 1600
rect 4222 1604 4230 1606
rect 4222 1600 4224 1604
rect 4228 1600 4230 1604
rect 4222 1598 4230 1600
rect 4246 1604 4254 1606
rect 4246 1600 4248 1604
rect 4252 1600 4254 1604
rect 4246 1598 4254 1600
rect 4270 1604 4278 1606
rect 4270 1600 4272 1604
rect 4276 1600 4278 1604
rect 4270 1598 4278 1600
rect 4294 1604 4302 1606
rect 4294 1600 4296 1604
rect 4300 1600 4302 1604
rect 4294 1598 4302 1600
rect 4510 1604 4518 1606
rect 4510 1600 4512 1604
rect 4516 1600 4518 1604
rect 4510 1598 4518 1600
rect 4534 1604 4542 1606
rect 4534 1600 4536 1604
rect 4540 1600 4542 1604
rect 4534 1598 4542 1600
rect 4558 1604 4566 1606
rect 4558 1600 4560 1604
rect 4564 1600 4566 1604
rect 4558 1598 4566 1600
rect 4582 1604 4590 1606
rect 4582 1600 4584 1604
rect 4588 1600 4590 1604
rect 4582 1598 4590 1600
rect 4606 1604 4614 1606
rect 4606 1600 4608 1604
rect 4612 1600 4614 1604
rect 4606 1598 4614 1600
rect 4630 1604 4638 1606
rect 4630 1600 4632 1604
rect 4636 1600 4638 1604
rect 4630 1598 4638 1600
rect 4654 1604 4662 1606
rect 4654 1600 4656 1604
rect 4660 1600 4662 1604
rect 4654 1598 4662 1600
rect 4678 1604 4686 1606
rect 4678 1600 4680 1604
rect 4684 1600 4686 1604
rect 4678 1598 4686 1600
rect 4702 1604 4710 1606
rect 4702 1600 4704 1604
rect 4708 1600 4710 1604
rect 4702 1598 4710 1600
rect 4726 1604 4734 1606
rect 4726 1600 4728 1604
rect 4732 1600 4734 1604
rect 4726 1598 4734 1600
rect 4750 1604 4758 1606
rect 4750 1600 4752 1604
rect 4756 1600 4758 1604
rect 4750 1598 4758 1600
rect 4774 1604 4782 1606
rect 4774 1600 4776 1604
rect 4780 1600 4782 1604
rect 4774 1598 4782 1600
rect 4798 1600 4800 1606
rect 5710 1604 5718 1606
rect 5710 1600 5712 1604
rect 5716 1600 5718 1604
rect 4798 1598 4806 1600
rect 4822 1598 4830 1600
rect 4846 1598 4854 1600
rect 4870 1598 4878 1600
rect 4894 1598 4902 1600
rect 5710 1598 5718 1600
rect 5734 1604 5742 1606
rect 5734 1600 5736 1604
rect 5740 1600 5742 1604
rect 5734 1598 5742 1600
rect 5758 1604 5766 1606
rect 5758 1600 5760 1604
rect 5764 1600 5766 1604
rect 5758 1598 5766 1600
rect 5782 1604 5790 1606
rect 5782 1600 5784 1604
rect 5788 1600 5790 1604
rect 5782 1598 5790 1600
rect 5806 1604 5814 1606
rect 5806 1600 5808 1604
rect 5812 1600 5814 1604
rect 5806 1598 5814 1600
rect 5830 1604 5838 1606
rect 5830 1600 5832 1604
rect 5836 1600 5838 1604
rect 5830 1598 5838 1600
rect 5854 1604 5862 1606
rect 5854 1600 5856 1604
rect 5860 1600 5862 1604
rect 5854 1598 5862 1600
rect 5878 1604 5886 1606
rect 5878 1600 5880 1604
rect 5884 1600 5886 1604
rect 5878 1598 5886 1600
rect 5902 1604 5910 1606
rect 5902 1600 5904 1604
rect 5908 1600 5910 1604
rect 5902 1598 5910 1600
rect 5926 1604 5934 1606
rect 5926 1600 5928 1604
rect 5932 1600 5934 1604
rect 5926 1598 5934 1600
rect 5950 1604 5958 1606
rect 5950 1600 5952 1604
rect 5956 1600 5958 1604
rect 5950 1598 5958 1600
rect 5974 1604 5982 1606
rect 5974 1600 5976 1604
rect 5980 1600 5982 1604
rect 5974 1598 5982 1600
rect 5998 1604 6006 1606
rect 5998 1600 6000 1604
rect 6004 1600 6006 1604
rect 5998 1598 6006 1600
rect 6022 1604 6030 1606
rect 6022 1600 6024 1604
rect 6028 1600 6030 1604
rect 6022 1598 6030 1600
rect 6046 1604 6054 1606
rect 6046 1600 6048 1604
rect 6052 1600 6054 1604
rect 6046 1598 6054 1600
rect 6070 1604 6078 1606
rect 6070 1600 6072 1604
rect 6076 1600 6078 1604
rect 6070 1598 6078 1600
rect 6094 1604 6102 1606
rect 6094 1600 6096 1604
rect 6100 1600 6102 1604
rect 6094 1598 6102 1600
rect 6310 1604 6318 1606
rect 6310 1600 6312 1604
rect 6316 1600 6318 1604
rect 6310 1598 6318 1600
rect 6334 1604 6342 1606
rect 6334 1600 6336 1604
rect 6340 1600 6342 1604
rect 6334 1598 6342 1600
rect 6358 1604 6366 1606
rect 6358 1600 6360 1604
rect 6364 1600 6366 1604
rect 6358 1598 6366 1600
rect 6382 1604 6390 1606
rect 6382 1600 6384 1604
rect 6388 1600 6390 1604
rect 6382 1598 6390 1600
rect 6406 1604 6414 1606
rect 6406 1600 6408 1604
rect 6412 1600 6414 1604
rect 6406 1598 6414 1600
rect 6430 1604 6438 1606
rect 6430 1600 6432 1604
rect 6436 1600 6438 1604
rect 6430 1598 6438 1600
rect 6454 1604 6462 1606
rect 6454 1600 6456 1604
rect 6460 1600 6462 1604
rect 6454 1598 6462 1600
rect 6478 1604 6486 1606
rect 6478 1600 6480 1604
rect 6484 1600 6486 1604
rect 6478 1598 6486 1600
rect 6502 1604 6510 1606
rect 6502 1600 6504 1604
rect 6508 1600 6510 1604
rect 6502 1598 6510 1600
rect 6526 1604 6534 1606
rect 6526 1600 6528 1604
rect 6532 1600 6534 1604
rect 6526 1598 6534 1600
rect 6550 1604 6558 1606
rect 6550 1600 6552 1604
rect 6556 1600 6558 1604
rect 6550 1598 6558 1600
rect 6574 1604 6582 1606
rect 6574 1600 6576 1604
rect 6580 1600 6582 1604
rect 6574 1598 6582 1600
rect 6598 1604 6606 1606
rect 6598 1600 6600 1604
rect 6604 1600 6606 1604
rect 6598 1598 6606 1600
rect 6622 1604 6630 1606
rect 6622 1600 6624 1604
rect 6628 1600 6630 1604
rect 6622 1598 6630 1600
rect 6646 1604 6654 1606
rect 6646 1600 6648 1604
rect 6652 1600 6654 1604
rect 6646 1598 6654 1600
rect 6670 1604 6678 1606
rect 6670 1600 6672 1604
rect 6676 1600 6678 1604
rect 6670 1598 6678 1600
rect 6694 1604 6702 1606
rect 6694 1600 6696 1604
rect 6700 1600 6702 1604
rect 6694 1598 6702 1600
rect 6910 1604 6918 1606
rect 6910 1600 6912 1604
rect 6916 1600 6918 1604
rect 6910 1598 6918 1600
rect 6934 1604 6942 1606
rect 6934 1600 6936 1604
rect 6940 1600 6942 1604
rect 6934 1598 6942 1600
rect 6958 1604 6966 1606
rect 6958 1600 6960 1604
rect 6964 1600 6966 1604
rect 6958 1598 6966 1600
rect 6982 1604 6990 1606
rect 6982 1600 6984 1604
rect 6988 1600 6990 1604
rect 6982 1598 6990 1600
rect 7006 1604 7014 1606
rect 7006 1600 7008 1604
rect 7012 1600 7014 1604
rect 7006 1598 7014 1600
rect 7030 1604 7038 1606
rect 7030 1600 7032 1604
rect 7036 1600 7038 1604
rect 7030 1598 7038 1600
rect 7054 1604 7062 1606
rect 7054 1600 7056 1604
rect 7060 1600 7062 1604
rect 7054 1598 7062 1600
rect 7078 1604 7086 1606
rect 7078 1600 7080 1604
rect 7084 1600 7086 1604
rect 7078 1598 7086 1600
rect 7102 1604 7110 1606
rect 7102 1600 7104 1604
rect 7108 1600 7110 1604
rect 7102 1598 7110 1600
rect 7126 1604 7134 1606
rect 7126 1600 7128 1604
rect 7132 1600 7134 1604
rect 7126 1598 7134 1600
rect 7150 1604 7158 1606
rect 7150 1600 7152 1604
rect 7156 1600 7158 1604
rect 7150 1598 7158 1600
rect 7174 1604 7182 1606
rect 7174 1600 7176 1604
rect 7180 1600 7182 1604
rect 7174 1598 7182 1600
rect 7198 1598 7200 1606
rect 2098 1592 2106 1594
rect 2098 1588 2100 1592
rect 2104 1588 2106 1592
rect 2098 1586 2106 1588
rect 2122 1592 2130 1594
rect 2122 1588 2124 1592
rect 2128 1588 2130 1592
rect 2122 1586 2130 1588
rect 2146 1592 2154 1594
rect 2146 1588 2148 1592
rect 2152 1588 2154 1592
rect 2146 1586 2154 1588
rect 2170 1592 2178 1594
rect 2170 1588 2172 1592
rect 2176 1588 2178 1592
rect 2170 1586 2178 1588
rect 2194 1592 2202 1594
rect 2194 1588 2196 1592
rect 2200 1588 2202 1592
rect 2194 1586 2202 1588
rect 2218 1592 2226 1594
rect 2218 1588 2220 1592
rect 2224 1588 2226 1592
rect 2218 1586 2226 1588
rect 2242 1592 2250 1594
rect 2242 1588 2244 1592
rect 2248 1588 2250 1592
rect 2242 1586 2250 1588
rect 2266 1592 2274 1594
rect 2266 1588 2268 1592
rect 2272 1588 2274 1592
rect 2266 1586 2274 1588
rect 2290 1592 2298 1594
rect 2290 1588 2292 1592
rect 2296 1588 2298 1592
rect 2290 1586 2298 1588
rect 2314 1592 2322 1594
rect 2314 1588 2316 1592
rect 2320 1588 2322 1592
rect 2314 1586 2322 1588
rect 2338 1592 2346 1594
rect 2338 1588 2340 1592
rect 2344 1588 2346 1592
rect 2338 1586 2346 1588
rect 2362 1592 2370 1594
rect 2362 1588 2364 1592
rect 2368 1588 2370 1592
rect 2362 1586 2370 1588
rect 2386 1592 2394 1594
rect 2386 1588 2388 1592
rect 2392 1588 2394 1592
rect 2386 1586 2394 1588
rect 2410 1592 2418 1594
rect 2410 1588 2412 1592
rect 2416 1588 2418 1592
rect 2410 1586 2418 1588
rect 2434 1592 2442 1594
rect 2434 1588 2436 1592
rect 2440 1588 2442 1592
rect 2434 1586 2442 1588
rect 2458 1592 2466 1594
rect 2458 1588 2460 1592
rect 2464 1588 2466 1592
rect 2458 1586 2466 1588
rect 2482 1592 2490 1594
rect 2482 1588 2484 1592
rect 2488 1588 2490 1592
rect 2482 1586 2490 1588
rect 2698 1592 2706 1594
rect 2698 1588 2700 1592
rect 2704 1588 2706 1592
rect 2698 1586 2706 1588
rect 2722 1592 2730 1594
rect 2722 1588 2724 1592
rect 2728 1588 2730 1592
rect 2722 1586 2730 1588
rect 2746 1592 2754 1594
rect 2746 1588 2748 1592
rect 2752 1588 2754 1592
rect 2746 1586 2754 1588
rect 2770 1592 2778 1594
rect 2770 1588 2772 1592
rect 2776 1588 2778 1592
rect 2770 1586 2778 1588
rect 2794 1592 2802 1594
rect 2794 1588 2796 1592
rect 2800 1588 2802 1592
rect 2794 1586 2802 1588
rect 2818 1592 2826 1594
rect 2818 1588 2820 1592
rect 2824 1588 2826 1592
rect 2818 1586 2826 1588
rect 2842 1592 2850 1594
rect 2842 1588 2844 1592
rect 2848 1588 2850 1592
rect 2842 1586 2850 1588
rect 2866 1592 2874 1594
rect 2866 1588 2868 1592
rect 2872 1588 2874 1592
rect 2866 1586 2874 1588
rect 2890 1592 2898 1594
rect 2890 1588 2892 1592
rect 2896 1588 2898 1592
rect 2890 1586 2898 1588
rect 2914 1592 2922 1594
rect 2914 1588 2916 1592
rect 2920 1588 2922 1592
rect 2914 1586 2922 1588
rect 2938 1592 2946 1594
rect 2938 1588 2940 1592
rect 2944 1588 2946 1592
rect 2938 1586 2946 1588
rect 2962 1592 2970 1594
rect 2962 1588 2964 1592
rect 2968 1588 2970 1592
rect 2962 1586 2970 1588
rect 2986 1592 2994 1594
rect 2986 1588 2988 1592
rect 2992 1588 2994 1592
rect 2986 1586 2994 1588
rect 3010 1592 3018 1594
rect 3010 1588 3012 1592
rect 3016 1588 3018 1592
rect 3010 1586 3018 1588
rect 3034 1592 3042 1594
rect 3034 1588 3036 1592
rect 3040 1588 3042 1592
rect 3034 1586 3042 1588
rect 3058 1592 3066 1594
rect 3058 1588 3060 1592
rect 3064 1588 3066 1592
rect 3058 1586 3066 1588
rect 3082 1592 3090 1594
rect 3082 1588 3084 1592
rect 3088 1588 3090 1592
rect 3082 1586 3090 1588
rect 3298 1592 3306 1594
rect 3298 1588 3300 1592
rect 3304 1588 3306 1592
rect 3298 1586 3306 1588
rect 3322 1592 3330 1594
rect 3322 1588 3324 1592
rect 3328 1588 3330 1592
rect 3322 1586 3330 1588
rect 3346 1592 3354 1594
rect 3346 1588 3348 1592
rect 3352 1588 3354 1592
rect 3346 1586 3354 1588
rect 3370 1592 3378 1594
rect 3370 1588 3372 1592
rect 3376 1588 3378 1592
rect 3370 1586 3378 1588
rect 3394 1592 3402 1594
rect 3394 1588 3396 1592
rect 3400 1588 3402 1592
rect 3394 1586 3402 1588
rect 3418 1592 3426 1594
rect 3418 1588 3420 1592
rect 3424 1588 3426 1592
rect 3418 1586 3426 1588
rect 3442 1592 3450 1594
rect 3442 1588 3444 1592
rect 3448 1588 3450 1592
rect 3442 1586 3450 1588
rect 3466 1592 3474 1594
rect 3466 1588 3468 1592
rect 3472 1588 3474 1592
rect 3466 1586 3474 1588
rect 3490 1592 3498 1594
rect 3490 1588 3492 1592
rect 3496 1588 3498 1592
rect 3490 1586 3498 1588
rect 3514 1592 3522 1594
rect 3514 1588 3516 1592
rect 3520 1588 3522 1592
rect 3514 1586 3522 1588
rect 3538 1592 3546 1594
rect 3538 1588 3540 1592
rect 3544 1588 3546 1592
rect 3538 1586 3546 1588
rect 3562 1592 3570 1594
rect 3562 1588 3564 1592
rect 3568 1588 3570 1592
rect 3562 1586 3570 1588
rect 3586 1592 3594 1594
rect 3586 1588 3588 1592
rect 3592 1588 3594 1592
rect 3586 1586 3594 1588
rect 3610 1592 3618 1594
rect 3610 1588 3612 1592
rect 3616 1588 3618 1592
rect 3610 1586 3618 1588
rect 3634 1592 3642 1594
rect 3634 1588 3636 1592
rect 3640 1588 3642 1592
rect 3634 1586 3642 1588
rect 3658 1592 3666 1594
rect 3658 1588 3660 1592
rect 3664 1588 3666 1592
rect 3658 1586 3666 1588
rect 3682 1592 3690 1594
rect 3682 1588 3684 1592
rect 3688 1588 3690 1592
rect 3682 1586 3690 1588
rect 3898 1592 3906 1594
rect 3898 1588 3900 1592
rect 3904 1588 3906 1592
rect 3898 1586 3906 1588
rect 3922 1592 3930 1594
rect 3922 1588 3924 1592
rect 3928 1588 3930 1592
rect 3922 1586 3930 1588
rect 3946 1592 3954 1594
rect 3946 1588 3948 1592
rect 3952 1588 3954 1592
rect 3946 1586 3954 1588
rect 3970 1592 3978 1594
rect 3970 1588 3972 1592
rect 3976 1588 3978 1592
rect 3970 1586 3978 1588
rect 3994 1592 4002 1594
rect 3994 1588 3996 1592
rect 4000 1588 4002 1592
rect 3994 1586 4002 1588
rect 4018 1592 4026 1594
rect 4018 1588 4020 1592
rect 4024 1588 4026 1592
rect 4018 1586 4026 1588
rect 4042 1592 4050 1594
rect 4042 1588 4044 1592
rect 4048 1588 4050 1592
rect 4042 1586 4050 1588
rect 4066 1592 4074 1594
rect 4066 1588 4068 1592
rect 4072 1588 4074 1592
rect 4066 1586 4074 1588
rect 4090 1592 4098 1594
rect 4090 1588 4092 1592
rect 4096 1588 4098 1592
rect 4090 1586 4098 1588
rect 4114 1592 4122 1594
rect 4114 1588 4116 1592
rect 4120 1588 4122 1592
rect 4114 1586 4122 1588
rect 4138 1592 4146 1594
rect 4138 1588 4140 1592
rect 4144 1588 4146 1592
rect 4138 1586 4146 1588
rect 4162 1592 4170 1594
rect 4162 1588 4164 1592
rect 4168 1588 4170 1592
rect 4162 1586 4170 1588
rect 4186 1592 4194 1594
rect 4186 1588 4188 1592
rect 4192 1588 4194 1592
rect 4186 1586 4194 1588
rect 4210 1592 4218 1594
rect 4210 1588 4212 1592
rect 4216 1588 4218 1592
rect 4210 1586 4218 1588
rect 4234 1592 4242 1594
rect 4234 1588 4236 1592
rect 4240 1588 4242 1592
rect 4234 1586 4242 1588
rect 4258 1592 4266 1594
rect 4258 1588 4260 1592
rect 4264 1588 4266 1592
rect 4258 1586 4266 1588
rect 4282 1592 4290 1594
rect 4282 1588 4284 1592
rect 4288 1588 4290 1592
rect 4282 1586 4290 1588
rect 4498 1592 4506 1594
rect 4498 1588 4500 1592
rect 4504 1588 4506 1592
rect 4498 1586 4506 1588
rect 4522 1592 4530 1594
rect 4522 1588 4524 1592
rect 4528 1588 4530 1592
rect 4522 1586 4530 1588
rect 4546 1592 4554 1594
rect 4546 1588 4548 1592
rect 4552 1588 4554 1592
rect 4546 1586 4554 1588
rect 4570 1592 4578 1594
rect 4570 1588 4572 1592
rect 4576 1588 4578 1592
rect 4570 1586 4578 1588
rect 4594 1592 4602 1594
rect 4594 1588 4596 1592
rect 4600 1588 4602 1592
rect 4594 1586 4602 1588
rect 4618 1592 4626 1594
rect 4618 1588 4620 1592
rect 4624 1588 4626 1592
rect 4618 1586 4626 1588
rect 4642 1592 4650 1594
rect 4642 1588 4644 1592
rect 4648 1588 4650 1592
rect 4642 1586 4650 1588
rect 4666 1592 4674 1594
rect 4666 1588 4668 1592
rect 4672 1588 4674 1592
rect 4666 1586 4674 1588
rect 4690 1592 4698 1594
rect 4690 1588 4692 1592
rect 4696 1588 4698 1592
rect 4690 1586 4698 1588
rect 4714 1592 4722 1594
rect 4714 1588 4716 1592
rect 4720 1588 4722 1592
rect 4714 1586 4722 1588
rect 4738 1592 4746 1594
rect 4738 1588 4740 1592
rect 4744 1588 4746 1592
rect 4738 1586 4746 1588
rect 4762 1592 4770 1594
rect 4762 1588 4764 1592
rect 4768 1588 4770 1592
rect 4762 1586 4770 1588
rect 4786 1592 4794 1594
rect 4786 1588 4788 1592
rect 4792 1588 4794 1592
rect 4786 1586 4794 1588
rect 4810 1592 4818 1594
rect 4810 1588 4812 1592
rect 4816 1588 4818 1592
rect 4810 1586 4818 1588
rect 4834 1592 4842 1594
rect 4834 1588 4836 1592
rect 4840 1588 4842 1592
rect 4834 1586 4842 1588
rect 4858 1592 4866 1594
rect 4858 1588 4860 1592
rect 4864 1588 4866 1592
rect 4858 1586 4866 1588
rect 4882 1592 4890 1594
rect 4882 1588 4884 1592
rect 4888 1588 4890 1592
rect 4882 1586 4890 1588
rect 5698 1592 5706 1594
rect 5698 1588 5700 1592
rect 5704 1588 5706 1592
rect 5698 1586 5706 1588
rect 5722 1592 5730 1594
rect 5722 1588 5724 1592
rect 5728 1588 5730 1592
rect 5722 1586 5730 1588
rect 5746 1592 5754 1594
rect 5746 1588 5748 1592
rect 5752 1588 5754 1592
rect 5746 1586 5754 1588
rect 5770 1592 5778 1594
rect 5770 1588 5772 1592
rect 5776 1588 5778 1592
rect 5770 1586 5778 1588
rect 5794 1592 5802 1594
rect 5794 1588 5796 1592
rect 5800 1588 5802 1592
rect 5794 1586 5802 1588
rect 5818 1592 5826 1594
rect 5818 1588 5820 1592
rect 5824 1588 5826 1592
rect 5818 1586 5826 1588
rect 5842 1592 5850 1594
rect 5842 1588 5844 1592
rect 5848 1588 5850 1592
rect 5842 1586 5850 1588
rect 5866 1592 5874 1594
rect 5866 1588 5868 1592
rect 5872 1588 5874 1592
rect 5866 1586 5874 1588
rect 5890 1592 5898 1594
rect 5890 1588 5892 1592
rect 5896 1588 5898 1592
rect 5890 1586 5898 1588
rect 5914 1592 5922 1594
rect 5914 1588 5916 1592
rect 5920 1588 5922 1592
rect 5914 1586 5922 1588
rect 5938 1592 5946 1594
rect 5938 1588 5940 1592
rect 5944 1588 5946 1592
rect 5938 1586 5946 1588
rect 5962 1592 5970 1594
rect 5962 1588 5964 1592
rect 5968 1588 5970 1592
rect 5962 1586 5970 1588
rect 5986 1592 5994 1594
rect 5986 1588 5988 1592
rect 5992 1588 5994 1592
rect 5986 1586 5994 1588
rect 6010 1592 6018 1594
rect 6010 1588 6012 1592
rect 6016 1588 6018 1592
rect 6010 1586 6018 1588
rect 6034 1592 6042 1594
rect 6034 1588 6036 1592
rect 6040 1588 6042 1592
rect 6034 1586 6042 1588
rect 6058 1592 6066 1594
rect 6058 1588 6060 1592
rect 6064 1588 6066 1592
rect 6058 1586 6066 1588
rect 6082 1592 6090 1594
rect 6082 1588 6084 1592
rect 6088 1588 6090 1592
rect 6082 1586 6090 1588
rect 6298 1592 6306 1594
rect 6298 1588 6300 1592
rect 6304 1588 6306 1592
rect 6298 1586 6306 1588
rect 6322 1592 6330 1594
rect 6322 1588 6324 1592
rect 6328 1588 6330 1592
rect 6322 1586 6330 1588
rect 6346 1592 6354 1594
rect 6346 1588 6348 1592
rect 6352 1588 6354 1592
rect 6346 1586 6354 1588
rect 6370 1592 6378 1594
rect 6370 1588 6372 1592
rect 6376 1588 6378 1592
rect 6370 1586 6378 1588
rect 6394 1592 6402 1594
rect 6394 1588 6396 1592
rect 6400 1588 6402 1592
rect 6394 1586 6402 1588
rect 6418 1592 6426 1594
rect 6418 1588 6420 1592
rect 6424 1588 6426 1592
rect 6418 1586 6426 1588
rect 6442 1592 6450 1594
rect 6442 1588 6444 1592
rect 6448 1588 6450 1592
rect 6442 1586 6450 1588
rect 6466 1592 6474 1594
rect 6466 1588 6468 1592
rect 6472 1588 6474 1592
rect 6466 1586 6474 1588
rect 6490 1592 6498 1594
rect 6490 1588 6492 1592
rect 6496 1588 6498 1592
rect 6490 1586 6498 1588
rect 6514 1592 6522 1594
rect 6514 1588 6516 1592
rect 6520 1588 6522 1592
rect 6514 1586 6522 1588
rect 6538 1592 6546 1594
rect 6538 1588 6540 1592
rect 6544 1588 6546 1592
rect 6538 1586 6546 1588
rect 6562 1592 6570 1594
rect 6562 1588 6564 1592
rect 6568 1588 6570 1592
rect 6562 1586 6570 1588
rect 6586 1592 6594 1594
rect 6586 1588 6588 1592
rect 6592 1588 6594 1592
rect 6586 1586 6594 1588
rect 6610 1592 6618 1594
rect 6610 1588 6612 1592
rect 6616 1588 6618 1592
rect 6610 1586 6618 1588
rect 6634 1592 6642 1594
rect 6634 1588 6636 1592
rect 6640 1588 6642 1592
rect 6634 1586 6642 1588
rect 6658 1592 6666 1594
rect 6658 1588 6660 1592
rect 6664 1588 6666 1592
rect 6658 1586 6666 1588
rect 6682 1592 6690 1594
rect 6682 1588 6684 1592
rect 6688 1588 6690 1592
rect 6682 1586 6690 1588
rect 6898 1592 6906 1594
rect 6898 1588 6900 1592
rect 6904 1588 6906 1592
rect 6898 1586 6906 1588
rect 6922 1592 6930 1594
rect 6922 1588 6924 1592
rect 6928 1588 6930 1592
rect 6922 1586 6930 1588
rect 6946 1592 6954 1594
rect 6946 1588 6948 1592
rect 6952 1588 6954 1592
rect 6946 1586 6954 1588
rect 6970 1592 6978 1594
rect 6970 1588 6972 1592
rect 6976 1588 6978 1592
rect 6970 1586 6978 1588
rect 6994 1592 7002 1594
rect 6994 1588 6996 1592
rect 7000 1588 7002 1592
rect 6994 1586 7002 1588
rect 7018 1592 7026 1594
rect 7018 1588 7020 1592
rect 7024 1588 7026 1592
rect 7018 1586 7026 1588
rect 7042 1592 7050 1594
rect 7042 1588 7044 1592
rect 7048 1588 7050 1592
rect 7042 1586 7050 1588
rect 7066 1592 7074 1594
rect 7066 1588 7068 1592
rect 7072 1588 7074 1592
rect 7066 1586 7074 1588
rect 7090 1592 7098 1594
rect 7090 1588 7092 1592
rect 7096 1588 7098 1592
rect 7090 1586 7098 1588
rect 7114 1592 7122 1594
rect 7114 1588 7116 1592
rect 7120 1588 7122 1592
rect 7114 1586 7122 1588
rect 7138 1592 7146 1594
rect 7138 1588 7140 1592
rect 7144 1588 7146 1592
rect 7138 1586 7146 1588
rect 7162 1592 7170 1594
rect 7162 1588 7164 1592
rect 7168 1588 7170 1592
rect 7162 1586 7170 1588
rect 7186 1592 7194 1594
rect 7186 1588 7188 1592
rect 7192 1588 7194 1592
rect 7186 1586 7194 1588
rect 2110 1580 2118 1582
rect 2110 1576 2112 1580
rect 2116 1576 2118 1580
rect 2110 1574 2118 1576
rect 2134 1580 2142 1582
rect 2134 1576 2136 1580
rect 2140 1576 2142 1580
rect 2134 1574 2142 1576
rect 2158 1580 2166 1582
rect 2158 1576 2160 1580
rect 2164 1576 2166 1580
rect 2158 1574 2166 1576
rect 2182 1580 2190 1582
rect 2182 1576 2184 1580
rect 2188 1576 2190 1580
rect 2182 1574 2190 1576
rect 2206 1580 2214 1582
rect 2206 1576 2208 1580
rect 2212 1576 2214 1580
rect 2206 1574 2214 1576
rect 2230 1580 2238 1582
rect 2230 1576 2232 1580
rect 2236 1576 2238 1580
rect 2230 1574 2238 1576
rect 2254 1580 2262 1582
rect 2254 1576 2256 1580
rect 2260 1576 2262 1580
rect 2254 1574 2262 1576
rect 2278 1580 2286 1582
rect 2278 1576 2280 1580
rect 2284 1576 2286 1580
rect 2278 1574 2286 1576
rect 2302 1580 2310 1582
rect 2302 1576 2304 1580
rect 2308 1576 2310 1580
rect 2302 1574 2310 1576
rect 2326 1580 2334 1582
rect 2326 1576 2328 1580
rect 2332 1576 2334 1580
rect 2326 1574 2334 1576
rect 2350 1580 2358 1582
rect 2350 1576 2352 1580
rect 2356 1576 2358 1580
rect 2350 1574 2358 1576
rect 2374 1580 2382 1582
rect 2374 1576 2376 1580
rect 2380 1576 2382 1580
rect 2374 1574 2382 1576
rect 2398 1580 2406 1582
rect 2398 1576 2400 1580
rect 2404 1576 2406 1580
rect 2398 1574 2406 1576
rect 2422 1580 2430 1582
rect 2422 1576 2424 1580
rect 2428 1576 2430 1580
rect 2422 1574 2430 1576
rect 2446 1580 2454 1582
rect 2446 1576 2448 1580
rect 2452 1576 2454 1580
rect 2446 1574 2454 1576
rect 2470 1580 2478 1582
rect 2470 1576 2472 1580
rect 2476 1576 2478 1580
rect 2470 1574 2478 1576
rect 2494 1580 2502 1582
rect 2494 1576 2496 1580
rect 2500 1576 2502 1580
rect 2494 1574 2502 1576
rect 2710 1580 2718 1582
rect 2710 1576 2712 1580
rect 2716 1576 2718 1580
rect 2710 1574 2718 1576
rect 2734 1580 2742 1582
rect 2734 1576 2736 1580
rect 2740 1576 2742 1580
rect 2734 1574 2742 1576
rect 2758 1580 2766 1582
rect 2758 1576 2760 1580
rect 2764 1576 2766 1580
rect 2758 1574 2766 1576
rect 2782 1580 2790 1582
rect 2782 1576 2784 1580
rect 2788 1576 2790 1580
rect 2782 1574 2790 1576
rect 2806 1580 2814 1582
rect 2806 1576 2808 1580
rect 2812 1576 2814 1580
rect 2806 1574 2814 1576
rect 2830 1580 2838 1582
rect 2830 1576 2832 1580
rect 2836 1576 2838 1580
rect 2830 1574 2838 1576
rect 2854 1580 2862 1582
rect 2854 1576 2856 1580
rect 2860 1576 2862 1580
rect 2854 1574 2862 1576
rect 2878 1580 2886 1582
rect 2878 1576 2880 1580
rect 2884 1576 2886 1580
rect 2878 1574 2886 1576
rect 2902 1580 2910 1582
rect 2902 1576 2904 1580
rect 2908 1576 2910 1580
rect 2902 1574 2910 1576
rect 2926 1580 2934 1582
rect 2926 1576 2928 1580
rect 2932 1576 2934 1580
rect 2926 1574 2934 1576
rect 2950 1580 2958 1582
rect 2950 1576 2952 1580
rect 2956 1576 2958 1580
rect 2950 1574 2958 1576
rect 2974 1580 2982 1582
rect 2974 1576 2976 1580
rect 2980 1576 2982 1580
rect 2974 1574 2982 1576
rect 2998 1580 3006 1582
rect 2998 1576 3000 1580
rect 3004 1576 3006 1580
rect 2998 1574 3006 1576
rect 3022 1580 3030 1582
rect 3022 1576 3024 1580
rect 3028 1576 3030 1580
rect 3022 1574 3030 1576
rect 3046 1580 3054 1582
rect 3046 1576 3048 1580
rect 3052 1576 3054 1580
rect 3046 1574 3054 1576
rect 3070 1580 3078 1582
rect 3070 1576 3072 1580
rect 3076 1576 3078 1580
rect 3070 1574 3078 1576
rect 3094 1580 3102 1582
rect 3094 1576 3096 1580
rect 3100 1576 3102 1580
rect 3094 1574 3102 1576
rect 3310 1580 3318 1582
rect 3310 1576 3312 1580
rect 3316 1576 3318 1580
rect 3310 1574 3318 1576
rect 3334 1580 3342 1582
rect 3334 1576 3336 1580
rect 3340 1576 3342 1580
rect 3334 1574 3342 1576
rect 3358 1580 3366 1582
rect 3358 1576 3360 1580
rect 3364 1576 3366 1580
rect 3358 1574 3366 1576
rect 3382 1580 3390 1582
rect 3382 1576 3384 1580
rect 3388 1576 3390 1580
rect 3382 1574 3390 1576
rect 3406 1580 3414 1582
rect 3406 1576 3408 1580
rect 3412 1576 3414 1580
rect 3406 1574 3414 1576
rect 3430 1580 3438 1582
rect 3430 1576 3432 1580
rect 3436 1576 3438 1580
rect 3430 1574 3438 1576
rect 3454 1580 3462 1582
rect 3454 1576 3456 1580
rect 3460 1576 3462 1580
rect 3454 1574 3462 1576
rect 3478 1580 3486 1582
rect 3478 1576 3480 1580
rect 3484 1576 3486 1580
rect 3478 1574 3486 1576
rect 3502 1580 3510 1582
rect 3502 1576 3504 1580
rect 3508 1576 3510 1580
rect 3502 1574 3510 1576
rect 3526 1580 3534 1582
rect 3526 1576 3528 1580
rect 3532 1576 3534 1580
rect 3526 1574 3534 1576
rect 3550 1580 3558 1582
rect 3550 1576 3552 1580
rect 3556 1576 3558 1580
rect 3550 1574 3558 1576
rect 3574 1580 3582 1582
rect 3574 1576 3576 1580
rect 3580 1576 3582 1580
rect 3574 1574 3582 1576
rect 3598 1580 3606 1582
rect 3598 1576 3600 1580
rect 3604 1576 3606 1580
rect 3598 1574 3606 1576
rect 3622 1580 3630 1582
rect 3622 1576 3624 1580
rect 3628 1576 3630 1580
rect 3622 1574 3630 1576
rect 3646 1580 3654 1582
rect 3646 1576 3648 1580
rect 3652 1576 3654 1580
rect 3646 1574 3654 1576
rect 3670 1580 3678 1582
rect 3670 1576 3672 1580
rect 3676 1576 3678 1580
rect 3670 1574 3678 1576
rect 3694 1580 3702 1582
rect 3694 1576 3696 1580
rect 3700 1576 3702 1580
rect 3694 1574 3702 1576
rect 3910 1580 3918 1582
rect 3910 1576 3912 1580
rect 3916 1576 3918 1580
rect 3910 1574 3918 1576
rect 3934 1580 3942 1582
rect 3934 1576 3936 1580
rect 3940 1576 3942 1580
rect 3934 1574 3942 1576
rect 3958 1580 3966 1582
rect 3958 1576 3960 1580
rect 3964 1576 3966 1580
rect 3958 1574 3966 1576
rect 3982 1580 3990 1582
rect 3982 1576 3984 1580
rect 3988 1576 3990 1580
rect 3982 1574 3990 1576
rect 4006 1580 4014 1582
rect 4006 1576 4008 1580
rect 4012 1576 4014 1580
rect 4006 1574 4014 1576
rect 4030 1580 4038 1582
rect 4030 1576 4032 1580
rect 4036 1576 4038 1580
rect 4030 1574 4038 1576
rect 4054 1580 4062 1582
rect 4054 1576 4056 1580
rect 4060 1576 4062 1580
rect 4054 1574 4062 1576
rect 4078 1580 4086 1582
rect 4078 1576 4080 1580
rect 4084 1576 4086 1580
rect 4078 1574 4086 1576
rect 4102 1580 4110 1582
rect 4102 1576 4104 1580
rect 4108 1576 4110 1580
rect 4102 1574 4110 1576
rect 4126 1580 4134 1582
rect 4126 1576 4128 1580
rect 4132 1576 4134 1580
rect 4126 1574 4134 1576
rect 4150 1580 4158 1582
rect 4150 1576 4152 1580
rect 4156 1576 4158 1580
rect 4150 1574 4158 1576
rect 4174 1580 4182 1582
rect 4174 1576 4176 1580
rect 4180 1576 4182 1580
rect 4174 1574 4182 1576
rect 4198 1580 4206 1582
rect 4198 1576 4200 1580
rect 4204 1576 4206 1580
rect 4198 1574 4206 1576
rect 4222 1580 4230 1582
rect 4222 1576 4224 1580
rect 4228 1576 4230 1580
rect 4222 1574 4230 1576
rect 4246 1580 4254 1582
rect 4246 1576 4248 1580
rect 4252 1576 4254 1580
rect 4246 1574 4254 1576
rect 4270 1580 4278 1582
rect 4270 1576 4272 1580
rect 4276 1576 4278 1580
rect 4270 1574 4278 1576
rect 4294 1580 4302 1582
rect 4294 1576 4296 1580
rect 4300 1576 4302 1580
rect 4294 1574 4302 1576
rect 4510 1580 4518 1582
rect 4510 1576 4512 1580
rect 4516 1576 4518 1580
rect 4510 1574 4518 1576
rect 4534 1580 4542 1582
rect 4534 1576 4536 1580
rect 4540 1576 4542 1580
rect 4534 1574 4542 1576
rect 4558 1580 4566 1582
rect 4558 1576 4560 1580
rect 4564 1576 4566 1580
rect 4558 1574 4566 1576
rect 4582 1580 4590 1582
rect 4582 1576 4584 1580
rect 4588 1576 4590 1580
rect 4582 1574 4590 1576
rect 4606 1580 4614 1582
rect 4606 1576 4608 1580
rect 4612 1576 4614 1580
rect 4606 1574 4614 1576
rect 4630 1580 4638 1582
rect 4630 1576 4632 1580
rect 4636 1576 4638 1580
rect 4630 1574 4638 1576
rect 4654 1580 4662 1582
rect 4654 1576 4656 1580
rect 4660 1576 4662 1580
rect 4654 1574 4662 1576
rect 4678 1580 4686 1582
rect 4678 1576 4680 1580
rect 4684 1576 4686 1580
rect 4678 1574 4686 1576
rect 4702 1580 4710 1582
rect 4702 1576 4704 1580
rect 4708 1576 4710 1580
rect 4702 1574 4710 1576
rect 4726 1580 4734 1582
rect 4726 1576 4728 1580
rect 4732 1576 4734 1580
rect 4726 1574 4734 1576
rect 4750 1580 4758 1582
rect 4750 1576 4752 1580
rect 4756 1576 4758 1580
rect 4750 1574 4758 1576
rect 4774 1580 4782 1582
rect 4774 1576 4776 1580
rect 4780 1576 4782 1580
rect 4774 1574 4782 1576
rect 4798 1580 4806 1582
rect 4798 1576 4800 1580
rect 4804 1576 4806 1580
rect 4798 1574 4806 1576
rect 4822 1580 4830 1582
rect 4822 1576 4824 1580
rect 4828 1576 4830 1580
rect 4822 1574 4830 1576
rect 4846 1580 4854 1582
rect 4846 1576 4848 1580
rect 4852 1576 4854 1580
rect 4846 1574 4854 1576
rect 4870 1580 4878 1582
rect 4870 1576 4872 1580
rect 4876 1576 4878 1580
rect 4870 1574 4878 1576
rect 4894 1580 4902 1582
rect 4894 1576 4896 1580
rect 4900 1576 4902 1580
rect 4894 1574 4902 1576
rect 5710 1580 5718 1582
rect 5710 1576 5712 1580
rect 5716 1576 5718 1580
rect 5710 1574 5718 1576
rect 5734 1580 5742 1582
rect 5734 1576 5736 1580
rect 5740 1576 5742 1580
rect 5734 1574 5742 1576
rect 5758 1580 5766 1582
rect 5758 1576 5760 1580
rect 5764 1576 5766 1580
rect 5758 1574 5766 1576
rect 5782 1580 5790 1582
rect 5782 1576 5784 1580
rect 5788 1576 5790 1580
rect 5782 1574 5790 1576
rect 5806 1580 5814 1582
rect 5806 1576 5808 1580
rect 5812 1576 5814 1580
rect 5806 1574 5814 1576
rect 5830 1580 5838 1582
rect 5830 1576 5832 1580
rect 5836 1576 5838 1580
rect 5830 1574 5838 1576
rect 5854 1580 5862 1582
rect 5854 1576 5856 1580
rect 5860 1576 5862 1580
rect 5854 1574 5862 1576
rect 5878 1580 5886 1582
rect 5878 1576 5880 1580
rect 5884 1576 5886 1580
rect 5878 1574 5886 1576
rect 5902 1580 5910 1582
rect 5902 1576 5904 1580
rect 5908 1576 5910 1580
rect 5902 1574 5910 1576
rect 5926 1580 5934 1582
rect 5926 1576 5928 1580
rect 5932 1576 5934 1580
rect 5926 1574 5934 1576
rect 5950 1580 5958 1582
rect 5950 1576 5952 1580
rect 5956 1576 5958 1580
rect 5950 1574 5958 1576
rect 5974 1580 5982 1582
rect 5974 1576 5976 1580
rect 5980 1576 5982 1580
rect 5974 1574 5982 1576
rect 5998 1580 6006 1582
rect 5998 1576 6000 1580
rect 6004 1576 6006 1580
rect 5998 1574 6006 1576
rect 6022 1580 6030 1582
rect 6022 1576 6024 1580
rect 6028 1576 6030 1580
rect 6022 1574 6030 1576
rect 6046 1580 6054 1582
rect 6046 1576 6048 1580
rect 6052 1576 6054 1580
rect 6046 1574 6054 1576
rect 6070 1580 6078 1582
rect 6070 1576 6072 1580
rect 6076 1576 6078 1580
rect 6070 1574 6078 1576
rect 6094 1580 6102 1582
rect 6094 1576 6096 1580
rect 6100 1576 6102 1580
rect 6094 1574 6102 1576
rect 6310 1580 6318 1582
rect 6310 1576 6312 1580
rect 6316 1576 6318 1580
rect 6310 1574 6318 1576
rect 6334 1580 6342 1582
rect 6334 1576 6336 1580
rect 6340 1576 6342 1580
rect 6334 1574 6342 1576
rect 6358 1580 6366 1582
rect 6358 1576 6360 1580
rect 6364 1576 6366 1580
rect 6358 1574 6366 1576
rect 6382 1580 6390 1582
rect 6382 1576 6384 1580
rect 6388 1576 6390 1580
rect 6382 1574 6390 1576
rect 6406 1580 6414 1582
rect 6406 1576 6408 1580
rect 6412 1576 6414 1580
rect 6406 1574 6414 1576
rect 6430 1580 6438 1582
rect 6430 1576 6432 1580
rect 6436 1576 6438 1580
rect 6430 1574 6438 1576
rect 6454 1580 6462 1582
rect 6454 1576 6456 1580
rect 6460 1576 6462 1580
rect 6454 1574 6462 1576
rect 6478 1580 6486 1582
rect 6478 1576 6480 1580
rect 6484 1576 6486 1580
rect 6478 1574 6486 1576
rect 6502 1580 6510 1582
rect 6502 1576 6504 1580
rect 6508 1576 6510 1580
rect 6502 1574 6510 1576
rect 6526 1580 6534 1582
rect 6526 1576 6528 1580
rect 6532 1576 6534 1580
rect 6526 1574 6534 1576
rect 6550 1580 6558 1582
rect 6550 1576 6552 1580
rect 6556 1576 6558 1580
rect 6550 1574 6558 1576
rect 6574 1580 6582 1582
rect 6574 1576 6576 1580
rect 6580 1576 6582 1580
rect 6574 1574 6582 1576
rect 6598 1580 6606 1582
rect 6598 1576 6600 1580
rect 6604 1576 6606 1580
rect 6598 1574 6606 1576
rect 6622 1580 6630 1582
rect 6622 1576 6624 1580
rect 6628 1576 6630 1580
rect 6622 1574 6630 1576
rect 6646 1580 6654 1582
rect 6646 1576 6648 1580
rect 6652 1576 6654 1580
rect 6646 1574 6654 1576
rect 6670 1580 6678 1582
rect 6670 1576 6672 1580
rect 6676 1576 6678 1580
rect 6670 1574 6678 1576
rect 6694 1580 6702 1582
rect 6694 1576 6696 1580
rect 6700 1576 6702 1580
rect 6694 1574 6702 1576
rect 6910 1580 6918 1582
rect 6910 1576 6912 1580
rect 6916 1576 6918 1580
rect 6910 1574 6918 1576
rect 6934 1580 6942 1582
rect 6934 1576 6936 1580
rect 6940 1576 6942 1580
rect 6934 1574 6942 1576
rect 6958 1580 6966 1582
rect 6958 1576 6960 1580
rect 6964 1576 6966 1580
rect 6958 1574 6966 1576
rect 6982 1580 6990 1582
rect 6982 1576 6984 1580
rect 6988 1576 6990 1580
rect 6982 1574 6990 1576
rect 7006 1580 7014 1582
rect 7006 1576 7008 1580
rect 7012 1576 7014 1580
rect 7006 1574 7014 1576
rect 7030 1580 7038 1582
rect 7030 1576 7032 1580
rect 7036 1576 7038 1580
rect 7030 1574 7038 1576
rect 7054 1580 7062 1582
rect 7054 1576 7056 1580
rect 7060 1576 7062 1580
rect 7054 1574 7062 1576
rect 7078 1580 7086 1582
rect 7078 1576 7080 1580
rect 7084 1576 7086 1580
rect 7078 1574 7086 1576
rect 7102 1580 7110 1582
rect 7102 1576 7104 1580
rect 7108 1576 7110 1580
rect 7102 1574 7110 1576
rect 7126 1580 7134 1582
rect 7126 1576 7128 1580
rect 7132 1576 7134 1580
rect 7126 1574 7134 1576
rect 7150 1580 7158 1582
rect 7150 1576 7152 1580
rect 7156 1576 7158 1580
rect 7150 1574 7158 1576
rect 7174 1580 7182 1582
rect 7174 1576 7176 1580
rect 7180 1576 7182 1580
rect 7174 1574 7182 1576
rect 7198 1574 7200 1582
rect 2098 1568 2106 1570
rect 2098 1564 2100 1568
rect 2104 1564 2106 1568
rect 2098 1562 2106 1564
rect 2122 1568 2130 1570
rect 2122 1564 2124 1568
rect 2128 1564 2130 1568
rect 2122 1562 2130 1564
rect 2146 1568 2154 1570
rect 2146 1564 2148 1568
rect 2152 1564 2154 1568
rect 2146 1562 2154 1564
rect 2170 1568 2178 1570
rect 2170 1564 2172 1568
rect 2176 1564 2178 1568
rect 2170 1562 2178 1564
rect 2194 1568 2202 1570
rect 2194 1564 2196 1568
rect 2200 1564 2202 1568
rect 2194 1562 2202 1564
rect 2218 1568 2226 1570
rect 2218 1564 2220 1568
rect 2224 1564 2226 1568
rect 2218 1562 2226 1564
rect 2242 1568 2250 1570
rect 2242 1564 2244 1568
rect 2248 1564 2250 1568
rect 2242 1562 2250 1564
rect 2266 1568 2274 1570
rect 2266 1564 2268 1568
rect 2272 1564 2274 1568
rect 2266 1562 2274 1564
rect 2290 1568 2298 1570
rect 2290 1564 2292 1568
rect 2296 1564 2298 1568
rect 2290 1562 2298 1564
rect 2314 1568 2322 1570
rect 2314 1564 2316 1568
rect 2320 1564 2322 1568
rect 2314 1562 2322 1564
rect 2338 1568 2346 1570
rect 2338 1564 2340 1568
rect 2344 1564 2346 1568
rect 2338 1562 2346 1564
rect 2362 1568 2370 1570
rect 2362 1564 2364 1568
rect 2368 1564 2370 1568
rect 2362 1562 2370 1564
rect 2386 1568 2394 1570
rect 2386 1564 2388 1568
rect 2392 1564 2394 1568
rect 2386 1562 2394 1564
rect 2410 1568 2418 1570
rect 2410 1564 2412 1568
rect 2416 1564 2418 1568
rect 2410 1562 2418 1564
rect 2434 1568 2442 1570
rect 2434 1564 2436 1568
rect 2440 1564 2442 1568
rect 2434 1562 2442 1564
rect 2458 1568 2466 1570
rect 2458 1564 2460 1568
rect 2464 1564 2466 1568
rect 2458 1562 2466 1564
rect 2482 1568 2490 1570
rect 2482 1564 2484 1568
rect 2488 1564 2490 1568
rect 2482 1562 2490 1564
rect 2698 1568 2706 1570
rect 2698 1564 2700 1568
rect 2704 1564 2706 1568
rect 2698 1562 2706 1564
rect 2722 1568 2730 1570
rect 2722 1564 2724 1568
rect 2728 1564 2730 1568
rect 2722 1562 2730 1564
rect 2746 1568 2754 1570
rect 2746 1564 2748 1568
rect 2752 1564 2754 1568
rect 2746 1562 2754 1564
rect 2770 1568 2778 1570
rect 2770 1564 2772 1568
rect 2776 1564 2778 1568
rect 2770 1562 2778 1564
rect 2794 1568 2802 1570
rect 2794 1564 2796 1568
rect 2800 1564 2802 1568
rect 2794 1562 2802 1564
rect 2818 1568 2826 1570
rect 2818 1564 2820 1568
rect 2824 1564 2826 1568
rect 2818 1562 2826 1564
rect 2842 1568 2850 1570
rect 2842 1564 2844 1568
rect 2848 1564 2850 1568
rect 2842 1562 2850 1564
rect 2866 1568 2874 1570
rect 2866 1564 2868 1568
rect 2872 1564 2874 1568
rect 2866 1562 2874 1564
rect 2890 1568 2898 1570
rect 2890 1564 2892 1568
rect 2896 1564 2898 1568
rect 2890 1562 2898 1564
rect 2914 1568 2922 1570
rect 2914 1564 2916 1568
rect 2920 1564 2922 1568
rect 2914 1562 2922 1564
rect 2938 1568 2946 1570
rect 2938 1564 2940 1568
rect 2944 1564 2946 1568
rect 2938 1562 2946 1564
rect 2962 1568 2970 1570
rect 2962 1564 2964 1568
rect 2968 1564 2970 1568
rect 2962 1562 2970 1564
rect 2986 1568 2994 1570
rect 2986 1564 2988 1568
rect 2992 1564 2994 1568
rect 2986 1562 2994 1564
rect 3010 1568 3018 1570
rect 3010 1564 3012 1568
rect 3016 1564 3018 1568
rect 3010 1562 3018 1564
rect 3034 1568 3042 1570
rect 3034 1564 3036 1568
rect 3040 1564 3042 1568
rect 3034 1562 3042 1564
rect 3058 1568 3066 1570
rect 3058 1564 3060 1568
rect 3064 1564 3066 1568
rect 3058 1562 3066 1564
rect 3082 1568 3090 1570
rect 3082 1564 3084 1568
rect 3088 1564 3090 1568
rect 3082 1562 3090 1564
rect 3298 1568 3306 1570
rect 3298 1564 3300 1568
rect 3304 1564 3306 1568
rect 3298 1562 3306 1564
rect 3322 1568 3330 1570
rect 3322 1564 3324 1568
rect 3328 1564 3330 1568
rect 3322 1562 3330 1564
rect 3346 1568 3354 1570
rect 3346 1564 3348 1568
rect 3352 1564 3354 1568
rect 3346 1562 3354 1564
rect 3370 1568 3378 1570
rect 3370 1564 3372 1568
rect 3376 1564 3378 1568
rect 3370 1562 3378 1564
rect 3394 1568 3402 1570
rect 3394 1564 3396 1568
rect 3400 1564 3402 1568
rect 3394 1562 3402 1564
rect 3418 1568 3426 1570
rect 3418 1564 3420 1568
rect 3424 1564 3426 1568
rect 3418 1562 3426 1564
rect 3442 1568 3450 1570
rect 3442 1564 3444 1568
rect 3448 1564 3450 1568
rect 3442 1562 3450 1564
rect 3466 1568 3474 1570
rect 3466 1564 3468 1568
rect 3472 1564 3474 1568
rect 3466 1562 3474 1564
rect 3490 1568 3498 1570
rect 3490 1564 3492 1568
rect 3496 1564 3498 1568
rect 3490 1562 3498 1564
rect 3514 1568 3522 1570
rect 3514 1564 3516 1568
rect 3520 1564 3522 1568
rect 3514 1562 3522 1564
rect 3538 1568 3546 1570
rect 3538 1564 3540 1568
rect 3544 1564 3546 1568
rect 3538 1562 3546 1564
rect 3562 1568 3570 1570
rect 3562 1564 3564 1568
rect 3568 1564 3570 1568
rect 3562 1562 3570 1564
rect 3586 1568 3594 1570
rect 3586 1564 3588 1568
rect 3592 1564 3594 1568
rect 3586 1562 3594 1564
rect 3610 1568 3618 1570
rect 3610 1564 3612 1568
rect 3616 1564 3618 1568
rect 3610 1562 3618 1564
rect 3634 1568 3642 1570
rect 3634 1564 3636 1568
rect 3640 1564 3642 1568
rect 3634 1562 3642 1564
rect 3658 1568 3666 1570
rect 3658 1564 3660 1568
rect 3664 1564 3666 1568
rect 3658 1562 3666 1564
rect 3682 1568 3690 1570
rect 3682 1564 3684 1568
rect 3688 1564 3690 1568
rect 3682 1562 3690 1564
rect 3898 1568 3906 1570
rect 3898 1564 3900 1568
rect 3904 1564 3906 1568
rect 3898 1562 3906 1564
rect 3922 1568 3930 1570
rect 3922 1564 3924 1568
rect 3928 1564 3930 1568
rect 3922 1562 3930 1564
rect 3946 1568 3954 1570
rect 3946 1564 3948 1568
rect 3952 1564 3954 1568
rect 3946 1562 3954 1564
rect 3970 1568 3978 1570
rect 3970 1564 3972 1568
rect 3976 1564 3978 1568
rect 3970 1562 3978 1564
rect 3994 1568 4002 1570
rect 3994 1564 3996 1568
rect 4000 1564 4002 1568
rect 3994 1562 4002 1564
rect 4018 1568 4026 1570
rect 4018 1564 4020 1568
rect 4024 1564 4026 1568
rect 4018 1562 4026 1564
rect 4042 1568 4050 1570
rect 4042 1564 4044 1568
rect 4048 1564 4050 1568
rect 4042 1562 4050 1564
rect 4066 1568 4074 1570
rect 4066 1564 4068 1568
rect 4072 1564 4074 1568
rect 4066 1562 4074 1564
rect 4090 1568 4098 1570
rect 4090 1564 4092 1568
rect 4096 1564 4098 1568
rect 4090 1562 4098 1564
rect 4114 1568 4122 1570
rect 4114 1564 4116 1568
rect 4120 1564 4122 1568
rect 4114 1562 4122 1564
rect 4138 1568 4146 1570
rect 4138 1564 4140 1568
rect 4144 1564 4146 1568
rect 4138 1562 4146 1564
rect 4162 1568 4170 1570
rect 4162 1564 4164 1568
rect 4168 1564 4170 1568
rect 4162 1562 4170 1564
rect 4186 1568 4194 1570
rect 4186 1564 4188 1568
rect 4192 1564 4194 1568
rect 4186 1562 4194 1564
rect 4210 1568 4218 1570
rect 4210 1564 4212 1568
rect 4216 1564 4218 1568
rect 4210 1562 4218 1564
rect 4234 1568 4242 1570
rect 4234 1564 4236 1568
rect 4240 1564 4242 1568
rect 4234 1562 4242 1564
rect 4258 1568 4266 1570
rect 4258 1564 4260 1568
rect 4264 1564 4266 1568
rect 4258 1562 4266 1564
rect 4282 1568 4290 1570
rect 4282 1564 4284 1568
rect 4288 1564 4290 1568
rect 4282 1562 4290 1564
rect 4498 1568 4506 1570
rect 4498 1564 4500 1568
rect 4504 1564 4506 1568
rect 4498 1562 4506 1564
rect 4522 1568 4530 1570
rect 4522 1564 4524 1568
rect 4528 1564 4530 1568
rect 4522 1562 4530 1564
rect 4546 1568 4554 1570
rect 4546 1564 4548 1568
rect 4552 1564 4554 1568
rect 4546 1562 4554 1564
rect 4570 1568 4578 1570
rect 4570 1564 4572 1568
rect 4576 1564 4578 1568
rect 4570 1562 4578 1564
rect 4594 1568 4602 1570
rect 4594 1564 4596 1568
rect 4600 1564 4602 1568
rect 4594 1562 4602 1564
rect 4618 1568 4626 1570
rect 4618 1564 4620 1568
rect 4624 1564 4626 1568
rect 4618 1562 4626 1564
rect 4642 1568 4650 1570
rect 4642 1564 4644 1568
rect 4648 1564 4650 1568
rect 4642 1562 4650 1564
rect 4666 1568 4674 1570
rect 4666 1564 4668 1568
rect 4672 1564 4674 1568
rect 4666 1562 4674 1564
rect 4690 1568 4698 1570
rect 4690 1564 4692 1568
rect 4696 1564 4698 1568
rect 4690 1562 4698 1564
rect 4714 1568 4722 1570
rect 4714 1564 4716 1568
rect 4720 1564 4722 1568
rect 4714 1562 4722 1564
rect 4738 1568 4746 1570
rect 4738 1564 4740 1568
rect 4744 1564 4746 1568
rect 4738 1562 4746 1564
rect 4762 1568 4770 1570
rect 4762 1564 4764 1568
rect 4768 1564 4770 1568
rect 4762 1562 4770 1564
rect 4786 1568 4794 1570
rect 4786 1564 4788 1568
rect 4792 1564 4794 1568
rect 4786 1562 4794 1564
rect 4810 1568 4818 1570
rect 4810 1564 4812 1568
rect 4816 1564 4818 1568
rect 4810 1562 4818 1564
rect 4834 1568 4842 1570
rect 4834 1564 4836 1568
rect 4840 1564 4842 1568
rect 4834 1562 4842 1564
rect 4858 1568 4866 1570
rect 4858 1564 4860 1568
rect 4864 1564 4866 1568
rect 4858 1562 4866 1564
rect 4882 1568 4890 1570
rect 4882 1564 4884 1568
rect 4888 1564 4890 1568
rect 4882 1562 4890 1564
rect 5698 1568 5706 1570
rect 5698 1564 5700 1568
rect 5704 1564 5706 1568
rect 5698 1562 5706 1564
rect 5722 1568 5730 1570
rect 5722 1564 5724 1568
rect 5728 1564 5730 1568
rect 5722 1562 5730 1564
rect 5746 1568 5754 1570
rect 5746 1564 5748 1568
rect 5752 1564 5754 1568
rect 5746 1562 5754 1564
rect 5770 1568 5778 1570
rect 5770 1564 5772 1568
rect 5776 1564 5778 1568
rect 5770 1562 5778 1564
rect 5794 1568 5802 1570
rect 5794 1564 5796 1568
rect 5800 1564 5802 1568
rect 5794 1562 5802 1564
rect 5818 1568 5826 1570
rect 5818 1564 5820 1568
rect 5824 1564 5826 1568
rect 5818 1562 5826 1564
rect 5842 1568 5850 1570
rect 5842 1564 5844 1568
rect 5848 1564 5850 1568
rect 5842 1562 5850 1564
rect 5866 1568 5874 1570
rect 5866 1564 5868 1568
rect 5872 1564 5874 1568
rect 5866 1562 5874 1564
rect 5890 1568 5898 1570
rect 5890 1564 5892 1568
rect 5896 1564 5898 1568
rect 5890 1562 5898 1564
rect 5914 1568 5922 1570
rect 5914 1564 5916 1568
rect 5920 1564 5922 1568
rect 5914 1562 5922 1564
rect 5938 1568 5946 1570
rect 5938 1564 5940 1568
rect 5944 1564 5946 1568
rect 5938 1562 5946 1564
rect 5962 1568 5970 1570
rect 5962 1564 5964 1568
rect 5968 1564 5970 1568
rect 5962 1562 5970 1564
rect 5986 1568 5994 1570
rect 5986 1564 5988 1568
rect 5992 1564 5994 1568
rect 5986 1562 5994 1564
rect 6010 1568 6018 1570
rect 6010 1564 6012 1568
rect 6016 1564 6018 1568
rect 6010 1562 6018 1564
rect 6034 1568 6042 1570
rect 6034 1564 6036 1568
rect 6040 1564 6042 1568
rect 6034 1562 6042 1564
rect 6058 1568 6066 1570
rect 6058 1564 6060 1568
rect 6064 1564 6066 1568
rect 6058 1562 6066 1564
rect 6082 1568 6090 1570
rect 6082 1564 6084 1568
rect 6088 1564 6090 1568
rect 6082 1562 6090 1564
rect 6298 1568 6306 1570
rect 6298 1564 6300 1568
rect 6304 1564 6306 1568
rect 6298 1562 6306 1564
rect 6322 1568 6330 1570
rect 6322 1564 6324 1568
rect 6328 1564 6330 1568
rect 6322 1562 6330 1564
rect 6346 1568 6354 1570
rect 6346 1564 6348 1568
rect 6352 1564 6354 1568
rect 6346 1562 6354 1564
rect 6370 1568 6378 1570
rect 6370 1564 6372 1568
rect 6376 1564 6378 1568
rect 6370 1562 6378 1564
rect 6394 1568 6402 1570
rect 6394 1564 6396 1568
rect 6400 1564 6402 1568
rect 6394 1562 6402 1564
rect 6418 1568 6426 1570
rect 6418 1564 6420 1568
rect 6424 1564 6426 1568
rect 6418 1562 6426 1564
rect 6442 1568 6450 1570
rect 6442 1564 6444 1568
rect 6448 1564 6450 1568
rect 6442 1562 6450 1564
rect 6466 1568 6474 1570
rect 6466 1564 6468 1568
rect 6472 1564 6474 1568
rect 6466 1562 6474 1564
rect 6490 1568 6498 1570
rect 6490 1564 6492 1568
rect 6496 1564 6498 1568
rect 6490 1562 6498 1564
rect 6514 1568 6522 1570
rect 6514 1564 6516 1568
rect 6520 1564 6522 1568
rect 6514 1562 6522 1564
rect 6538 1568 6546 1570
rect 6538 1564 6540 1568
rect 6544 1564 6546 1568
rect 6538 1562 6546 1564
rect 6562 1568 6570 1570
rect 6562 1564 6564 1568
rect 6568 1564 6570 1568
rect 6562 1562 6570 1564
rect 6586 1568 6594 1570
rect 6586 1564 6588 1568
rect 6592 1564 6594 1568
rect 6586 1562 6594 1564
rect 6610 1568 6618 1570
rect 6610 1564 6612 1568
rect 6616 1564 6618 1568
rect 6610 1562 6618 1564
rect 6634 1568 6642 1570
rect 6634 1564 6636 1568
rect 6640 1564 6642 1568
rect 6634 1562 6642 1564
rect 6658 1568 6666 1570
rect 6658 1564 6660 1568
rect 6664 1564 6666 1568
rect 6658 1562 6666 1564
rect 6682 1568 6690 1570
rect 6682 1564 6684 1568
rect 6688 1564 6690 1568
rect 6682 1562 6690 1564
rect 6898 1568 6906 1570
rect 6898 1564 6900 1568
rect 6904 1564 6906 1568
rect 6898 1562 6906 1564
rect 6922 1568 6930 1570
rect 6922 1564 6924 1568
rect 6928 1564 6930 1568
rect 6922 1562 6930 1564
rect 6946 1568 6954 1570
rect 6946 1564 6948 1568
rect 6952 1564 6954 1568
rect 6946 1562 6954 1564
rect 6970 1568 6978 1570
rect 6970 1564 6972 1568
rect 6976 1564 6978 1568
rect 6970 1562 6978 1564
rect 6994 1568 7002 1570
rect 6994 1564 6996 1568
rect 7000 1564 7002 1568
rect 6994 1562 7002 1564
rect 7018 1568 7026 1570
rect 7018 1564 7020 1568
rect 7024 1564 7026 1568
rect 7018 1562 7026 1564
rect 7042 1568 7050 1570
rect 7042 1564 7044 1568
rect 7048 1564 7050 1568
rect 7042 1562 7050 1564
rect 7066 1568 7074 1570
rect 7066 1564 7068 1568
rect 7072 1564 7074 1568
rect 7066 1562 7074 1564
rect 7090 1568 7098 1570
rect 7090 1564 7092 1568
rect 7096 1564 7098 1568
rect 7090 1562 7098 1564
rect 7114 1568 7122 1570
rect 7114 1564 7116 1568
rect 7120 1564 7122 1568
rect 7114 1562 7122 1564
rect 7138 1568 7146 1570
rect 7138 1564 7140 1568
rect 7144 1564 7146 1568
rect 7138 1562 7146 1564
rect 7162 1568 7170 1570
rect 7162 1564 7164 1568
rect 7168 1564 7170 1568
rect 7162 1562 7170 1564
rect 7186 1568 7194 1570
rect 7186 1564 7188 1568
rect 7192 1564 7194 1568
rect 7186 1562 7194 1564
rect 2110 1556 2118 1558
rect 2110 1552 2112 1556
rect 2116 1552 2118 1556
rect 2110 1550 2118 1552
rect 2134 1556 2142 1558
rect 2134 1552 2136 1556
rect 2140 1552 2142 1556
rect 2134 1550 2142 1552
rect 2158 1556 2166 1558
rect 2158 1552 2160 1556
rect 2164 1552 2166 1556
rect 2158 1550 2166 1552
rect 2182 1556 2190 1558
rect 2182 1552 2184 1556
rect 2188 1552 2190 1556
rect 2182 1550 2190 1552
rect 2206 1556 2214 1558
rect 2206 1552 2208 1556
rect 2212 1552 2214 1556
rect 2206 1550 2214 1552
rect 2230 1556 2238 1558
rect 2230 1552 2232 1556
rect 2236 1552 2238 1556
rect 2230 1550 2238 1552
rect 2254 1556 2262 1558
rect 2254 1552 2256 1556
rect 2260 1552 2262 1556
rect 2254 1550 2262 1552
rect 2278 1556 2286 1558
rect 2278 1552 2280 1556
rect 2284 1552 2286 1556
rect 2278 1550 2286 1552
rect 2302 1556 2310 1558
rect 2302 1552 2304 1556
rect 2308 1552 2310 1556
rect 2302 1550 2310 1552
rect 2326 1556 2334 1558
rect 2326 1552 2328 1556
rect 2332 1552 2334 1556
rect 2326 1550 2334 1552
rect 2350 1556 2358 1558
rect 2350 1552 2352 1556
rect 2356 1552 2358 1556
rect 2350 1550 2358 1552
rect 2374 1556 2382 1558
rect 2374 1552 2376 1556
rect 2380 1552 2382 1556
rect 2374 1550 2382 1552
rect 2398 1556 2406 1558
rect 2398 1552 2400 1556
rect 2404 1552 2406 1556
rect 2398 1550 2406 1552
rect 2422 1556 2430 1558
rect 2422 1552 2424 1556
rect 2428 1552 2430 1556
rect 2422 1550 2430 1552
rect 2446 1556 2454 1558
rect 2446 1552 2448 1556
rect 2452 1552 2454 1556
rect 2446 1550 2454 1552
rect 2470 1556 2478 1558
rect 2470 1552 2472 1556
rect 2476 1552 2478 1556
rect 2470 1550 2478 1552
rect 2494 1556 2502 1558
rect 2494 1552 2496 1556
rect 2500 1552 2502 1556
rect 2494 1550 2502 1552
rect 2710 1556 2718 1558
rect 2710 1552 2712 1556
rect 2716 1552 2718 1556
rect 2710 1550 2718 1552
rect 2734 1556 2742 1558
rect 2734 1552 2736 1556
rect 2740 1552 2742 1556
rect 2734 1550 2742 1552
rect 2758 1556 2766 1558
rect 2758 1552 2760 1556
rect 2764 1552 2766 1556
rect 2758 1550 2766 1552
rect 2782 1556 2790 1558
rect 2782 1552 2784 1556
rect 2788 1552 2790 1556
rect 2782 1550 2790 1552
rect 2806 1556 2814 1558
rect 2806 1552 2808 1556
rect 2812 1552 2814 1556
rect 2806 1550 2814 1552
rect 2830 1556 2838 1558
rect 2830 1552 2832 1556
rect 2836 1552 2838 1556
rect 2830 1550 2838 1552
rect 2854 1556 2862 1558
rect 2854 1552 2856 1556
rect 2860 1552 2862 1556
rect 2854 1550 2862 1552
rect 2878 1556 2886 1558
rect 2878 1552 2880 1556
rect 2884 1552 2886 1556
rect 2878 1550 2886 1552
rect 2902 1556 2910 1558
rect 2902 1552 2904 1556
rect 2908 1552 2910 1556
rect 2902 1550 2910 1552
rect 2926 1556 2934 1558
rect 2926 1552 2928 1556
rect 2932 1552 2934 1556
rect 2926 1550 2934 1552
rect 2950 1556 2958 1558
rect 2950 1552 2952 1556
rect 2956 1552 2958 1556
rect 2950 1550 2958 1552
rect 2974 1556 2982 1558
rect 2974 1552 2976 1556
rect 2980 1552 2982 1556
rect 2974 1550 2982 1552
rect 2998 1556 3006 1558
rect 2998 1552 3000 1556
rect 3004 1552 3006 1556
rect 2998 1550 3006 1552
rect 3022 1556 3030 1558
rect 3022 1552 3024 1556
rect 3028 1552 3030 1556
rect 3022 1550 3030 1552
rect 3046 1556 3054 1558
rect 3046 1552 3048 1556
rect 3052 1552 3054 1556
rect 3046 1550 3054 1552
rect 3070 1556 3078 1558
rect 3070 1552 3072 1556
rect 3076 1552 3078 1556
rect 3070 1550 3078 1552
rect 3094 1556 3102 1558
rect 3094 1552 3096 1556
rect 3100 1552 3102 1556
rect 3094 1550 3102 1552
rect 3310 1556 3318 1558
rect 3310 1552 3312 1556
rect 3316 1552 3318 1556
rect 3310 1550 3318 1552
rect 3334 1556 3342 1558
rect 3334 1552 3336 1556
rect 3340 1552 3342 1556
rect 3334 1550 3342 1552
rect 3358 1556 3366 1558
rect 3358 1552 3360 1556
rect 3364 1552 3366 1556
rect 3358 1550 3366 1552
rect 3382 1556 3390 1558
rect 3382 1552 3384 1556
rect 3388 1552 3390 1556
rect 3382 1550 3390 1552
rect 3406 1556 3414 1558
rect 3406 1552 3408 1556
rect 3412 1552 3414 1556
rect 3406 1550 3414 1552
rect 3430 1556 3438 1558
rect 3430 1552 3432 1556
rect 3436 1552 3438 1556
rect 3430 1550 3438 1552
rect 3454 1556 3462 1558
rect 3454 1552 3456 1556
rect 3460 1552 3462 1556
rect 3454 1550 3462 1552
rect 3478 1556 3486 1558
rect 3478 1552 3480 1556
rect 3484 1552 3486 1556
rect 3478 1550 3486 1552
rect 3502 1556 3510 1558
rect 3502 1552 3504 1556
rect 3508 1552 3510 1556
rect 3502 1550 3510 1552
rect 3526 1556 3534 1558
rect 3526 1552 3528 1556
rect 3532 1552 3534 1556
rect 3526 1550 3534 1552
rect 3550 1556 3558 1558
rect 3550 1552 3552 1556
rect 3556 1552 3558 1556
rect 3550 1550 3558 1552
rect 3574 1556 3582 1558
rect 3574 1552 3576 1556
rect 3580 1552 3582 1556
rect 3574 1550 3582 1552
rect 3598 1556 3606 1558
rect 3598 1552 3600 1556
rect 3604 1552 3606 1556
rect 3598 1550 3606 1552
rect 3622 1556 3630 1558
rect 3622 1552 3624 1556
rect 3628 1552 3630 1556
rect 3622 1550 3630 1552
rect 3646 1556 3654 1558
rect 3646 1552 3648 1556
rect 3652 1552 3654 1556
rect 3646 1550 3654 1552
rect 3670 1556 3678 1558
rect 3670 1552 3672 1556
rect 3676 1552 3678 1556
rect 3670 1550 3678 1552
rect 3694 1556 3702 1558
rect 3694 1552 3696 1556
rect 3700 1552 3702 1556
rect 3694 1550 3702 1552
rect 3910 1556 3918 1558
rect 3910 1552 3912 1556
rect 3916 1552 3918 1556
rect 3910 1550 3918 1552
rect 3934 1556 3942 1558
rect 3934 1552 3936 1556
rect 3940 1552 3942 1556
rect 3934 1550 3942 1552
rect 3958 1556 3966 1558
rect 3958 1552 3960 1556
rect 3964 1552 3966 1556
rect 3958 1550 3966 1552
rect 3982 1556 3990 1558
rect 3982 1552 3984 1556
rect 3988 1552 3990 1556
rect 3982 1550 3990 1552
rect 4006 1556 4014 1558
rect 4006 1552 4008 1556
rect 4012 1552 4014 1556
rect 4006 1550 4014 1552
rect 4030 1556 4038 1558
rect 4030 1552 4032 1556
rect 4036 1552 4038 1556
rect 4030 1550 4038 1552
rect 4054 1556 4062 1558
rect 4054 1552 4056 1556
rect 4060 1552 4062 1556
rect 4054 1550 4062 1552
rect 4078 1556 4086 1558
rect 4078 1552 4080 1556
rect 4084 1552 4086 1556
rect 4078 1550 4086 1552
rect 4102 1556 4110 1558
rect 4102 1552 4104 1556
rect 4108 1552 4110 1556
rect 4102 1550 4110 1552
rect 4126 1556 4134 1558
rect 4126 1552 4128 1556
rect 4132 1552 4134 1556
rect 4126 1550 4134 1552
rect 4150 1556 4158 1558
rect 4150 1552 4152 1556
rect 4156 1552 4158 1556
rect 4150 1550 4158 1552
rect 4174 1556 4182 1558
rect 4174 1552 4176 1556
rect 4180 1552 4182 1556
rect 4174 1550 4182 1552
rect 4198 1556 4206 1558
rect 4198 1552 4200 1556
rect 4204 1552 4206 1556
rect 4198 1550 4206 1552
rect 4222 1556 4230 1558
rect 4222 1552 4224 1556
rect 4228 1552 4230 1556
rect 4222 1550 4230 1552
rect 4246 1556 4254 1558
rect 4246 1552 4248 1556
rect 4252 1552 4254 1556
rect 4246 1550 4254 1552
rect 4270 1556 4278 1558
rect 4270 1552 4272 1556
rect 4276 1552 4278 1556
rect 4270 1550 4278 1552
rect 4294 1556 4302 1558
rect 4294 1552 4296 1556
rect 4300 1552 4302 1556
rect 4294 1550 4302 1552
rect 4510 1556 4518 1558
rect 4510 1552 4512 1556
rect 4516 1552 4518 1556
rect 4510 1550 4518 1552
rect 4534 1556 4542 1558
rect 4534 1552 4536 1556
rect 4540 1552 4542 1556
rect 4534 1550 4542 1552
rect 4558 1556 4566 1558
rect 4558 1552 4560 1556
rect 4564 1552 4566 1556
rect 4558 1550 4566 1552
rect 4582 1556 4590 1558
rect 4582 1552 4584 1556
rect 4588 1552 4590 1556
rect 4582 1550 4590 1552
rect 4606 1556 4614 1558
rect 4606 1552 4608 1556
rect 4612 1552 4614 1556
rect 4606 1550 4614 1552
rect 4630 1556 4638 1558
rect 4630 1552 4632 1556
rect 4636 1552 4638 1556
rect 4630 1550 4638 1552
rect 4654 1556 4662 1558
rect 4654 1552 4656 1556
rect 4660 1552 4662 1556
rect 4654 1550 4662 1552
rect 4678 1556 4686 1558
rect 4678 1552 4680 1556
rect 4684 1552 4686 1556
rect 4678 1550 4686 1552
rect 4702 1556 4710 1558
rect 4702 1552 4704 1556
rect 4708 1552 4710 1556
rect 4702 1550 4710 1552
rect 4726 1556 4734 1558
rect 4726 1552 4728 1556
rect 4732 1552 4734 1556
rect 4726 1550 4734 1552
rect 4750 1556 4758 1558
rect 4750 1552 4752 1556
rect 4756 1552 4758 1556
rect 4750 1550 4758 1552
rect 4774 1556 4782 1558
rect 4774 1552 4776 1556
rect 4780 1552 4782 1556
rect 4774 1550 4782 1552
rect 4798 1556 4806 1558
rect 4798 1552 4800 1556
rect 4804 1552 4806 1556
rect 4798 1550 4806 1552
rect 4822 1556 4830 1558
rect 4822 1552 4824 1556
rect 4828 1552 4830 1556
rect 4822 1550 4830 1552
rect 4846 1556 4854 1558
rect 4846 1552 4848 1556
rect 4852 1552 4854 1556
rect 4846 1550 4854 1552
rect 4870 1556 4878 1558
rect 4870 1552 4872 1556
rect 4876 1552 4878 1556
rect 4870 1550 4878 1552
rect 4894 1556 4902 1558
rect 4894 1552 4896 1556
rect 4900 1552 4902 1556
rect 4894 1550 4902 1552
rect 5710 1556 5718 1558
rect 5710 1552 5712 1556
rect 5716 1552 5718 1556
rect 5710 1550 5718 1552
rect 5734 1556 5742 1558
rect 5734 1552 5736 1556
rect 5740 1552 5742 1556
rect 5734 1550 5742 1552
rect 5758 1556 5766 1558
rect 5758 1552 5760 1556
rect 5764 1552 5766 1556
rect 5758 1550 5766 1552
rect 5782 1556 5790 1558
rect 5782 1552 5784 1556
rect 5788 1552 5790 1556
rect 5782 1550 5790 1552
rect 5806 1556 5814 1558
rect 5806 1552 5808 1556
rect 5812 1552 5814 1556
rect 5806 1550 5814 1552
rect 5830 1556 5838 1558
rect 5830 1552 5832 1556
rect 5836 1552 5838 1556
rect 5830 1550 5838 1552
rect 5854 1556 5862 1558
rect 5854 1552 5856 1556
rect 5860 1552 5862 1556
rect 5854 1550 5862 1552
rect 5878 1556 5886 1558
rect 5878 1552 5880 1556
rect 5884 1552 5886 1556
rect 5878 1550 5886 1552
rect 5902 1556 5910 1558
rect 5902 1552 5904 1556
rect 5908 1552 5910 1556
rect 5902 1550 5910 1552
rect 5926 1556 5934 1558
rect 5926 1552 5928 1556
rect 5932 1552 5934 1556
rect 5926 1550 5934 1552
rect 5950 1556 5958 1558
rect 5950 1552 5952 1556
rect 5956 1552 5958 1556
rect 5950 1550 5958 1552
rect 5974 1556 5982 1558
rect 5974 1552 5976 1556
rect 5980 1552 5982 1556
rect 5974 1550 5982 1552
rect 5998 1556 6006 1558
rect 5998 1552 6000 1556
rect 6004 1552 6006 1556
rect 5998 1550 6006 1552
rect 6022 1556 6030 1558
rect 6022 1552 6024 1556
rect 6028 1552 6030 1556
rect 6022 1550 6030 1552
rect 6046 1556 6054 1558
rect 6046 1552 6048 1556
rect 6052 1552 6054 1556
rect 6046 1550 6054 1552
rect 6070 1556 6078 1558
rect 6070 1552 6072 1556
rect 6076 1552 6078 1556
rect 6070 1550 6078 1552
rect 6094 1556 6102 1558
rect 6094 1552 6096 1556
rect 6100 1552 6102 1556
rect 6094 1550 6102 1552
rect 6310 1556 6318 1558
rect 6310 1552 6312 1556
rect 6316 1552 6318 1556
rect 6310 1550 6318 1552
rect 6334 1556 6342 1558
rect 6334 1552 6336 1556
rect 6340 1552 6342 1556
rect 6334 1550 6342 1552
rect 6358 1556 6366 1558
rect 6358 1552 6360 1556
rect 6364 1552 6366 1556
rect 6358 1550 6366 1552
rect 6382 1556 6390 1558
rect 6382 1552 6384 1556
rect 6388 1552 6390 1556
rect 6382 1550 6390 1552
rect 6406 1556 6414 1558
rect 6406 1552 6408 1556
rect 6412 1552 6414 1556
rect 6406 1550 6414 1552
rect 6430 1556 6438 1558
rect 6430 1552 6432 1556
rect 6436 1552 6438 1556
rect 6430 1550 6438 1552
rect 6454 1556 6462 1558
rect 6454 1552 6456 1556
rect 6460 1552 6462 1556
rect 6454 1550 6462 1552
rect 6478 1556 6486 1558
rect 6478 1552 6480 1556
rect 6484 1552 6486 1556
rect 6478 1550 6486 1552
rect 6502 1556 6510 1558
rect 6502 1552 6504 1556
rect 6508 1552 6510 1556
rect 6502 1550 6510 1552
rect 6526 1556 6534 1558
rect 6526 1552 6528 1556
rect 6532 1552 6534 1556
rect 6526 1550 6534 1552
rect 6550 1556 6558 1558
rect 6550 1552 6552 1556
rect 6556 1552 6558 1556
rect 6550 1550 6558 1552
rect 6574 1556 6582 1558
rect 6574 1552 6576 1556
rect 6580 1552 6582 1556
rect 6574 1550 6582 1552
rect 6598 1556 6606 1558
rect 6598 1552 6600 1556
rect 6604 1552 6606 1556
rect 6598 1550 6606 1552
rect 6622 1556 6630 1558
rect 6622 1552 6624 1556
rect 6628 1552 6630 1556
rect 6622 1550 6630 1552
rect 6646 1556 6654 1558
rect 6646 1552 6648 1556
rect 6652 1552 6654 1556
rect 6646 1550 6654 1552
rect 6670 1556 6678 1558
rect 6670 1552 6672 1556
rect 6676 1552 6678 1556
rect 6670 1550 6678 1552
rect 6694 1556 6702 1558
rect 6694 1552 6696 1556
rect 6700 1552 6702 1556
rect 6694 1550 6702 1552
rect 6910 1556 6918 1558
rect 6910 1552 6912 1556
rect 6916 1552 6918 1556
rect 6910 1550 6918 1552
rect 6934 1556 6942 1558
rect 6934 1552 6936 1556
rect 6940 1552 6942 1556
rect 6934 1550 6942 1552
rect 6958 1556 6966 1558
rect 6958 1552 6960 1556
rect 6964 1552 6966 1556
rect 6958 1550 6966 1552
rect 6982 1556 6990 1558
rect 6982 1552 6984 1556
rect 6988 1552 6990 1556
rect 6982 1550 6990 1552
rect 7006 1556 7014 1558
rect 7006 1552 7008 1556
rect 7012 1552 7014 1556
rect 7006 1550 7014 1552
rect 7030 1556 7038 1558
rect 7030 1552 7032 1556
rect 7036 1552 7038 1556
rect 7030 1550 7038 1552
rect 7054 1556 7062 1558
rect 7054 1552 7056 1556
rect 7060 1552 7062 1556
rect 7054 1550 7062 1552
rect 7078 1556 7086 1558
rect 7078 1552 7080 1556
rect 7084 1552 7086 1556
rect 7078 1550 7086 1552
rect 7102 1556 7110 1558
rect 7102 1552 7104 1556
rect 7108 1552 7110 1556
rect 7102 1550 7110 1552
rect 7126 1556 7134 1558
rect 7126 1552 7128 1556
rect 7132 1552 7134 1556
rect 7126 1550 7134 1552
rect 7150 1556 7158 1558
rect 7150 1552 7152 1556
rect 7156 1552 7158 1556
rect 7150 1550 7158 1552
rect 7174 1556 7182 1558
rect 7174 1552 7176 1556
rect 7180 1552 7182 1556
rect 7174 1550 7182 1552
rect 7198 1550 7200 1558
rect 2098 1544 2106 1546
rect 2098 1540 2100 1544
rect 2104 1540 2106 1544
rect 2098 1538 2106 1540
rect 2122 1544 2130 1546
rect 2122 1540 2124 1544
rect 2128 1540 2130 1544
rect 2122 1538 2130 1540
rect 2146 1544 2154 1546
rect 2146 1540 2148 1544
rect 2152 1540 2154 1544
rect 2146 1538 2154 1540
rect 2170 1544 2178 1546
rect 2170 1540 2172 1544
rect 2176 1540 2178 1544
rect 2170 1538 2178 1540
rect 2194 1544 2202 1546
rect 2194 1540 2196 1544
rect 2200 1540 2202 1544
rect 2194 1538 2202 1540
rect 2218 1544 2226 1546
rect 2218 1540 2220 1544
rect 2224 1540 2226 1544
rect 2218 1538 2226 1540
rect 2242 1544 2250 1546
rect 2242 1540 2244 1544
rect 2248 1540 2250 1544
rect 2242 1538 2250 1540
rect 2266 1544 2274 1546
rect 2266 1540 2268 1544
rect 2272 1540 2274 1544
rect 2266 1538 2274 1540
rect 2290 1544 2298 1546
rect 2290 1540 2292 1544
rect 2296 1540 2298 1544
rect 2290 1538 2298 1540
rect 2314 1544 2322 1546
rect 2314 1540 2316 1544
rect 2320 1540 2322 1544
rect 2314 1538 2322 1540
rect 2338 1544 2346 1546
rect 2338 1540 2340 1544
rect 2344 1540 2346 1544
rect 2338 1538 2346 1540
rect 2362 1544 2370 1546
rect 2362 1540 2364 1544
rect 2368 1540 2370 1544
rect 2362 1538 2370 1540
rect 2386 1544 2394 1546
rect 2386 1540 2388 1544
rect 2392 1540 2394 1544
rect 2386 1538 2394 1540
rect 2410 1544 2418 1546
rect 2410 1540 2412 1544
rect 2416 1540 2418 1544
rect 2410 1538 2418 1540
rect 2434 1544 2442 1546
rect 2434 1540 2436 1544
rect 2440 1540 2442 1544
rect 2434 1538 2442 1540
rect 2458 1544 2466 1546
rect 2458 1540 2460 1544
rect 2464 1540 2466 1544
rect 2458 1538 2466 1540
rect 2482 1544 2490 1546
rect 2482 1540 2484 1544
rect 2488 1540 2490 1544
rect 2482 1538 2490 1540
rect 2698 1544 2706 1546
rect 2698 1540 2700 1544
rect 2704 1540 2706 1544
rect 2698 1538 2706 1540
rect 2722 1544 2730 1546
rect 2722 1540 2724 1544
rect 2728 1540 2730 1544
rect 2722 1538 2730 1540
rect 2746 1544 2754 1546
rect 2746 1540 2748 1544
rect 2752 1540 2754 1544
rect 2746 1538 2754 1540
rect 2770 1544 2778 1546
rect 2770 1540 2772 1544
rect 2776 1540 2778 1544
rect 2770 1538 2778 1540
rect 2794 1544 2802 1546
rect 2794 1540 2796 1544
rect 2800 1540 2802 1544
rect 2794 1538 2802 1540
rect 2818 1544 2826 1546
rect 2818 1540 2820 1544
rect 2824 1540 2826 1544
rect 2818 1538 2826 1540
rect 2842 1544 2850 1546
rect 2842 1540 2844 1544
rect 2848 1540 2850 1544
rect 2842 1538 2850 1540
rect 2866 1544 2874 1546
rect 2866 1540 2868 1544
rect 2872 1540 2874 1544
rect 2866 1538 2874 1540
rect 2890 1544 2898 1546
rect 2890 1540 2892 1544
rect 2896 1540 2898 1544
rect 2890 1538 2898 1540
rect 2914 1544 2922 1546
rect 2914 1540 2916 1544
rect 2920 1540 2922 1544
rect 2914 1538 2922 1540
rect 2938 1544 2946 1546
rect 2938 1540 2940 1544
rect 2944 1540 2946 1544
rect 2938 1538 2946 1540
rect 2962 1544 2970 1546
rect 2962 1540 2964 1544
rect 2968 1540 2970 1544
rect 2962 1538 2970 1540
rect 2986 1544 2994 1546
rect 2986 1540 2988 1544
rect 2992 1540 2994 1544
rect 2986 1538 2994 1540
rect 3010 1544 3018 1546
rect 3010 1540 3012 1544
rect 3016 1540 3018 1544
rect 3010 1538 3018 1540
rect 3034 1544 3042 1546
rect 3034 1540 3036 1544
rect 3040 1540 3042 1544
rect 3034 1538 3042 1540
rect 3058 1544 3066 1546
rect 3058 1540 3060 1544
rect 3064 1540 3066 1544
rect 3058 1538 3066 1540
rect 3082 1544 3090 1546
rect 3082 1540 3084 1544
rect 3088 1540 3090 1544
rect 3082 1538 3090 1540
rect 3298 1544 3306 1546
rect 3298 1540 3300 1544
rect 3304 1540 3306 1544
rect 3298 1538 3306 1540
rect 3322 1544 3330 1546
rect 3322 1540 3324 1544
rect 3328 1540 3330 1544
rect 3322 1538 3330 1540
rect 3346 1544 3354 1546
rect 3346 1540 3348 1544
rect 3352 1540 3354 1544
rect 3346 1538 3354 1540
rect 3370 1544 3378 1546
rect 3370 1540 3372 1544
rect 3376 1540 3378 1544
rect 3370 1538 3378 1540
rect 3394 1544 3402 1546
rect 3394 1540 3396 1544
rect 3400 1540 3402 1544
rect 3394 1538 3402 1540
rect 3418 1544 3426 1546
rect 3418 1540 3420 1544
rect 3424 1540 3426 1544
rect 3418 1538 3426 1540
rect 3442 1544 3450 1546
rect 3442 1540 3444 1544
rect 3448 1540 3450 1544
rect 3442 1538 3450 1540
rect 3466 1544 3474 1546
rect 3466 1540 3468 1544
rect 3472 1540 3474 1544
rect 3466 1538 3474 1540
rect 3490 1544 3498 1546
rect 3490 1540 3492 1544
rect 3496 1540 3498 1544
rect 3490 1538 3498 1540
rect 3514 1544 3522 1546
rect 3514 1540 3516 1544
rect 3520 1540 3522 1544
rect 3514 1538 3522 1540
rect 3538 1544 3546 1546
rect 3538 1540 3540 1544
rect 3544 1540 3546 1544
rect 3538 1538 3546 1540
rect 3562 1544 3570 1546
rect 3562 1540 3564 1544
rect 3568 1540 3570 1544
rect 3562 1538 3570 1540
rect 3586 1544 3594 1546
rect 3586 1540 3588 1544
rect 3592 1540 3594 1544
rect 3586 1538 3594 1540
rect 3610 1544 3618 1546
rect 3610 1540 3612 1544
rect 3616 1540 3618 1544
rect 3610 1538 3618 1540
rect 3634 1544 3642 1546
rect 3634 1540 3636 1544
rect 3640 1540 3642 1544
rect 3634 1538 3642 1540
rect 3658 1544 3666 1546
rect 3658 1540 3660 1544
rect 3664 1540 3666 1544
rect 3658 1538 3666 1540
rect 3682 1544 3690 1546
rect 3682 1540 3684 1544
rect 3688 1540 3690 1544
rect 3682 1538 3690 1540
rect 3898 1544 3906 1546
rect 3898 1540 3900 1544
rect 3904 1540 3906 1544
rect 3898 1538 3906 1540
rect 3922 1544 3930 1546
rect 3922 1540 3924 1544
rect 3928 1540 3930 1544
rect 3922 1538 3930 1540
rect 3946 1544 3954 1546
rect 3946 1540 3948 1544
rect 3952 1540 3954 1544
rect 3946 1538 3954 1540
rect 3970 1544 3978 1546
rect 3970 1540 3972 1544
rect 3976 1540 3978 1544
rect 3970 1538 3978 1540
rect 3994 1544 4002 1546
rect 3994 1540 3996 1544
rect 4000 1540 4002 1544
rect 3994 1538 4002 1540
rect 4018 1544 4026 1546
rect 4018 1540 4020 1544
rect 4024 1540 4026 1544
rect 4018 1538 4026 1540
rect 4042 1544 4050 1546
rect 4042 1540 4044 1544
rect 4048 1540 4050 1544
rect 4042 1538 4050 1540
rect 4066 1544 4074 1546
rect 4066 1540 4068 1544
rect 4072 1540 4074 1544
rect 4066 1538 4074 1540
rect 4090 1544 4098 1546
rect 4090 1540 4092 1544
rect 4096 1540 4098 1544
rect 4090 1538 4098 1540
rect 4114 1544 4122 1546
rect 4114 1540 4116 1544
rect 4120 1540 4122 1544
rect 4114 1538 4122 1540
rect 4138 1544 4146 1546
rect 4138 1540 4140 1544
rect 4144 1540 4146 1544
rect 4138 1538 4146 1540
rect 4162 1544 4170 1546
rect 4162 1540 4164 1544
rect 4168 1540 4170 1544
rect 4162 1538 4170 1540
rect 4186 1544 4194 1546
rect 4186 1540 4188 1544
rect 4192 1540 4194 1544
rect 4186 1538 4194 1540
rect 4210 1544 4218 1546
rect 4210 1540 4212 1544
rect 4216 1540 4218 1544
rect 4210 1538 4218 1540
rect 4234 1544 4242 1546
rect 4234 1540 4236 1544
rect 4240 1540 4242 1544
rect 4234 1538 4242 1540
rect 4258 1544 4266 1546
rect 4258 1540 4260 1544
rect 4264 1540 4266 1544
rect 4258 1538 4266 1540
rect 4282 1544 4290 1546
rect 4282 1540 4284 1544
rect 4288 1540 4290 1544
rect 4282 1538 4290 1540
rect 4498 1544 4506 1546
rect 4498 1540 4500 1544
rect 4504 1540 4506 1544
rect 4498 1538 4506 1540
rect 4522 1544 4530 1546
rect 4522 1540 4524 1544
rect 4528 1540 4530 1544
rect 4522 1538 4530 1540
rect 4546 1544 4554 1546
rect 4546 1540 4548 1544
rect 4552 1540 4554 1544
rect 4546 1538 4554 1540
rect 4570 1544 4578 1546
rect 4570 1540 4572 1544
rect 4576 1540 4578 1544
rect 4570 1538 4578 1540
rect 4594 1544 4602 1546
rect 4594 1540 4596 1544
rect 4600 1540 4602 1544
rect 4594 1538 4602 1540
rect 4618 1544 4626 1546
rect 4618 1540 4620 1544
rect 4624 1540 4626 1544
rect 4618 1538 4626 1540
rect 4642 1544 4650 1546
rect 4642 1540 4644 1544
rect 4648 1540 4650 1544
rect 4642 1538 4650 1540
rect 4666 1544 4674 1546
rect 4666 1540 4668 1544
rect 4672 1540 4674 1544
rect 4666 1538 4674 1540
rect 4690 1544 4698 1546
rect 4690 1540 4692 1544
rect 4696 1540 4698 1544
rect 4690 1538 4698 1540
rect 4714 1544 4722 1546
rect 4714 1540 4716 1544
rect 4720 1540 4722 1544
rect 4714 1538 4722 1540
rect 4738 1544 4746 1546
rect 4738 1540 4740 1544
rect 4744 1540 4746 1544
rect 4738 1538 4746 1540
rect 4762 1544 4770 1546
rect 4762 1540 4764 1544
rect 4768 1540 4770 1544
rect 4762 1538 4770 1540
rect 4786 1544 4794 1546
rect 4786 1540 4788 1544
rect 4792 1540 4794 1544
rect 4786 1538 4794 1540
rect 4810 1544 4818 1546
rect 4810 1540 4812 1544
rect 4816 1540 4818 1544
rect 4810 1538 4818 1540
rect 4834 1544 4842 1546
rect 4834 1540 4836 1544
rect 4840 1540 4842 1544
rect 4834 1538 4842 1540
rect 4858 1544 4866 1546
rect 4858 1540 4860 1544
rect 4864 1540 4866 1544
rect 4858 1538 4866 1540
rect 4882 1544 4890 1546
rect 4882 1540 4884 1544
rect 4888 1540 4890 1544
rect 4882 1538 4890 1540
rect 5698 1544 5706 1546
rect 5698 1540 5700 1544
rect 5704 1540 5706 1544
rect 5698 1538 5706 1540
rect 5722 1544 5730 1546
rect 5722 1540 5724 1544
rect 5728 1540 5730 1544
rect 5722 1538 5730 1540
rect 5746 1544 5754 1546
rect 5746 1540 5748 1544
rect 5752 1540 5754 1544
rect 5746 1538 5754 1540
rect 5770 1544 5778 1546
rect 5770 1540 5772 1544
rect 5776 1540 5778 1544
rect 5770 1538 5778 1540
rect 5794 1544 5802 1546
rect 5794 1540 5796 1544
rect 5800 1540 5802 1544
rect 5794 1538 5802 1540
rect 5818 1544 5826 1546
rect 5818 1540 5820 1544
rect 5824 1540 5826 1544
rect 5818 1538 5826 1540
rect 5842 1544 5850 1546
rect 5842 1540 5844 1544
rect 5848 1540 5850 1544
rect 5842 1538 5850 1540
rect 5866 1544 5874 1546
rect 5866 1540 5868 1544
rect 5872 1540 5874 1544
rect 5866 1538 5874 1540
rect 5890 1544 5898 1546
rect 5890 1540 5892 1544
rect 5896 1540 5898 1544
rect 5890 1538 5898 1540
rect 5914 1544 5922 1546
rect 5914 1540 5916 1544
rect 5920 1540 5922 1544
rect 5914 1538 5922 1540
rect 5938 1544 5946 1546
rect 5938 1540 5940 1544
rect 5944 1540 5946 1544
rect 5938 1538 5946 1540
rect 5962 1544 5970 1546
rect 5962 1540 5964 1544
rect 5968 1540 5970 1544
rect 5962 1538 5970 1540
rect 5986 1544 5994 1546
rect 5986 1540 5988 1544
rect 5992 1540 5994 1544
rect 5986 1538 5994 1540
rect 6010 1544 6018 1546
rect 6010 1540 6012 1544
rect 6016 1540 6018 1544
rect 6010 1538 6018 1540
rect 6034 1544 6042 1546
rect 6034 1540 6036 1544
rect 6040 1540 6042 1544
rect 6034 1538 6042 1540
rect 6058 1544 6066 1546
rect 6058 1540 6060 1544
rect 6064 1540 6066 1544
rect 6058 1538 6066 1540
rect 6082 1544 6090 1546
rect 6082 1540 6084 1544
rect 6088 1540 6090 1544
rect 6082 1538 6090 1540
rect 6298 1544 6306 1546
rect 6298 1540 6300 1544
rect 6304 1540 6306 1544
rect 6298 1538 6306 1540
rect 6322 1544 6330 1546
rect 6322 1540 6324 1544
rect 6328 1540 6330 1544
rect 6322 1538 6330 1540
rect 6346 1544 6354 1546
rect 6346 1540 6348 1544
rect 6352 1540 6354 1544
rect 6346 1538 6354 1540
rect 6370 1544 6378 1546
rect 6370 1540 6372 1544
rect 6376 1540 6378 1544
rect 6370 1538 6378 1540
rect 6394 1544 6402 1546
rect 6394 1540 6396 1544
rect 6400 1540 6402 1544
rect 6394 1538 6402 1540
rect 6418 1544 6426 1546
rect 6418 1540 6420 1544
rect 6424 1540 6426 1544
rect 6418 1538 6426 1540
rect 6442 1544 6450 1546
rect 6442 1540 6444 1544
rect 6448 1540 6450 1544
rect 6442 1538 6450 1540
rect 6466 1544 6474 1546
rect 6466 1540 6468 1544
rect 6472 1540 6474 1544
rect 6466 1538 6474 1540
rect 6490 1544 6498 1546
rect 6490 1540 6492 1544
rect 6496 1540 6498 1544
rect 6490 1538 6498 1540
rect 6514 1544 6522 1546
rect 6514 1540 6516 1544
rect 6520 1540 6522 1544
rect 6514 1538 6522 1540
rect 6538 1544 6546 1546
rect 6538 1540 6540 1544
rect 6544 1540 6546 1544
rect 6538 1538 6546 1540
rect 6562 1544 6570 1546
rect 6562 1540 6564 1544
rect 6568 1540 6570 1544
rect 6562 1538 6570 1540
rect 6586 1544 6594 1546
rect 6586 1540 6588 1544
rect 6592 1540 6594 1544
rect 6586 1538 6594 1540
rect 6610 1544 6618 1546
rect 6610 1540 6612 1544
rect 6616 1540 6618 1544
rect 6610 1538 6618 1540
rect 6634 1544 6642 1546
rect 6634 1540 6636 1544
rect 6640 1540 6642 1544
rect 6634 1538 6642 1540
rect 6658 1544 6666 1546
rect 6658 1540 6660 1544
rect 6664 1540 6666 1544
rect 6658 1538 6666 1540
rect 6682 1544 6690 1546
rect 6682 1540 6684 1544
rect 6688 1540 6690 1544
rect 6682 1538 6690 1540
rect 6898 1544 6906 1546
rect 6898 1540 6900 1544
rect 6904 1540 6906 1544
rect 6898 1538 6906 1540
rect 6922 1544 6930 1546
rect 6922 1540 6924 1544
rect 6928 1540 6930 1544
rect 6922 1538 6930 1540
rect 6946 1544 6954 1546
rect 6946 1540 6948 1544
rect 6952 1540 6954 1544
rect 6946 1538 6954 1540
rect 6970 1544 6978 1546
rect 6970 1540 6972 1544
rect 6976 1540 6978 1544
rect 6970 1538 6978 1540
rect 6994 1544 7002 1546
rect 6994 1540 6996 1544
rect 7000 1540 7002 1544
rect 6994 1538 7002 1540
rect 7018 1544 7026 1546
rect 7018 1540 7020 1544
rect 7024 1540 7026 1544
rect 7018 1538 7026 1540
rect 7042 1544 7050 1546
rect 7042 1540 7044 1544
rect 7048 1540 7050 1544
rect 7042 1538 7050 1540
rect 7066 1544 7074 1546
rect 7066 1540 7068 1544
rect 7072 1540 7074 1544
rect 7066 1538 7074 1540
rect 7090 1544 7098 1546
rect 7090 1540 7092 1544
rect 7096 1540 7098 1544
rect 7090 1538 7098 1540
rect 7114 1544 7122 1546
rect 7114 1540 7116 1544
rect 7120 1540 7122 1544
rect 7114 1538 7122 1540
rect 7138 1544 7146 1546
rect 7138 1540 7140 1544
rect 7144 1540 7146 1544
rect 7138 1538 7146 1540
rect 7162 1544 7170 1546
rect 7162 1540 7164 1544
rect 7168 1540 7170 1544
rect 7162 1538 7170 1540
rect 7186 1544 7194 1546
rect 7186 1540 7188 1544
rect 7192 1540 7194 1544
rect 7186 1538 7194 1540
rect 4412 1328 4414 1330
rect 4986 1328 4988 1330
rect 5012 1328 5014 1330
rect 5586 1328 5588 1330
rect 4410 1326 4412 1328
rect 4988 1326 4990 1328
rect 5010 1326 5012 1328
rect 5588 1326 5590 1328
rect 2012 1316 2014 1324
rect 2020 1316 2022 1318
rect 2612 1316 2614 1324
rect 3220 1320 3222 1322
rect 3778 1320 3780 1322
rect 3820 1320 3822 1322
rect 4378 1320 4380 1322
rect 5620 1320 5622 1322
rect 6220 1320 6222 1322
rect 6778 1320 6780 1322
rect 3218 1318 3220 1320
rect 3780 1318 3782 1320
rect 3818 1318 3820 1320
rect 4380 1318 4382 1320
rect 5618 1318 5620 1320
rect 6218 1318 6220 1320
rect 6780 1318 6782 1320
rect 2620 1316 2622 1318
rect 6812 1316 6814 1324
rect 6820 1316 6822 1318
rect 2008 1314 2010 1316
rect 2014 1314 2016 1316
rect 2018 1314 2022 1316
rect 2608 1314 2610 1316
rect 2614 1314 2616 1316
rect 2618 1314 2622 1316
rect 6808 1314 6810 1316
rect 6814 1314 6816 1316
rect 6818 1314 6822 1316
rect 2010 1312 2014 1314
rect 2610 1312 2614 1314
rect 6810 1312 6814 1314
rect 2562 1302 2564 1304
rect 3162 1302 3164 1304
rect 2036 1300 2038 1302
rect 2564 1300 2566 1302
rect 2636 1300 2638 1302
rect 3164 1300 3166 1302
rect 6836 1300 6838 1302
rect 2034 1298 2036 1300
rect 2634 1298 2636 1300
rect 6834 1298 6836 1300
rect 3280 1296 3290 1298
rect 3278 1294 3290 1296
rect 3710 1296 3720 1298
rect 3880 1296 3890 1298
rect 3710 1294 3722 1296
rect 3878 1294 3890 1296
rect 4310 1296 4320 1298
rect 6280 1296 6290 1298
rect 4310 1294 4322 1296
rect 6278 1294 6290 1296
rect 6710 1296 6720 1298
rect 6710 1294 6722 1296
rect 3280 1290 3282 1294
rect 3718 1290 3720 1294
rect 3280 1286 3290 1290
rect 3278 1284 3290 1286
rect 3710 1286 3720 1290
rect 3880 1290 3882 1294
rect 4318 1290 4320 1294
rect 4474 1290 4476 1292
rect 4504 1290 4506 1292
rect 4534 1290 4536 1292
rect 4564 1290 4566 1292
rect 4594 1290 4596 1292
rect 4624 1290 4626 1292
rect 4654 1290 4656 1292
rect 4684 1290 4686 1292
rect 4714 1290 4716 1292
rect 4744 1290 4746 1292
rect 4774 1290 4776 1292
rect 4804 1290 4806 1292
rect 4834 1290 4836 1292
rect 4864 1290 4866 1292
rect 4894 1290 4896 1292
rect 4924 1290 4926 1292
rect 5074 1290 5076 1292
rect 5104 1290 5106 1292
rect 5134 1290 5136 1292
rect 5164 1290 5166 1292
rect 5194 1290 5196 1292
rect 5224 1290 5226 1292
rect 5254 1290 5256 1292
rect 5284 1290 5286 1292
rect 5314 1290 5316 1292
rect 5344 1290 5346 1292
rect 5374 1290 5376 1292
rect 5404 1290 5406 1292
rect 5434 1290 5436 1292
rect 5464 1290 5466 1292
rect 5494 1290 5496 1292
rect 5524 1290 5526 1292
rect 5674 1290 5676 1292
rect 5704 1290 5706 1292
rect 5734 1290 5736 1292
rect 5764 1290 5766 1292
rect 5794 1290 5796 1292
rect 5824 1290 5826 1292
rect 5854 1290 5856 1292
rect 5884 1290 5886 1292
rect 5914 1290 5916 1292
rect 5944 1290 5946 1292
rect 5974 1290 5976 1292
rect 6004 1290 6006 1292
rect 6034 1290 6036 1292
rect 6064 1290 6066 1292
rect 6094 1290 6096 1292
rect 6124 1290 6126 1292
rect 6280 1290 6282 1294
rect 6718 1290 6720 1294
rect 3880 1286 3890 1290
rect 3710 1284 3722 1286
rect 3878 1284 3890 1286
rect 4310 1286 4320 1290
rect 4476 1288 4478 1290
rect 4482 1288 4484 1290
rect 4506 1288 4508 1290
rect 4512 1288 4514 1290
rect 4536 1288 4538 1290
rect 4542 1288 4544 1290
rect 4566 1288 4568 1290
rect 4572 1288 4574 1290
rect 4596 1288 4598 1290
rect 4602 1288 4604 1290
rect 4626 1288 4628 1290
rect 4632 1288 4634 1290
rect 4656 1288 4658 1290
rect 4662 1288 4664 1290
rect 4686 1288 4688 1290
rect 4692 1288 4694 1290
rect 4716 1288 4718 1290
rect 4722 1288 4724 1290
rect 4746 1288 4748 1290
rect 4752 1288 4754 1290
rect 4776 1288 4778 1290
rect 4782 1288 4784 1290
rect 4806 1288 4808 1290
rect 4812 1288 4814 1290
rect 4836 1288 4838 1290
rect 4842 1288 4844 1290
rect 4866 1288 4868 1290
rect 4872 1288 4874 1290
rect 4896 1288 4898 1290
rect 4902 1288 4904 1290
rect 4926 1288 4928 1290
rect 4932 1288 4934 1290
rect 5076 1288 5078 1290
rect 5082 1288 5084 1290
rect 5106 1288 5108 1290
rect 5112 1288 5114 1290
rect 5136 1288 5138 1290
rect 5142 1288 5144 1290
rect 5166 1288 5168 1290
rect 5172 1288 5174 1290
rect 5196 1288 5198 1290
rect 5202 1288 5204 1290
rect 5226 1288 5228 1290
rect 5232 1288 5234 1290
rect 5256 1288 5258 1290
rect 5262 1288 5264 1290
rect 5286 1288 5288 1290
rect 5292 1288 5294 1290
rect 5316 1288 5318 1290
rect 5322 1288 5324 1290
rect 5346 1288 5348 1290
rect 5352 1288 5354 1290
rect 5376 1288 5378 1290
rect 5382 1288 5384 1290
rect 5406 1288 5408 1290
rect 5412 1288 5414 1290
rect 5436 1288 5438 1290
rect 5442 1288 5444 1290
rect 5466 1288 5468 1290
rect 5472 1288 5474 1290
rect 5496 1288 5498 1290
rect 5502 1288 5504 1290
rect 5526 1288 5528 1290
rect 5532 1288 5534 1290
rect 5676 1288 5678 1290
rect 5682 1288 5684 1290
rect 5706 1288 5708 1290
rect 5712 1288 5714 1290
rect 5736 1288 5738 1290
rect 5742 1288 5744 1290
rect 5766 1288 5768 1290
rect 5772 1288 5774 1290
rect 5796 1288 5798 1290
rect 5802 1288 5804 1290
rect 5826 1288 5828 1290
rect 5832 1288 5834 1290
rect 5856 1288 5858 1290
rect 5862 1288 5864 1290
rect 5886 1288 5888 1290
rect 5892 1288 5894 1290
rect 5916 1288 5918 1290
rect 5922 1288 5924 1290
rect 5946 1288 5948 1290
rect 5952 1288 5954 1290
rect 5976 1288 5978 1290
rect 5982 1288 5984 1290
rect 6006 1288 6008 1290
rect 6012 1288 6014 1290
rect 6036 1288 6038 1290
rect 6042 1288 6044 1290
rect 6066 1288 6068 1290
rect 6072 1288 6074 1290
rect 6096 1288 6098 1290
rect 6102 1288 6104 1290
rect 6126 1288 6128 1290
rect 6132 1288 6134 1290
rect 4484 1286 4486 1288
rect 4514 1286 4516 1288
rect 4544 1286 4546 1288
rect 4574 1286 4576 1288
rect 4604 1286 4606 1288
rect 4634 1286 4636 1288
rect 4664 1286 4666 1288
rect 4694 1286 4696 1288
rect 4724 1286 4726 1288
rect 4754 1286 4756 1288
rect 4784 1286 4786 1288
rect 4814 1286 4816 1288
rect 4844 1286 4846 1288
rect 4874 1286 4876 1288
rect 4904 1286 4906 1288
rect 4934 1286 4936 1288
rect 5084 1286 5086 1288
rect 5114 1286 5116 1288
rect 5144 1286 5146 1288
rect 5174 1286 5176 1288
rect 5204 1286 5206 1288
rect 5234 1286 5236 1288
rect 5264 1286 5266 1288
rect 5294 1286 5296 1288
rect 5324 1286 5326 1288
rect 5354 1286 5356 1288
rect 5384 1286 5386 1288
rect 5414 1286 5416 1288
rect 5444 1286 5446 1288
rect 5474 1286 5476 1288
rect 5504 1286 5506 1288
rect 5534 1286 5536 1288
rect 5684 1286 5686 1288
rect 5714 1286 5716 1288
rect 5744 1286 5746 1288
rect 5774 1286 5776 1288
rect 5804 1286 5806 1288
rect 5834 1286 5836 1288
rect 5864 1286 5866 1288
rect 5894 1286 5896 1288
rect 5924 1286 5926 1288
rect 5954 1286 5956 1288
rect 5984 1286 5986 1288
rect 6014 1286 6016 1288
rect 6044 1286 6046 1288
rect 6074 1286 6076 1288
rect 6104 1286 6106 1288
rect 6134 1286 6136 1288
rect 6280 1286 6290 1290
rect 4310 1284 4322 1286
rect 6278 1284 6290 1286
rect 6710 1286 6720 1290
rect 6710 1284 6722 1286
rect 2058 1282 2060 1284
rect 2658 1282 2660 1284
rect 3280 1282 3282 1284
rect 3718 1282 3720 1284
rect 3880 1282 3882 1284
rect 4318 1282 4320 1284
rect 6280 1282 6282 1284
rect 6718 1282 6720 1284
rect 6858 1282 6860 1284
rect 2060 1280 2062 1282
rect 2660 1280 2662 1282
rect 3282 1280 3284 1282
rect 3716 1280 3718 1282
rect 3882 1280 3884 1282
rect 4316 1280 4318 1282
rect 4484 1280 4486 1282
rect 4514 1280 4516 1282
rect 4544 1280 4546 1282
rect 4574 1280 4576 1282
rect 4604 1280 4606 1282
rect 4634 1280 4636 1282
rect 4664 1280 4666 1282
rect 4694 1280 4696 1282
rect 4724 1280 4726 1282
rect 4754 1280 4756 1282
rect 4784 1280 4786 1282
rect 4814 1280 4816 1282
rect 4844 1280 4846 1282
rect 4874 1280 4876 1282
rect 4904 1280 4906 1282
rect 4934 1280 4936 1282
rect 5084 1280 5086 1282
rect 5114 1280 5116 1282
rect 5144 1280 5146 1282
rect 5174 1280 5176 1282
rect 5204 1280 5206 1282
rect 5234 1280 5236 1282
rect 5264 1280 5266 1282
rect 5294 1280 5296 1282
rect 5324 1280 5326 1282
rect 5354 1280 5356 1282
rect 5384 1280 5386 1282
rect 5414 1280 5416 1282
rect 5444 1280 5446 1282
rect 5474 1280 5476 1282
rect 5504 1280 5506 1282
rect 5534 1280 5536 1282
rect 5684 1280 5686 1282
rect 5714 1280 5716 1282
rect 5744 1280 5746 1282
rect 5774 1280 5776 1282
rect 5804 1280 5806 1282
rect 5834 1280 5836 1282
rect 5864 1280 5866 1282
rect 5894 1280 5896 1282
rect 5924 1280 5926 1282
rect 5954 1280 5956 1282
rect 5984 1280 5986 1282
rect 6014 1280 6016 1282
rect 6044 1280 6046 1282
rect 6074 1280 6076 1282
rect 6104 1280 6106 1282
rect 6134 1280 6136 1282
rect 6282 1280 6284 1282
rect 6716 1280 6718 1282
rect 6860 1280 6862 1282
rect 3250 1279 3252 1280
rect 3748 1279 3750 1280
rect 3850 1279 3852 1280
rect 4348 1279 4350 1280
rect 4476 1278 4478 1280
rect 4482 1278 4484 1280
rect 4506 1278 4508 1280
rect 4512 1278 4514 1280
rect 4536 1278 4538 1280
rect 4542 1278 4544 1280
rect 4566 1278 4568 1280
rect 4572 1278 4574 1280
rect 4596 1278 4598 1280
rect 4602 1278 4604 1280
rect 4626 1278 4628 1280
rect 4632 1278 4634 1280
rect 4656 1278 4658 1280
rect 4662 1278 4664 1280
rect 4686 1278 4688 1280
rect 4692 1278 4694 1280
rect 4716 1278 4718 1280
rect 4722 1278 4724 1280
rect 4746 1278 4748 1280
rect 4752 1278 4754 1280
rect 4776 1278 4778 1280
rect 4782 1278 4784 1280
rect 4806 1278 4808 1280
rect 4812 1278 4814 1280
rect 4836 1278 4838 1280
rect 4842 1278 4844 1280
rect 4866 1278 4868 1280
rect 4872 1278 4874 1280
rect 4896 1278 4898 1280
rect 4902 1278 4904 1280
rect 4926 1278 4928 1280
rect 4932 1278 4934 1280
rect 5076 1278 5078 1280
rect 5082 1278 5084 1280
rect 5106 1278 5108 1280
rect 5112 1278 5114 1280
rect 5136 1278 5138 1280
rect 5142 1278 5144 1280
rect 5166 1278 5168 1280
rect 5172 1278 5174 1280
rect 5196 1278 5198 1280
rect 5202 1278 5204 1280
rect 5226 1278 5228 1280
rect 5232 1278 5234 1280
rect 5256 1278 5258 1280
rect 5262 1278 5264 1280
rect 5286 1278 5288 1280
rect 5292 1278 5294 1280
rect 5316 1278 5318 1280
rect 5322 1278 5324 1280
rect 5346 1278 5348 1280
rect 5352 1278 5354 1280
rect 5376 1278 5378 1280
rect 5382 1278 5384 1280
rect 5406 1278 5408 1280
rect 5412 1278 5414 1280
rect 5436 1278 5438 1280
rect 5442 1278 5444 1280
rect 5466 1278 5468 1280
rect 5472 1278 5474 1280
rect 5496 1278 5498 1280
rect 5502 1278 5504 1280
rect 5526 1278 5528 1280
rect 5532 1278 5534 1280
rect 5676 1278 5678 1280
rect 5682 1278 5684 1280
rect 5706 1278 5708 1280
rect 5712 1278 5714 1280
rect 5736 1278 5738 1280
rect 5742 1278 5744 1280
rect 5766 1278 5768 1280
rect 5772 1278 5774 1280
rect 5796 1278 5798 1280
rect 5802 1278 5804 1280
rect 5826 1278 5828 1280
rect 5832 1278 5834 1280
rect 5856 1278 5858 1280
rect 5862 1278 5864 1280
rect 5886 1278 5888 1280
rect 5892 1278 5894 1280
rect 5916 1278 5918 1280
rect 5922 1278 5924 1280
rect 5946 1278 5948 1280
rect 5952 1278 5954 1280
rect 5976 1278 5978 1280
rect 5982 1278 5984 1280
rect 6006 1278 6008 1280
rect 6012 1278 6014 1280
rect 6036 1278 6038 1280
rect 6042 1278 6044 1280
rect 6066 1278 6068 1280
rect 6072 1278 6074 1280
rect 6096 1278 6098 1280
rect 6102 1278 6104 1280
rect 6126 1278 6128 1280
rect 6132 1278 6134 1280
rect 6250 1279 6252 1280
rect 6748 1279 6750 1280
rect 3248 1277 3250 1278
rect 3750 1277 3752 1278
rect 3848 1277 3850 1278
rect 4350 1277 4352 1278
rect 4474 1276 4476 1278
rect 4504 1276 4506 1278
rect 4534 1276 4536 1278
rect 4564 1276 4566 1278
rect 4594 1276 4596 1278
rect 4624 1276 4626 1278
rect 4654 1276 4656 1278
rect 4684 1276 4686 1278
rect 4714 1276 4716 1278
rect 4744 1276 4746 1278
rect 4774 1276 4776 1278
rect 4804 1276 4806 1278
rect 4834 1276 4836 1278
rect 4864 1276 4866 1278
rect 4894 1276 4896 1278
rect 4924 1276 4926 1278
rect 5074 1276 5076 1278
rect 5104 1276 5106 1278
rect 5134 1276 5136 1278
rect 5164 1276 5166 1278
rect 5194 1276 5196 1278
rect 5224 1276 5226 1278
rect 5254 1276 5256 1278
rect 5284 1276 5286 1278
rect 5314 1276 5316 1278
rect 5344 1276 5346 1278
rect 5374 1276 5376 1278
rect 5404 1276 5406 1278
rect 5434 1276 5436 1278
rect 5464 1276 5466 1278
rect 5494 1276 5496 1278
rect 5524 1276 5526 1278
rect 5674 1276 5676 1278
rect 5704 1276 5706 1278
rect 5734 1276 5736 1278
rect 5764 1276 5766 1278
rect 5794 1276 5796 1278
rect 5824 1276 5826 1278
rect 5854 1276 5856 1278
rect 5884 1276 5886 1278
rect 5914 1276 5916 1278
rect 5944 1276 5946 1278
rect 5974 1276 5976 1278
rect 6004 1276 6006 1278
rect 6034 1276 6036 1278
rect 6064 1276 6066 1278
rect 6094 1276 6096 1278
rect 6124 1276 6126 1278
rect 6248 1277 6250 1278
rect 6750 1277 6752 1278
rect 4474 1270 4476 1272
rect 4504 1270 4506 1272
rect 4534 1270 4536 1272
rect 4564 1270 4566 1272
rect 4594 1270 4596 1272
rect 4624 1270 4626 1272
rect 4654 1270 4656 1272
rect 4684 1270 4686 1272
rect 4714 1270 4716 1272
rect 4744 1270 4746 1272
rect 4774 1270 4776 1272
rect 4804 1270 4806 1272
rect 4834 1270 4836 1272
rect 4864 1270 4866 1272
rect 4894 1270 4896 1272
rect 4924 1270 4926 1272
rect 5074 1270 5076 1272
rect 5104 1270 5106 1272
rect 5134 1270 5136 1272
rect 5164 1270 5166 1272
rect 5194 1270 5196 1272
rect 5224 1270 5226 1272
rect 5254 1270 5256 1272
rect 5284 1270 5286 1272
rect 5314 1270 5316 1272
rect 5344 1270 5346 1272
rect 5374 1270 5376 1272
rect 5404 1270 5406 1272
rect 5434 1270 5436 1272
rect 5464 1270 5466 1272
rect 5494 1270 5496 1272
rect 5524 1270 5526 1272
rect 5674 1270 5676 1272
rect 5704 1270 5706 1272
rect 5734 1270 5736 1272
rect 5764 1270 5766 1272
rect 5794 1270 5796 1272
rect 5824 1270 5826 1272
rect 5854 1270 5856 1272
rect 5884 1270 5886 1272
rect 5914 1270 5916 1272
rect 5944 1270 5946 1272
rect 5974 1270 5976 1272
rect 6004 1270 6006 1272
rect 6034 1270 6036 1272
rect 6064 1270 6066 1272
rect 6094 1270 6096 1272
rect 6124 1270 6126 1272
rect 4476 1268 4478 1270
rect 4482 1268 4484 1270
rect 4506 1268 4508 1270
rect 4512 1268 4514 1270
rect 4536 1268 4538 1270
rect 4542 1268 4544 1270
rect 4566 1268 4568 1270
rect 4572 1268 4574 1270
rect 4596 1268 4598 1270
rect 4602 1268 4604 1270
rect 4626 1268 4628 1270
rect 4632 1268 4634 1270
rect 4656 1268 4658 1270
rect 4662 1268 4664 1270
rect 4686 1268 4688 1270
rect 4692 1268 4694 1270
rect 4716 1268 4718 1270
rect 4722 1268 4724 1270
rect 4746 1268 4748 1270
rect 4752 1268 4754 1270
rect 4776 1268 4778 1270
rect 4782 1268 4784 1270
rect 4806 1268 4808 1270
rect 4812 1268 4814 1270
rect 4836 1268 4838 1270
rect 4842 1268 4844 1270
rect 4866 1268 4868 1270
rect 4872 1268 4874 1270
rect 4896 1268 4898 1270
rect 4902 1268 4904 1270
rect 4926 1268 4928 1270
rect 4932 1268 4934 1270
rect 5076 1268 5078 1270
rect 5082 1268 5084 1270
rect 5106 1268 5108 1270
rect 5112 1268 5114 1270
rect 5136 1268 5138 1270
rect 5142 1268 5144 1270
rect 5166 1268 5168 1270
rect 5172 1268 5174 1270
rect 5196 1268 5198 1270
rect 5202 1268 5204 1270
rect 5226 1268 5228 1270
rect 5232 1268 5234 1270
rect 5256 1268 5258 1270
rect 5262 1268 5264 1270
rect 5286 1268 5288 1270
rect 5292 1268 5294 1270
rect 5316 1268 5318 1270
rect 5322 1268 5324 1270
rect 5346 1268 5348 1270
rect 5352 1268 5354 1270
rect 5376 1268 5378 1270
rect 5382 1268 5384 1270
rect 5406 1268 5408 1270
rect 5412 1268 5414 1270
rect 5436 1268 5438 1270
rect 5442 1268 5444 1270
rect 5466 1268 5468 1270
rect 5472 1268 5474 1270
rect 5496 1268 5498 1270
rect 5502 1268 5504 1270
rect 5526 1268 5528 1270
rect 5532 1268 5534 1270
rect 5676 1268 5678 1270
rect 5682 1268 5684 1270
rect 5706 1268 5708 1270
rect 5712 1268 5714 1270
rect 5736 1268 5738 1270
rect 5742 1268 5744 1270
rect 5766 1268 5768 1270
rect 5772 1268 5774 1270
rect 5796 1268 5798 1270
rect 5802 1268 5804 1270
rect 5826 1268 5828 1270
rect 5832 1268 5834 1270
rect 5856 1268 5858 1270
rect 5862 1268 5864 1270
rect 5886 1268 5888 1270
rect 5892 1268 5894 1270
rect 5916 1268 5918 1270
rect 5922 1268 5924 1270
rect 5946 1268 5948 1270
rect 5952 1268 5954 1270
rect 5976 1268 5978 1270
rect 5982 1268 5984 1270
rect 6006 1268 6008 1270
rect 6012 1268 6014 1270
rect 6036 1268 6038 1270
rect 6042 1268 6044 1270
rect 6066 1268 6068 1270
rect 6072 1268 6074 1270
rect 6096 1268 6098 1270
rect 6102 1268 6104 1270
rect 6126 1268 6128 1270
rect 6132 1268 6134 1270
rect 4484 1266 4486 1268
rect 4514 1266 4516 1268
rect 4544 1266 4546 1268
rect 4574 1266 4576 1268
rect 4604 1266 4606 1268
rect 4634 1266 4636 1268
rect 4664 1266 4666 1268
rect 4694 1266 4696 1268
rect 4724 1266 4726 1268
rect 4754 1266 4756 1268
rect 4784 1266 4786 1268
rect 4814 1266 4816 1268
rect 4844 1266 4846 1268
rect 4874 1266 4876 1268
rect 4904 1266 4906 1268
rect 4934 1266 4936 1268
rect 5084 1266 5086 1268
rect 5114 1266 5116 1268
rect 5144 1266 5146 1268
rect 5174 1266 5176 1268
rect 5204 1266 5206 1268
rect 5234 1266 5236 1268
rect 5264 1266 5266 1268
rect 5294 1266 5296 1268
rect 5324 1266 5326 1268
rect 5354 1266 5356 1268
rect 5384 1266 5386 1268
rect 5414 1266 5416 1268
rect 5444 1266 5446 1268
rect 5474 1266 5476 1268
rect 5504 1266 5506 1268
rect 5534 1266 5536 1268
rect 5684 1266 5686 1268
rect 5714 1266 5716 1268
rect 5744 1266 5746 1268
rect 5774 1266 5776 1268
rect 5804 1266 5806 1268
rect 5834 1266 5836 1268
rect 5864 1266 5866 1268
rect 5894 1266 5896 1268
rect 5924 1266 5926 1268
rect 5954 1266 5956 1268
rect 5984 1266 5986 1268
rect 6014 1266 6016 1268
rect 6044 1266 6046 1268
rect 6074 1266 6076 1268
rect 6104 1266 6106 1268
rect 6134 1266 6136 1268
rect 4484 1260 4486 1262
rect 4514 1260 4516 1262
rect 4544 1260 4546 1262
rect 4574 1260 4576 1262
rect 4604 1260 4606 1262
rect 4634 1260 4636 1262
rect 4664 1260 4666 1262
rect 4694 1260 4696 1262
rect 4724 1260 4726 1262
rect 4754 1260 4756 1262
rect 4784 1260 4786 1262
rect 4814 1260 4816 1262
rect 4844 1260 4846 1262
rect 4874 1260 4876 1262
rect 4904 1260 4906 1262
rect 4934 1260 4936 1262
rect 5084 1260 5086 1262
rect 5114 1260 5116 1262
rect 5144 1260 5146 1262
rect 5174 1260 5176 1262
rect 5204 1260 5206 1262
rect 5234 1260 5236 1262
rect 5264 1260 5266 1262
rect 5294 1260 5296 1262
rect 5324 1260 5326 1262
rect 5354 1260 5356 1262
rect 5384 1260 5386 1262
rect 5414 1260 5416 1262
rect 5444 1260 5446 1262
rect 5474 1260 5476 1262
rect 5504 1260 5506 1262
rect 5534 1260 5536 1262
rect 5684 1260 5686 1262
rect 5714 1260 5716 1262
rect 5744 1260 5746 1262
rect 5774 1260 5776 1262
rect 5804 1260 5806 1262
rect 5834 1260 5836 1262
rect 5864 1260 5866 1262
rect 5894 1260 5896 1262
rect 5924 1260 5926 1262
rect 5954 1260 5956 1262
rect 5984 1260 5986 1262
rect 6014 1260 6016 1262
rect 6044 1260 6046 1262
rect 6074 1260 6076 1262
rect 6104 1260 6106 1262
rect 6134 1260 6136 1262
rect 3250 1259 3252 1260
rect 3748 1259 3750 1260
rect 3850 1259 3852 1260
rect 4348 1259 4350 1260
rect 4476 1258 4478 1260
rect 4482 1258 4484 1260
rect 4506 1258 4508 1260
rect 4512 1258 4514 1260
rect 4536 1258 4538 1260
rect 4542 1258 4544 1260
rect 4566 1258 4568 1260
rect 4572 1258 4574 1260
rect 4596 1258 4598 1260
rect 4602 1258 4604 1260
rect 4626 1258 4628 1260
rect 4632 1258 4634 1260
rect 4656 1258 4658 1260
rect 4662 1258 4664 1260
rect 4686 1258 4688 1260
rect 4692 1258 4694 1260
rect 4716 1258 4718 1260
rect 4722 1258 4724 1260
rect 4746 1258 4748 1260
rect 4752 1258 4754 1260
rect 4776 1258 4778 1260
rect 4782 1258 4784 1260
rect 4806 1258 4808 1260
rect 4812 1258 4814 1260
rect 4836 1258 4838 1260
rect 4842 1258 4844 1260
rect 4866 1258 4868 1260
rect 4872 1258 4874 1260
rect 4896 1258 4898 1260
rect 4902 1258 4904 1260
rect 4926 1258 4928 1260
rect 4932 1258 4934 1260
rect 5076 1258 5078 1260
rect 5082 1258 5084 1260
rect 5106 1258 5108 1260
rect 5112 1258 5114 1260
rect 5136 1258 5138 1260
rect 5142 1258 5144 1260
rect 5166 1258 5168 1260
rect 5172 1258 5174 1260
rect 5196 1258 5198 1260
rect 5202 1258 5204 1260
rect 5226 1258 5228 1260
rect 5232 1258 5234 1260
rect 5256 1258 5258 1260
rect 5262 1258 5264 1260
rect 5286 1258 5288 1260
rect 5292 1258 5294 1260
rect 5316 1258 5318 1260
rect 5322 1258 5324 1260
rect 5346 1258 5348 1260
rect 5352 1258 5354 1260
rect 5376 1258 5378 1260
rect 5382 1258 5384 1260
rect 5406 1258 5408 1260
rect 5412 1258 5414 1260
rect 5436 1258 5438 1260
rect 5442 1258 5444 1260
rect 5466 1258 5468 1260
rect 5472 1258 5474 1260
rect 5496 1258 5498 1260
rect 5502 1258 5504 1260
rect 5526 1258 5528 1260
rect 5532 1258 5534 1260
rect 5676 1258 5678 1260
rect 5682 1258 5684 1260
rect 5706 1258 5708 1260
rect 5712 1258 5714 1260
rect 5736 1258 5738 1260
rect 5742 1258 5744 1260
rect 5766 1258 5768 1260
rect 5772 1258 5774 1260
rect 5796 1258 5798 1260
rect 5802 1258 5804 1260
rect 5826 1258 5828 1260
rect 5832 1258 5834 1260
rect 5856 1258 5858 1260
rect 5862 1258 5864 1260
rect 5886 1258 5888 1260
rect 5892 1258 5894 1260
rect 5916 1258 5918 1260
rect 5922 1258 5924 1260
rect 5946 1258 5948 1260
rect 5952 1258 5954 1260
rect 5976 1258 5978 1260
rect 5982 1258 5984 1260
rect 6006 1258 6008 1260
rect 6012 1258 6014 1260
rect 6036 1258 6038 1260
rect 6042 1258 6044 1260
rect 6066 1258 6068 1260
rect 6072 1258 6074 1260
rect 6096 1258 6098 1260
rect 6102 1258 6104 1260
rect 6126 1258 6128 1260
rect 6132 1258 6134 1260
rect 6250 1259 6252 1260
rect 6748 1259 6750 1260
rect 3248 1257 3250 1258
rect 3750 1257 3752 1258
rect 3848 1257 3850 1258
rect 4350 1257 4352 1258
rect 4474 1256 4476 1258
rect 4504 1256 4506 1258
rect 4534 1256 4536 1258
rect 4564 1256 4566 1258
rect 4594 1256 4596 1258
rect 4624 1256 4626 1258
rect 4654 1256 4656 1258
rect 4684 1256 4686 1258
rect 4714 1256 4716 1258
rect 4744 1256 4746 1258
rect 4774 1256 4776 1258
rect 4804 1256 4806 1258
rect 4834 1256 4836 1258
rect 4864 1256 4866 1258
rect 4894 1256 4896 1258
rect 4924 1256 4926 1258
rect 5074 1256 5076 1258
rect 5104 1256 5106 1258
rect 5134 1256 5136 1258
rect 5164 1256 5166 1258
rect 5194 1256 5196 1258
rect 5224 1256 5226 1258
rect 5254 1256 5256 1258
rect 5284 1256 5286 1258
rect 5314 1256 5316 1258
rect 5344 1256 5346 1258
rect 5374 1256 5376 1258
rect 5404 1256 5406 1258
rect 5434 1256 5436 1258
rect 5464 1256 5466 1258
rect 5494 1256 5496 1258
rect 5524 1256 5526 1258
rect 5674 1256 5676 1258
rect 5704 1256 5706 1258
rect 5734 1256 5736 1258
rect 5764 1256 5766 1258
rect 5794 1256 5796 1258
rect 5824 1256 5826 1258
rect 5854 1256 5856 1258
rect 5884 1256 5886 1258
rect 5914 1256 5916 1258
rect 5944 1256 5946 1258
rect 5974 1256 5976 1258
rect 6004 1256 6006 1258
rect 6034 1256 6036 1258
rect 6064 1256 6066 1258
rect 6094 1256 6096 1258
rect 6124 1256 6126 1258
rect 6248 1257 6250 1258
rect 6750 1257 6752 1258
rect 4474 1250 4476 1252
rect 4504 1250 4506 1252
rect 4534 1250 4536 1252
rect 4564 1250 4566 1252
rect 4594 1250 4596 1252
rect 4624 1250 4626 1252
rect 4654 1250 4656 1252
rect 4684 1250 4686 1252
rect 4714 1250 4716 1252
rect 4744 1250 4746 1252
rect 4774 1250 4776 1252
rect 4804 1250 4806 1252
rect 4834 1250 4836 1252
rect 4864 1250 4866 1252
rect 4894 1250 4896 1252
rect 4924 1250 4926 1252
rect 5074 1250 5076 1252
rect 5104 1250 5106 1252
rect 5134 1250 5136 1252
rect 5164 1250 5166 1252
rect 5194 1250 5196 1252
rect 5224 1250 5226 1252
rect 5254 1250 5256 1252
rect 5284 1250 5286 1252
rect 5314 1250 5316 1252
rect 5344 1250 5346 1252
rect 5374 1250 5376 1252
rect 5404 1250 5406 1252
rect 5434 1250 5436 1252
rect 5464 1250 5466 1252
rect 5494 1250 5496 1252
rect 5524 1250 5526 1252
rect 5674 1250 5676 1252
rect 5704 1250 5706 1252
rect 5734 1250 5736 1252
rect 5764 1250 5766 1252
rect 5794 1250 5796 1252
rect 5824 1250 5826 1252
rect 5854 1250 5856 1252
rect 5884 1250 5886 1252
rect 5914 1250 5916 1252
rect 5944 1250 5946 1252
rect 5974 1250 5976 1252
rect 6004 1250 6006 1252
rect 6034 1250 6036 1252
rect 6064 1250 6066 1252
rect 6094 1250 6096 1252
rect 6124 1250 6126 1252
rect 4476 1248 4478 1250
rect 4482 1248 4484 1250
rect 4506 1248 4508 1250
rect 4512 1248 4514 1250
rect 4536 1248 4538 1250
rect 4542 1248 4544 1250
rect 4566 1248 4568 1250
rect 4572 1248 4574 1250
rect 4596 1248 4598 1250
rect 4602 1248 4604 1250
rect 4626 1248 4628 1250
rect 4632 1248 4634 1250
rect 4656 1248 4658 1250
rect 4662 1248 4664 1250
rect 4686 1248 4688 1250
rect 4692 1248 4694 1250
rect 4716 1248 4718 1250
rect 4722 1248 4724 1250
rect 4746 1248 4748 1250
rect 4752 1248 4754 1250
rect 4776 1248 4778 1250
rect 4782 1248 4784 1250
rect 4806 1248 4808 1250
rect 4812 1248 4814 1250
rect 4836 1248 4838 1250
rect 4842 1248 4844 1250
rect 4866 1248 4868 1250
rect 4872 1248 4874 1250
rect 4896 1248 4898 1250
rect 4902 1248 4904 1250
rect 4926 1248 4928 1250
rect 4932 1248 4934 1250
rect 5076 1248 5078 1250
rect 5082 1248 5084 1250
rect 5106 1248 5108 1250
rect 5112 1248 5114 1250
rect 5136 1248 5138 1250
rect 5142 1248 5144 1250
rect 5166 1248 5168 1250
rect 5172 1248 5174 1250
rect 5196 1248 5198 1250
rect 5202 1248 5204 1250
rect 5226 1248 5228 1250
rect 5232 1248 5234 1250
rect 5256 1248 5258 1250
rect 5262 1248 5264 1250
rect 5286 1248 5288 1250
rect 5292 1248 5294 1250
rect 5316 1248 5318 1250
rect 5322 1248 5324 1250
rect 5346 1248 5348 1250
rect 5352 1248 5354 1250
rect 5376 1248 5378 1250
rect 5382 1248 5384 1250
rect 5406 1248 5408 1250
rect 5412 1248 5414 1250
rect 5436 1248 5438 1250
rect 5442 1248 5444 1250
rect 5466 1248 5468 1250
rect 5472 1248 5474 1250
rect 5496 1248 5498 1250
rect 5502 1248 5504 1250
rect 5526 1248 5528 1250
rect 5532 1248 5534 1250
rect 5676 1248 5678 1250
rect 5682 1248 5684 1250
rect 5706 1248 5708 1250
rect 5712 1248 5714 1250
rect 5736 1248 5738 1250
rect 5742 1248 5744 1250
rect 5766 1248 5768 1250
rect 5772 1248 5774 1250
rect 5796 1248 5798 1250
rect 5802 1248 5804 1250
rect 5826 1248 5828 1250
rect 5832 1248 5834 1250
rect 5856 1248 5858 1250
rect 5862 1248 5864 1250
rect 5886 1248 5888 1250
rect 5892 1248 5894 1250
rect 5916 1248 5918 1250
rect 5922 1248 5924 1250
rect 5946 1248 5948 1250
rect 5952 1248 5954 1250
rect 5976 1248 5978 1250
rect 5982 1248 5984 1250
rect 6006 1248 6008 1250
rect 6012 1248 6014 1250
rect 6036 1248 6038 1250
rect 6042 1248 6044 1250
rect 6066 1248 6068 1250
rect 6072 1248 6074 1250
rect 6096 1248 6098 1250
rect 6102 1248 6104 1250
rect 6126 1248 6128 1250
rect 6132 1248 6134 1250
rect 4484 1246 4486 1248
rect 4514 1246 4516 1248
rect 4544 1246 4546 1248
rect 4574 1246 4576 1248
rect 4604 1246 4606 1248
rect 4634 1246 4636 1248
rect 4664 1246 4666 1248
rect 4694 1246 4696 1248
rect 4724 1246 4726 1248
rect 4754 1246 4756 1248
rect 4784 1246 4786 1248
rect 4814 1246 4816 1248
rect 4844 1246 4846 1248
rect 4874 1246 4876 1248
rect 4904 1246 4906 1248
rect 4934 1246 4936 1248
rect 5084 1246 5086 1248
rect 5114 1246 5116 1248
rect 5144 1246 5146 1248
rect 5174 1246 5176 1248
rect 5204 1246 5206 1248
rect 5234 1246 5236 1248
rect 5264 1246 5266 1248
rect 5294 1246 5296 1248
rect 5324 1246 5326 1248
rect 5354 1246 5356 1248
rect 5384 1246 5386 1248
rect 5414 1246 5416 1248
rect 5444 1246 5446 1248
rect 5474 1246 5476 1248
rect 5504 1246 5506 1248
rect 5534 1246 5536 1248
rect 5684 1246 5686 1248
rect 5714 1246 5716 1248
rect 5744 1246 5746 1248
rect 5774 1246 5776 1248
rect 5804 1246 5806 1248
rect 5834 1246 5836 1248
rect 5864 1246 5866 1248
rect 5894 1246 5896 1248
rect 5924 1246 5926 1248
rect 5954 1246 5956 1248
rect 5984 1246 5986 1248
rect 6014 1246 6016 1248
rect 6044 1246 6046 1248
rect 6074 1246 6076 1248
rect 6104 1246 6106 1248
rect 6134 1246 6136 1248
rect 3296 1242 3298 1244
rect 3702 1242 3704 1244
rect 3896 1242 3898 1244
rect 4302 1242 4304 1244
rect 6296 1242 6298 1244
rect 6702 1242 6704 1244
rect 3294 1240 3296 1242
rect 3704 1240 3706 1242
rect 3894 1240 3896 1242
rect 4304 1240 4306 1242
rect 4484 1240 4486 1242
rect 4514 1240 4516 1242
rect 4544 1240 4546 1242
rect 4574 1240 4576 1242
rect 4604 1240 4606 1242
rect 4634 1240 4636 1242
rect 4664 1240 4666 1242
rect 4694 1240 4696 1242
rect 4724 1240 4726 1242
rect 4754 1240 4756 1242
rect 4784 1240 4786 1242
rect 4814 1240 4816 1242
rect 4844 1240 4846 1242
rect 4874 1240 4876 1242
rect 4904 1240 4906 1242
rect 4934 1240 4936 1242
rect 5084 1240 5086 1242
rect 5114 1240 5116 1242
rect 5144 1240 5146 1242
rect 5174 1240 5176 1242
rect 5204 1240 5206 1242
rect 5234 1240 5236 1242
rect 5264 1240 5266 1242
rect 5294 1240 5296 1242
rect 5324 1240 5326 1242
rect 5354 1240 5356 1242
rect 5384 1240 5386 1242
rect 5414 1240 5416 1242
rect 5444 1240 5446 1242
rect 5474 1240 5476 1242
rect 5504 1240 5506 1242
rect 5534 1240 5536 1242
rect 5684 1240 5686 1242
rect 5714 1240 5716 1242
rect 5744 1240 5746 1242
rect 5774 1240 5776 1242
rect 5804 1240 5806 1242
rect 5834 1240 5836 1242
rect 5864 1240 5866 1242
rect 5894 1240 5896 1242
rect 5924 1240 5926 1242
rect 5954 1240 5956 1242
rect 5984 1240 5986 1242
rect 6014 1240 6016 1242
rect 6044 1240 6046 1242
rect 6074 1240 6076 1242
rect 6104 1240 6106 1242
rect 6134 1240 6136 1242
rect 6294 1240 6296 1242
rect 6704 1240 6706 1242
rect 3250 1239 3252 1240
rect 3748 1239 3750 1240
rect 3850 1239 3852 1240
rect 4348 1239 4350 1240
rect 4476 1238 4478 1240
rect 4482 1238 4484 1240
rect 4506 1238 4508 1240
rect 4512 1238 4514 1240
rect 4536 1238 4538 1240
rect 4542 1238 4544 1240
rect 4566 1238 4568 1240
rect 4572 1238 4574 1240
rect 4596 1238 4598 1240
rect 4602 1238 4604 1240
rect 4626 1238 4628 1240
rect 4632 1238 4634 1240
rect 4656 1238 4658 1240
rect 4662 1238 4664 1240
rect 4686 1238 4688 1240
rect 4692 1238 4694 1240
rect 4716 1238 4718 1240
rect 4722 1238 4724 1240
rect 4746 1238 4748 1240
rect 4752 1238 4754 1240
rect 4776 1238 4778 1240
rect 4782 1238 4784 1240
rect 4806 1238 4808 1240
rect 4812 1238 4814 1240
rect 4836 1238 4838 1240
rect 4842 1238 4844 1240
rect 4866 1238 4868 1240
rect 4872 1238 4874 1240
rect 4896 1238 4898 1240
rect 4902 1238 4904 1240
rect 4926 1238 4928 1240
rect 4932 1238 4934 1240
rect 5076 1238 5078 1240
rect 5082 1238 5084 1240
rect 5106 1238 5108 1240
rect 5112 1238 5114 1240
rect 5136 1238 5138 1240
rect 5142 1238 5144 1240
rect 5166 1238 5168 1240
rect 5172 1238 5174 1240
rect 5196 1238 5198 1240
rect 5202 1238 5204 1240
rect 5226 1238 5228 1240
rect 5232 1238 5234 1240
rect 5256 1238 5258 1240
rect 5262 1238 5264 1240
rect 5286 1238 5288 1240
rect 5292 1238 5294 1240
rect 5316 1238 5318 1240
rect 5322 1238 5324 1240
rect 5346 1238 5348 1240
rect 5352 1238 5354 1240
rect 5376 1238 5378 1240
rect 5382 1238 5384 1240
rect 5406 1238 5408 1240
rect 5412 1238 5414 1240
rect 5436 1238 5438 1240
rect 5442 1238 5444 1240
rect 5466 1238 5468 1240
rect 5472 1238 5474 1240
rect 5496 1238 5498 1240
rect 5502 1238 5504 1240
rect 5526 1238 5528 1240
rect 5532 1238 5534 1240
rect 5676 1238 5678 1240
rect 5682 1238 5684 1240
rect 5706 1238 5708 1240
rect 5712 1238 5714 1240
rect 5736 1238 5738 1240
rect 5742 1238 5744 1240
rect 5766 1238 5768 1240
rect 5772 1238 5774 1240
rect 5796 1238 5798 1240
rect 5802 1238 5804 1240
rect 5826 1238 5828 1240
rect 5832 1238 5834 1240
rect 5856 1238 5858 1240
rect 5862 1238 5864 1240
rect 5886 1238 5888 1240
rect 5892 1238 5894 1240
rect 5916 1238 5918 1240
rect 5922 1238 5924 1240
rect 5946 1238 5948 1240
rect 5952 1238 5954 1240
rect 5976 1238 5978 1240
rect 5982 1238 5984 1240
rect 6006 1238 6008 1240
rect 6012 1238 6014 1240
rect 6036 1238 6038 1240
rect 6042 1238 6044 1240
rect 6066 1238 6068 1240
rect 6072 1238 6074 1240
rect 6096 1238 6098 1240
rect 6102 1238 6104 1240
rect 6126 1238 6128 1240
rect 6132 1238 6134 1240
rect 6250 1239 6252 1240
rect 6748 1239 6750 1240
rect 3248 1237 3250 1238
rect 3750 1237 3752 1238
rect 3848 1237 3850 1238
rect 4350 1237 4352 1238
rect 4474 1236 4476 1238
rect 4504 1236 4506 1238
rect 4534 1236 4536 1238
rect 4564 1236 4566 1238
rect 4594 1236 4596 1238
rect 4624 1236 4626 1238
rect 4654 1236 4656 1238
rect 4684 1236 4686 1238
rect 4714 1236 4716 1238
rect 4744 1236 4746 1238
rect 4774 1236 4776 1238
rect 4804 1236 4806 1238
rect 4834 1236 4836 1238
rect 4864 1236 4866 1238
rect 4894 1236 4896 1238
rect 4924 1236 4926 1238
rect 5074 1236 5076 1238
rect 5104 1236 5106 1238
rect 5134 1236 5136 1238
rect 5164 1236 5166 1238
rect 5194 1236 5196 1238
rect 5224 1236 5226 1238
rect 5254 1236 5256 1238
rect 5284 1236 5286 1238
rect 5314 1236 5316 1238
rect 5344 1236 5346 1238
rect 5374 1236 5376 1238
rect 5404 1236 5406 1238
rect 5434 1236 5436 1238
rect 5464 1236 5466 1238
rect 5494 1236 5496 1238
rect 5524 1236 5526 1238
rect 5674 1236 5676 1238
rect 5704 1236 5706 1238
rect 5734 1236 5736 1238
rect 5764 1236 5766 1238
rect 5794 1236 5796 1238
rect 5824 1236 5826 1238
rect 5854 1236 5856 1238
rect 5884 1236 5886 1238
rect 5914 1236 5916 1238
rect 5944 1236 5946 1238
rect 5974 1236 5976 1238
rect 6004 1236 6006 1238
rect 6034 1236 6036 1238
rect 6064 1236 6066 1238
rect 6094 1236 6096 1238
rect 6124 1236 6126 1238
rect 6248 1237 6250 1238
rect 6750 1237 6752 1238
rect 4474 1230 4476 1232
rect 4504 1230 4506 1232
rect 4534 1230 4536 1232
rect 4564 1230 4566 1232
rect 4594 1230 4596 1232
rect 4624 1230 4626 1232
rect 4654 1230 4656 1232
rect 4684 1230 4686 1232
rect 4714 1230 4716 1232
rect 4744 1230 4746 1232
rect 4774 1230 4776 1232
rect 4804 1230 4806 1232
rect 4834 1230 4836 1232
rect 4864 1230 4866 1232
rect 4894 1230 4896 1232
rect 4924 1230 4926 1232
rect 5074 1230 5076 1232
rect 5104 1230 5106 1232
rect 5134 1230 5136 1232
rect 5164 1230 5166 1232
rect 5194 1230 5196 1232
rect 5224 1230 5226 1232
rect 5254 1230 5256 1232
rect 5284 1230 5286 1232
rect 5314 1230 5316 1232
rect 5344 1230 5346 1232
rect 5374 1230 5376 1232
rect 5404 1230 5406 1232
rect 5434 1230 5436 1232
rect 5464 1230 5466 1232
rect 5494 1230 5496 1232
rect 5524 1230 5526 1232
rect 5674 1230 5676 1232
rect 5704 1230 5706 1232
rect 5734 1230 5736 1232
rect 5764 1230 5766 1232
rect 5794 1230 5796 1232
rect 5824 1230 5826 1232
rect 5854 1230 5856 1232
rect 5884 1230 5886 1232
rect 5914 1230 5916 1232
rect 5944 1230 5946 1232
rect 5974 1230 5976 1232
rect 6004 1230 6006 1232
rect 6034 1230 6036 1232
rect 6064 1230 6066 1232
rect 6094 1230 6096 1232
rect 6124 1230 6126 1232
rect 4476 1228 4478 1230
rect 4482 1228 4484 1230
rect 4506 1228 4508 1230
rect 4512 1228 4514 1230
rect 4536 1228 4538 1230
rect 4542 1228 4544 1230
rect 4566 1228 4568 1230
rect 4572 1228 4574 1230
rect 4596 1228 4598 1230
rect 4602 1228 4604 1230
rect 4626 1228 4628 1230
rect 4632 1228 4634 1230
rect 4656 1228 4658 1230
rect 4662 1228 4664 1230
rect 4686 1228 4688 1230
rect 4692 1228 4694 1230
rect 4716 1228 4718 1230
rect 4722 1228 4724 1230
rect 4746 1228 4748 1230
rect 4752 1228 4754 1230
rect 4776 1228 4778 1230
rect 4782 1228 4784 1230
rect 4806 1228 4808 1230
rect 4812 1228 4814 1230
rect 4836 1228 4838 1230
rect 4842 1228 4844 1230
rect 4866 1228 4868 1230
rect 4872 1228 4874 1230
rect 4896 1228 4898 1230
rect 4902 1228 4904 1230
rect 4926 1228 4928 1230
rect 4932 1228 4934 1230
rect 5076 1228 5078 1230
rect 5082 1228 5084 1230
rect 5106 1228 5108 1230
rect 5112 1228 5114 1230
rect 5136 1228 5138 1230
rect 5142 1228 5144 1230
rect 5166 1228 5168 1230
rect 5172 1228 5174 1230
rect 5196 1228 5198 1230
rect 5202 1228 5204 1230
rect 5226 1228 5228 1230
rect 5232 1228 5234 1230
rect 5256 1228 5258 1230
rect 5262 1228 5264 1230
rect 5286 1228 5288 1230
rect 5292 1228 5294 1230
rect 5316 1228 5318 1230
rect 5322 1228 5324 1230
rect 5346 1228 5348 1230
rect 5352 1228 5354 1230
rect 5376 1228 5378 1230
rect 5382 1228 5384 1230
rect 5406 1228 5408 1230
rect 5412 1228 5414 1230
rect 5436 1228 5438 1230
rect 5442 1228 5444 1230
rect 5466 1228 5468 1230
rect 5472 1228 5474 1230
rect 5496 1228 5498 1230
rect 5502 1228 5504 1230
rect 5526 1228 5528 1230
rect 5532 1228 5534 1230
rect 5676 1228 5678 1230
rect 5682 1228 5684 1230
rect 5706 1228 5708 1230
rect 5712 1228 5714 1230
rect 5736 1228 5738 1230
rect 5742 1228 5744 1230
rect 5766 1228 5768 1230
rect 5772 1228 5774 1230
rect 5796 1228 5798 1230
rect 5802 1228 5804 1230
rect 5826 1228 5828 1230
rect 5832 1228 5834 1230
rect 5856 1228 5858 1230
rect 5862 1228 5864 1230
rect 5886 1228 5888 1230
rect 5892 1228 5894 1230
rect 5916 1228 5918 1230
rect 5922 1228 5924 1230
rect 5946 1228 5948 1230
rect 5952 1228 5954 1230
rect 5976 1228 5978 1230
rect 5982 1228 5984 1230
rect 6006 1228 6008 1230
rect 6012 1228 6014 1230
rect 6036 1228 6038 1230
rect 6042 1228 6044 1230
rect 6066 1228 6068 1230
rect 6072 1228 6074 1230
rect 6096 1228 6098 1230
rect 6102 1228 6104 1230
rect 6126 1228 6128 1230
rect 6132 1228 6134 1230
rect 4484 1226 4486 1228
rect 4514 1226 4516 1228
rect 4544 1226 4546 1228
rect 4574 1226 4576 1228
rect 4604 1226 4606 1228
rect 4634 1226 4636 1228
rect 4664 1226 4666 1228
rect 4694 1226 4696 1228
rect 4724 1226 4726 1228
rect 4754 1226 4756 1228
rect 4784 1226 4786 1228
rect 4814 1226 4816 1228
rect 4844 1226 4846 1228
rect 4874 1226 4876 1228
rect 4904 1226 4906 1228
rect 4934 1226 4936 1228
rect 5084 1226 5086 1228
rect 5114 1226 5116 1228
rect 5144 1226 5146 1228
rect 5174 1226 5176 1228
rect 5204 1226 5206 1228
rect 5234 1226 5236 1228
rect 5264 1226 5266 1228
rect 5294 1226 5296 1228
rect 5324 1226 5326 1228
rect 5354 1226 5356 1228
rect 5384 1226 5386 1228
rect 5414 1226 5416 1228
rect 5444 1226 5446 1228
rect 5474 1226 5476 1228
rect 5504 1226 5506 1228
rect 5534 1226 5536 1228
rect 5684 1226 5686 1228
rect 5714 1226 5716 1228
rect 5744 1226 5746 1228
rect 5774 1226 5776 1228
rect 5804 1226 5806 1228
rect 5834 1226 5836 1228
rect 5864 1226 5866 1228
rect 5894 1226 5896 1228
rect 5924 1226 5926 1228
rect 5954 1226 5956 1228
rect 5984 1226 5986 1228
rect 6014 1226 6016 1228
rect 6044 1226 6046 1228
rect 6074 1226 6076 1228
rect 6104 1226 6106 1228
rect 6134 1226 6136 1228
rect 4484 1220 4486 1222
rect 4514 1220 4516 1222
rect 4544 1220 4546 1222
rect 4574 1220 4576 1222
rect 4604 1220 4606 1222
rect 4634 1220 4636 1222
rect 4664 1220 4666 1222
rect 4694 1220 4696 1222
rect 4724 1220 4726 1222
rect 4754 1220 4756 1222
rect 4784 1220 4786 1222
rect 4814 1220 4816 1222
rect 4844 1220 4846 1222
rect 4874 1220 4876 1222
rect 4904 1220 4906 1222
rect 4934 1220 4936 1222
rect 5084 1220 5086 1222
rect 5114 1220 5116 1222
rect 5144 1220 5146 1222
rect 5174 1220 5176 1222
rect 5204 1220 5206 1222
rect 5234 1220 5236 1222
rect 5264 1220 5266 1222
rect 5294 1220 5296 1222
rect 5324 1220 5326 1222
rect 5354 1220 5356 1222
rect 5384 1220 5386 1222
rect 5414 1220 5416 1222
rect 5444 1220 5446 1222
rect 5474 1220 5476 1222
rect 5504 1220 5506 1222
rect 5534 1220 5536 1222
rect 5684 1220 5686 1222
rect 5714 1220 5716 1222
rect 5744 1220 5746 1222
rect 5774 1220 5776 1222
rect 5804 1220 5806 1222
rect 5834 1220 5836 1222
rect 5864 1220 5866 1222
rect 5894 1220 5896 1222
rect 5924 1220 5926 1222
rect 5954 1220 5956 1222
rect 5984 1220 5986 1222
rect 6014 1220 6016 1222
rect 6044 1220 6046 1222
rect 6074 1220 6076 1222
rect 6104 1220 6106 1222
rect 6134 1220 6136 1222
rect 3250 1219 3252 1220
rect 3748 1219 3750 1220
rect 3850 1219 3852 1220
rect 4348 1219 4350 1220
rect 4476 1218 4478 1220
rect 4482 1218 4484 1220
rect 4506 1218 4508 1220
rect 4512 1218 4514 1220
rect 4536 1218 4538 1220
rect 4542 1218 4544 1220
rect 4566 1218 4568 1220
rect 4572 1218 4574 1220
rect 4596 1218 4598 1220
rect 4602 1218 4604 1220
rect 4626 1218 4628 1220
rect 4632 1218 4634 1220
rect 4656 1218 4658 1220
rect 4662 1218 4664 1220
rect 4686 1218 4688 1220
rect 4692 1218 4694 1220
rect 4716 1218 4718 1220
rect 4722 1218 4724 1220
rect 4746 1218 4748 1220
rect 4752 1218 4754 1220
rect 4776 1218 4778 1220
rect 4782 1218 4784 1220
rect 4806 1218 4808 1220
rect 4812 1218 4814 1220
rect 4836 1218 4838 1220
rect 4842 1218 4844 1220
rect 4866 1218 4868 1220
rect 4872 1218 4874 1220
rect 4896 1218 4898 1220
rect 4902 1218 4904 1220
rect 4926 1218 4928 1220
rect 4932 1218 4934 1220
rect 5076 1218 5078 1220
rect 5082 1218 5084 1220
rect 5106 1218 5108 1220
rect 5112 1218 5114 1220
rect 5136 1218 5138 1220
rect 5142 1218 5144 1220
rect 5166 1218 5168 1220
rect 5172 1218 5174 1220
rect 5196 1218 5198 1220
rect 5202 1218 5204 1220
rect 5226 1218 5228 1220
rect 5232 1218 5234 1220
rect 5256 1218 5258 1220
rect 5262 1218 5264 1220
rect 5286 1218 5288 1220
rect 5292 1218 5294 1220
rect 5316 1218 5318 1220
rect 5322 1218 5324 1220
rect 5346 1218 5348 1220
rect 5352 1218 5354 1220
rect 5376 1218 5378 1220
rect 5382 1218 5384 1220
rect 5406 1218 5408 1220
rect 5412 1218 5414 1220
rect 5436 1218 5438 1220
rect 5442 1218 5444 1220
rect 5466 1218 5468 1220
rect 5472 1218 5474 1220
rect 5496 1218 5498 1220
rect 5502 1218 5504 1220
rect 5526 1218 5528 1220
rect 5532 1218 5534 1220
rect 5676 1218 5678 1220
rect 5682 1218 5684 1220
rect 5706 1218 5708 1220
rect 5712 1218 5714 1220
rect 5736 1218 5738 1220
rect 5742 1218 5744 1220
rect 5766 1218 5768 1220
rect 5772 1218 5774 1220
rect 5796 1218 5798 1220
rect 5802 1218 5804 1220
rect 5826 1218 5828 1220
rect 5832 1218 5834 1220
rect 5856 1218 5858 1220
rect 5862 1218 5864 1220
rect 5886 1218 5888 1220
rect 5892 1218 5894 1220
rect 5916 1218 5918 1220
rect 5922 1218 5924 1220
rect 5946 1218 5948 1220
rect 5952 1218 5954 1220
rect 5976 1218 5978 1220
rect 5982 1218 5984 1220
rect 6006 1218 6008 1220
rect 6012 1218 6014 1220
rect 6036 1218 6038 1220
rect 6042 1218 6044 1220
rect 6066 1218 6068 1220
rect 6072 1218 6074 1220
rect 6096 1218 6098 1220
rect 6102 1218 6104 1220
rect 6126 1218 6128 1220
rect 6132 1218 6134 1220
rect 6250 1219 6252 1220
rect 6748 1219 6750 1220
rect 3248 1217 3250 1218
rect 3750 1217 3752 1218
rect 3848 1217 3850 1218
rect 4350 1217 4352 1218
rect 4474 1216 4476 1218
rect 4504 1216 4506 1218
rect 4534 1216 4536 1218
rect 4564 1216 4566 1218
rect 4594 1216 4596 1218
rect 4624 1216 4626 1218
rect 4654 1216 4656 1218
rect 4684 1216 4686 1218
rect 4714 1216 4716 1218
rect 4744 1216 4746 1218
rect 4774 1216 4776 1218
rect 4804 1216 4806 1218
rect 4834 1216 4836 1218
rect 4864 1216 4866 1218
rect 4894 1216 4896 1218
rect 4924 1216 4926 1218
rect 5074 1216 5076 1218
rect 5104 1216 5106 1218
rect 5134 1216 5136 1218
rect 5164 1216 5166 1218
rect 5194 1216 5196 1218
rect 5224 1216 5226 1218
rect 5254 1216 5256 1218
rect 5284 1216 5286 1218
rect 5314 1216 5316 1218
rect 5344 1216 5346 1218
rect 5374 1216 5376 1218
rect 5404 1216 5406 1218
rect 5434 1216 5436 1218
rect 5464 1216 5466 1218
rect 5494 1216 5496 1218
rect 5524 1216 5526 1218
rect 5674 1216 5676 1218
rect 5704 1216 5706 1218
rect 5734 1216 5736 1218
rect 5764 1216 5766 1218
rect 5794 1216 5796 1218
rect 5824 1216 5826 1218
rect 5854 1216 5856 1218
rect 5884 1216 5886 1218
rect 5914 1216 5916 1218
rect 5944 1216 5946 1218
rect 5974 1216 5976 1218
rect 6004 1216 6006 1218
rect 6034 1216 6036 1218
rect 6064 1216 6066 1218
rect 6094 1216 6096 1218
rect 6124 1216 6126 1218
rect 6248 1217 6250 1218
rect 6750 1217 6752 1218
rect 4474 1210 4476 1212
rect 4504 1210 4506 1212
rect 4534 1210 4536 1212
rect 4564 1210 4566 1212
rect 4594 1210 4596 1212
rect 4624 1210 4626 1212
rect 4654 1210 4656 1212
rect 4684 1210 4686 1212
rect 4714 1210 4716 1212
rect 4744 1210 4746 1212
rect 4774 1210 4776 1212
rect 4804 1210 4806 1212
rect 4834 1210 4836 1212
rect 4864 1210 4866 1212
rect 4894 1210 4896 1212
rect 4924 1210 4926 1212
rect 5074 1210 5076 1212
rect 5104 1210 5106 1212
rect 5134 1210 5136 1212
rect 5164 1210 5166 1212
rect 5194 1210 5196 1212
rect 5224 1210 5226 1212
rect 5254 1210 5256 1212
rect 5284 1210 5286 1212
rect 5314 1210 5316 1212
rect 5344 1210 5346 1212
rect 5374 1210 5376 1212
rect 5404 1210 5406 1212
rect 5434 1210 5436 1212
rect 5464 1210 5466 1212
rect 5494 1210 5496 1212
rect 5524 1210 5526 1212
rect 5674 1210 5676 1212
rect 5704 1210 5706 1212
rect 5734 1210 5736 1212
rect 5764 1210 5766 1212
rect 5794 1210 5796 1212
rect 5824 1210 5826 1212
rect 5854 1210 5856 1212
rect 5884 1210 5886 1212
rect 5914 1210 5916 1212
rect 5944 1210 5946 1212
rect 5974 1210 5976 1212
rect 6004 1210 6006 1212
rect 6034 1210 6036 1212
rect 6064 1210 6066 1212
rect 6094 1210 6096 1212
rect 6124 1210 6126 1212
rect 4476 1208 4478 1210
rect 4482 1208 4484 1210
rect 4506 1208 4508 1210
rect 4512 1208 4514 1210
rect 4536 1208 4538 1210
rect 4542 1208 4544 1210
rect 4566 1208 4568 1210
rect 4572 1208 4574 1210
rect 4596 1208 4598 1210
rect 4602 1208 4604 1210
rect 4626 1208 4628 1210
rect 4632 1208 4634 1210
rect 4656 1208 4658 1210
rect 4662 1208 4664 1210
rect 4686 1208 4688 1210
rect 4692 1208 4694 1210
rect 4716 1208 4718 1210
rect 4722 1208 4724 1210
rect 4746 1208 4748 1210
rect 4752 1208 4754 1210
rect 4776 1208 4778 1210
rect 4782 1208 4784 1210
rect 4806 1208 4808 1210
rect 4812 1208 4814 1210
rect 4836 1208 4838 1210
rect 4842 1208 4844 1210
rect 4866 1208 4868 1210
rect 4872 1208 4874 1210
rect 4896 1208 4898 1210
rect 4902 1208 4904 1210
rect 4926 1208 4928 1210
rect 4932 1208 4934 1210
rect 5076 1208 5078 1210
rect 5082 1208 5084 1210
rect 5106 1208 5108 1210
rect 5112 1208 5114 1210
rect 5136 1208 5138 1210
rect 5142 1208 5144 1210
rect 5166 1208 5168 1210
rect 5172 1208 5174 1210
rect 5196 1208 5198 1210
rect 5202 1208 5204 1210
rect 5226 1208 5228 1210
rect 5232 1208 5234 1210
rect 5256 1208 5258 1210
rect 5262 1208 5264 1210
rect 5286 1208 5288 1210
rect 5292 1208 5294 1210
rect 5316 1208 5318 1210
rect 5322 1208 5324 1210
rect 5346 1208 5348 1210
rect 5352 1208 5354 1210
rect 5376 1208 5378 1210
rect 5382 1208 5384 1210
rect 5406 1208 5408 1210
rect 5412 1208 5414 1210
rect 5436 1208 5438 1210
rect 5442 1208 5444 1210
rect 5466 1208 5468 1210
rect 5472 1208 5474 1210
rect 5496 1208 5498 1210
rect 5502 1208 5504 1210
rect 5526 1208 5528 1210
rect 5532 1208 5534 1210
rect 5676 1208 5678 1210
rect 5682 1208 5684 1210
rect 5706 1208 5708 1210
rect 5712 1208 5714 1210
rect 5736 1208 5738 1210
rect 5742 1208 5744 1210
rect 5766 1208 5768 1210
rect 5772 1208 5774 1210
rect 5796 1208 5798 1210
rect 5802 1208 5804 1210
rect 5826 1208 5828 1210
rect 5832 1208 5834 1210
rect 5856 1208 5858 1210
rect 5862 1208 5864 1210
rect 5886 1208 5888 1210
rect 5892 1208 5894 1210
rect 5916 1208 5918 1210
rect 5922 1208 5924 1210
rect 5946 1208 5948 1210
rect 5952 1208 5954 1210
rect 5976 1208 5978 1210
rect 5982 1208 5984 1210
rect 6006 1208 6008 1210
rect 6012 1208 6014 1210
rect 6036 1208 6038 1210
rect 6042 1208 6044 1210
rect 6066 1208 6068 1210
rect 6072 1208 6074 1210
rect 6096 1208 6098 1210
rect 6102 1208 6104 1210
rect 6126 1208 6128 1210
rect 6132 1208 6134 1210
rect 4484 1206 4486 1208
rect 4514 1206 4516 1208
rect 4544 1206 4546 1208
rect 4574 1206 4576 1208
rect 4604 1206 4606 1208
rect 4634 1206 4636 1208
rect 4664 1206 4666 1208
rect 4694 1206 4696 1208
rect 4724 1206 4726 1208
rect 4754 1206 4756 1208
rect 4784 1206 4786 1208
rect 4814 1206 4816 1208
rect 4844 1206 4846 1208
rect 4874 1206 4876 1208
rect 4904 1206 4906 1208
rect 4934 1206 4936 1208
rect 5084 1206 5086 1208
rect 5114 1206 5116 1208
rect 5144 1206 5146 1208
rect 5174 1206 5176 1208
rect 5204 1206 5206 1208
rect 5234 1206 5236 1208
rect 5264 1206 5266 1208
rect 5294 1206 5296 1208
rect 5324 1206 5326 1208
rect 5354 1206 5356 1208
rect 5384 1206 5386 1208
rect 5414 1206 5416 1208
rect 5444 1206 5446 1208
rect 5474 1206 5476 1208
rect 5504 1206 5506 1208
rect 5534 1206 5536 1208
rect 5684 1206 5686 1208
rect 5714 1206 5716 1208
rect 5744 1206 5746 1208
rect 5774 1206 5776 1208
rect 5804 1206 5806 1208
rect 5834 1206 5836 1208
rect 5864 1206 5866 1208
rect 5894 1206 5896 1208
rect 5924 1206 5926 1208
rect 5954 1206 5956 1208
rect 5984 1206 5986 1208
rect 6014 1206 6016 1208
rect 6044 1206 6046 1208
rect 6074 1206 6076 1208
rect 6104 1206 6106 1208
rect 6134 1206 6136 1208
rect 4484 1200 4486 1202
rect 4514 1200 4516 1202
rect 4544 1200 4546 1202
rect 4574 1200 4576 1202
rect 4604 1200 4606 1202
rect 4634 1200 4636 1202
rect 4664 1200 4666 1202
rect 4694 1200 4696 1202
rect 4724 1200 4726 1202
rect 4754 1200 4756 1202
rect 4784 1200 4786 1202
rect 4814 1200 4816 1202
rect 4844 1200 4846 1202
rect 4874 1200 4876 1202
rect 4904 1200 4906 1202
rect 4934 1200 4936 1202
rect 5084 1200 5086 1202
rect 5114 1200 5116 1202
rect 5144 1200 5146 1202
rect 5174 1200 5176 1202
rect 5204 1200 5206 1202
rect 5234 1200 5236 1202
rect 5264 1200 5266 1202
rect 5294 1200 5296 1202
rect 5324 1200 5326 1202
rect 5354 1200 5356 1202
rect 5384 1200 5386 1202
rect 5414 1200 5416 1202
rect 5444 1200 5446 1202
rect 5474 1200 5476 1202
rect 5504 1200 5506 1202
rect 5534 1200 5536 1202
rect 5684 1200 5686 1202
rect 5714 1200 5716 1202
rect 5744 1200 5746 1202
rect 5774 1200 5776 1202
rect 5804 1200 5806 1202
rect 5834 1200 5836 1202
rect 5864 1200 5866 1202
rect 5894 1200 5896 1202
rect 5924 1200 5926 1202
rect 5954 1200 5956 1202
rect 5984 1200 5986 1202
rect 6014 1200 6016 1202
rect 6044 1200 6046 1202
rect 6074 1200 6076 1202
rect 6104 1200 6106 1202
rect 6134 1200 6136 1202
rect 3250 1199 3252 1200
rect 3748 1199 3750 1200
rect 3850 1199 3852 1200
rect 4348 1199 4350 1200
rect 4476 1198 4478 1200
rect 4482 1198 4484 1200
rect 4506 1198 4508 1200
rect 4512 1198 4514 1200
rect 4536 1198 4538 1200
rect 4542 1198 4544 1200
rect 4566 1198 4568 1200
rect 4572 1198 4574 1200
rect 4596 1198 4598 1200
rect 4602 1198 4604 1200
rect 4626 1198 4628 1200
rect 4632 1198 4634 1200
rect 4656 1198 4658 1200
rect 4662 1198 4664 1200
rect 4686 1198 4688 1200
rect 4692 1198 4694 1200
rect 4716 1198 4718 1200
rect 4722 1198 4724 1200
rect 4746 1198 4748 1200
rect 4752 1198 4754 1200
rect 4776 1198 4778 1200
rect 4782 1198 4784 1200
rect 4806 1198 4808 1200
rect 4812 1198 4814 1200
rect 4836 1198 4838 1200
rect 4842 1198 4844 1200
rect 4866 1198 4868 1200
rect 4872 1198 4874 1200
rect 4896 1198 4898 1200
rect 4902 1198 4904 1200
rect 4926 1198 4928 1200
rect 4932 1198 4934 1200
rect 5076 1198 5078 1200
rect 5082 1198 5084 1200
rect 5106 1198 5108 1200
rect 5112 1198 5114 1200
rect 5136 1198 5138 1200
rect 5142 1198 5144 1200
rect 5166 1198 5168 1200
rect 5172 1198 5174 1200
rect 5196 1198 5198 1200
rect 5202 1198 5204 1200
rect 5226 1198 5228 1200
rect 5232 1198 5234 1200
rect 5256 1198 5258 1200
rect 5262 1198 5264 1200
rect 5286 1198 5288 1200
rect 5292 1198 5294 1200
rect 5316 1198 5318 1200
rect 5322 1198 5324 1200
rect 5346 1198 5348 1200
rect 5352 1198 5354 1200
rect 5376 1198 5378 1200
rect 5382 1198 5384 1200
rect 5406 1198 5408 1200
rect 5412 1198 5414 1200
rect 5436 1198 5438 1200
rect 5442 1198 5444 1200
rect 5466 1198 5468 1200
rect 5472 1198 5474 1200
rect 5496 1198 5498 1200
rect 5502 1198 5504 1200
rect 5526 1198 5528 1200
rect 5532 1198 5534 1200
rect 5676 1198 5678 1200
rect 5682 1198 5684 1200
rect 5706 1198 5708 1200
rect 5712 1198 5714 1200
rect 5736 1198 5738 1200
rect 5742 1198 5744 1200
rect 5766 1198 5768 1200
rect 5772 1198 5774 1200
rect 5796 1198 5798 1200
rect 5802 1198 5804 1200
rect 5826 1198 5828 1200
rect 5832 1198 5834 1200
rect 5856 1198 5858 1200
rect 5862 1198 5864 1200
rect 5886 1198 5888 1200
rect 5892 1198 5894 1200
rect 5916 1198 5918 1200
rect 5922 1198 5924 1200
rect 5946 1198 5948 1200
rect 5952 1198 5954 1200
rect 5976 1198 5978 1200
rect 5982 1198 5984 1200
rect 6006 1198 6008 1200
rect 6012 1198 6014 1200
rect 6036 1198 6038 1200
rect 6042 1198 6044 1200
rect 6066 1198 6068 1200
rect 6072 1198 6074 1200
rect 6096 1198 6098 1200
rect 6102 1198 6104 1200
rect 6126 1198 6128 1200
rect 6132 1198 6134 1200
rect 6250 1199 6252 1200
rect 6748 1199 6750 1200
rect 3248 1197 3250 1198
rect 3750 1197 3752 1198
rect 3848 1197 3850 1198
rect 4350 1197 4352 1198
rect 4474 1196 4476 1198
rect 4504 1196 4506 1198
rect 4534 1196 4536 1198
rect 4564 1196 4566 1198
rect 4594 1196 4596 1198
rect 4624 1196 4626 1198
rect 4654 1196 4656 1198
rect 4684 1196 4686 1198
rect 4714 1196 4716 1198
rect 4744 1196 4746 1198
rect 4774 1196 4776 1198
rect 4804 1196 4806 1198
rect 4834 1196 4836 1198
rect 4864 1196 4866 1198
rect 4894 1196 4896 1198
rect 4924 1196 4926 1198
rect 5074 1196 5076 1198
rect 5104 1196 5106 1198
rect 5134 1196 5136 1198
rect 5164 1196 5166 1198
rect 5194 1196 5196 1198
rect 5224 1196 5226 1198
rect 5254 1196 5256 1198
rect 5284 1196 5286 1198
rect 5314 1196 5316 1198
rect 5344 1196 5346 1198
rect 5374 1196 5376 1198
rect 5404 1196 5406 1198
rect 5434 1196 5436 1198
rect 5464 1196 5466 1198
rect 5494 1196 5496 1198
rect 5524 1196 5526 1198
rect 5674 1196 5676 1198
rect 5704 1196 5706 1198
rect 5734 1196 5736 1198
rect 5764 1196 5766 1198
rect 5794 1196 5796 1198
rect 5824 1196 5826 1198
rect 5854 1196 5856 1198
rect 5884 1196 5886 1198
rect 5914 1196 5916 1198
rect 5944 1196 5946 1198
rect 5974 1196 5976 1198
rect 6004 1196 6006 1198
rect 6034 1196 6036 1198
rect 6064 1196 6066 1198
rect 6094 1196 6096 1198
rect 6124 1196 6126 1198
rect 6248 1197 6250 1198
rect 6750 1197 6752 1198
rect 4474 1190 4476 1192
rect 4924 1190 4926 1192
rect 5074 1190 5076 1192
rect 5524 1190 5526 1192
rect 5674 1190 5676 1192
rect 6124 1190 6126 1192
rect 4476 1188 4478 1190
rect 4482 1188 4484 1190
rect 4926 1188 4928 1190
rect 4932 1188 4934 1190
rect 5076 1188 5078 1190
rect 5082 1188 5084 1190
rect 5526 1188 5528 1190
rect 5532 1188 5534 1190
rect 5676 1188 5678 1190
rect 5682 1188 5684 1190
rect 6126 1188 6128 1190
rect 6132 1188 6134 1190
rect 4484 1186 4486 1188
rect 4934 1186 4936 1188
rect 5084 1186 5086 1188
rect 5534 1186 5536 1188
rect 5684 1186 5686 1188
rect 6134 1186 6136 1188
rect 3294 1180 3296 1182
rect 3704 1180 3706 1182
rect 3894 1180 3896 1182
rect 4304 1180 4306 1182
rect 4484 1180 4486 1182
rect 4934 1180 4936 1182
rect 5084 1180 5086 1182
rect 5534 1180 5536 1182
rect 5684 1180 5686 1182
rect 6134 1180 6136 1182
rect 6294 1180 6296 1182
rect 6704 1180 6706 1182
rect 3250 1179 3252 1180
rect 3296 1178 3298 1180
rect 3702 1178 3704 1180
rect 3748 1179 3750 1180
rect 3850 1179 3852 1180
rect 3896 1178 3898 1180
rect 4302 1178 4304 1180
rect 4348 1179 4350 1180
rect 4476 1178 4478 1180
rect 4482 1178 4484 1180
rect 4926 1178 4928 1180
rect 4932 1178 4934 1180
rect 5076 1178 5078 1180
rect 5082 1178 5084 1180
rect 5526 1178 5528 1180
rect 5532 1178 5534 1180
rect 5676 1178 5678 1180
rect 5682 1178 5684 1180
rect 6126 1178 6128 1180
rect 6132 1178 6134 1180
rect 6250 1179 6252 1180
rect 6296 1178 6298 1180
rect 6702 1178 6704 1180
rect 6748 1179 6750 1180
rect 3248 1177 3250 1178
rect 3750 1177 3752 1178
rect 3848 1177 3850 1178
rect 4350 1177 4352 1178
rect 4474 1176 4476 1178
rect 4924 1176 4926 1178
rect 5074 1176 5076 1178
rect 5524 1176 5526 1178
rect 5674 1176 5676 1178
rect 6124 1176 6126 1178
rect 6248 1177 6250 1178
rect 6750 1177 6752 1178
rect 4474 1170 4476 1172
rect 4504 1170 4506 1172
rect 4534 1170 4536 1172
rect 4564 1170 4566 1172
rect 4594 1170 4596 1172
rect 4624 1170 4626 1172
rect 4654 1170 4656 1172
rect 4684 1170 4686 1172
rect 4714 1170 4716 1172
rect 4744 1170 4746 1172
rect 4774 1170 4776 1172
rect 4804 1170 4806 1172
rect 4834 1170 4836 1172
rect 4864 1170 4866 1172
rect 4894 1170 4896 1172
rect 4924 1170 4926 1172
rect 5074 1170 5076 1172
rect 5104 1170 5106 1172
rect 5134 1170 5136 1172
rect 5164 1170 5166 1172
rect 5194 1170 5196 1172
rect 5224 1170 5226 1172
rect 5254 1170 5256 1172
rect 5284 1170 5286 1172
rect 5314 1170 5316 1172
rect 5344 1170 5346 1172
rect 5374 1170 5376 1172
rect 5404 1170 5406 1172
rect 5434 1170 5436 1172
rect 5464 1170 5466 1172
rect 5494 1170 5496 1172
rect 5524 1170 5526 1172
rect 5674 1170 5676 1172
rect 5704 1170 5706 1172
rect 5734 1170 5736 1172
rect 5764 1170 5766 1172
rect 5794 1170 5796 1172
rect 5824 1170 5826 1172
rect 5854 1170 5856 1172
rect 5884 1170 5886 1172
rect 5914 1170 5916 1172
rect 5944 1170 5946 1172
rect 5974 1170 5976 1172
rect 6004 1170 6006 1172
rect 6034 1170 6036 1172
rect 6064 1170 6066 1172
rect 6094 1170 6096 1172
rect 6124 1170 6126 1172
rect 4476 1168 4478 1170
rect 4482 1168 4484 1170
rect 4506 1168 4508 1170
rect 4512 1168 4514 1170
rect 4536 1168 4538 1170
rect 4542 1168 4544 1170
rect 4566 1168 4568 1170
rect 4572 1168 4574 1170
rect 4596 1168 4598 1170
rect 4602 1168 4604 1170
rect 4626 1168 4628 1170
rect 4632 1168 4634 1170
rect 4656 1168 4658 1170
rect 4662 1168 4664 1170
rect 4686 1168 4688 1170
rect 4692 1168 4694 1170
rect 4716 1168 4718 1170
rect 4722 1168 4724 1170
rect 4746 1168 4748 1170
rect 4752 1168 4754 1170
rect 4776 1168 4778 1170
rect 4782 1168 4784 1170
rect 4806 1168 4808 1170
rect 4812 1168 4814 1170
rect 4836 1168 4838 1170
rect 4842 1168 4844 1170
rect 4866 1168 4868 1170
rect 4872 1168 4874 1170
rect 4896 1168 4898 1170
rect 4902 1168 4904 1170
rect 4926 1168 4928 1170
rect 4932 1168 4934 1170
rect 5076 1168 5078 1170
rect 5082 1168 5084 1170
rect 5106 1168 5108 1170
rect 5112 1168 5114 1170
rect 5136 1168 5138 1170
rect 5142 1168 5144 1170
rect 5166 1168 5168 1170
rect 5172 1168 5174 1170
rect 5196 1168 5198 1170
rect 5202 1168 5204 1170
rect 5226 1168 5228 1170
rect 5232 1168 5234 1170
rect 5256 1168 5258 1170
rect 5262 1168 5264 1170
rect 5286 1168 5288 1170
rect 5292 1168 5294 1170
rect 5316 1168 5318 1170
rect 5322 1168 5324 1170
rect 5346 1168 5348 1170
rect 5352 1168 5354 1170
rect 5376 1168 5378 1170
rect 5382 1168 5384 1170
rect 5406 1168 5408 1170
rect 5412 1168 5414 1170
rect 5436 1168 5438 1170
rect 5442 1168 5444 1170
rect 5466 1168 5468 1170
rect 5472 1168 5474 1170
rect 5496 1168 5498 1170
rect 5502 1168 5504 1170
rect 5526 1168 5528 1170
rect 5532 1168 5534 1170
rect 5676 1168 5678 1170
rect 5682 1168 5684 1170
rect 5706 1168 5708 1170
rect 5712 1168 5714 1170
rect 5736 1168 5738 1170
rect 5742 1168 5744 1170
rect 5766 1168 5768 1170
rect 5772 1168 5774 1170
rect 5796 1168 5798 1170
rect 5802 1168 5804 1170
rect 5826 1168 5828 1170
rect 5832 1168 5834 1170
rect 5856 1168 5858 1170
rect 5862 1168 5864 1170
rect 5886 1168 5888 1170
rect 5892 1168 5894 1170
rect 5916 1168 5918 1170
rect 5922 1168 5924 1170
rect 5946 1168 5948 1170
rect 5952 1168 5954 1170
rect 5976 1168 5978 1170
rect 5982 1168 5984 1170
rect 6006 1168 6008 1170
rect 6012 1168 6014 1170
rect 6036 1168 6038 1170
rect 6042 1168 6044 1170
rect 6066 1168 6068 1170
rect 6072 1168 6074 1170
rect 6096 1168 6098 1170
rect 6102 1168 6104 1170
rect 6126 1168 6128 1170
rect 6132 1168 6134 1170
rect 4484 1166 4486 1168
rect 4514 1166 4516 1168
rect 4544 1166 4546 1168
rect 4574 1166 4576 1168
rect 4604 1166 4606 1168
rect 4634 1166 4636 1168
rect 4664 1166 4666 1168
rect 4694 1166 4696 1168
rect 4724 1166 4726 1168
rect 4754 1166 4756 1168
rect 4784 1166 4786 1168
rect 4814 1166 4816 1168
rect 4844 1166 4846 1168
rect 4874 1166 4876 1168
rect 4904 1166 4906 1168
rect 4934 1166 4936 1168
rect 5084 1166 5086 1168
rect 5114 1166 5116 1168
rect 5144 1166 5146 1168
rect 5174 1166 5176 1168
rect 5204 1166 5206 1168
rect 5234 1166 5236 1168
rect 5264 1166 5266 1168
rect 5294 1166 5296 1168
rect 5324 1166 5326 1168
rect 5354 1166 5356 1168
rect 5384 1166 5386 1168
rect 5414 1166 5416 1168
rect 5444 1166 5446 1168
rect 5474 1166 5476 1168
rect 5504 1166 5506 1168
rect 5534 1166 5536 1168
rect 5684 1166 5686 1168
rect 5714 1166 5716 1168
rect 5744 1166 5746 1168
rect 5774 1166 5776 1168
rect 5804 1166 5806 1168
rect 5834 1166 5836 1168
rect 5864 1166 5866 1168
rect 5894 1166 5896 1168
rect 5924 1166 5926 1168
rect 5954 1166 5956 1168
rect 5984 1166 5986 1168
rect 6014 1166 6016 1168
rect 6044 1166 6046 1168
rect 6074 1166 6076 1168
rect 6104 1166 6106 1168
rect 6134 1166 6136 1168
rect 4484 1160 4486 1162
rect 4514 1160 4516 1162
rect 4544 1160 4546 1162
rect 4574 1160 4576 1162
rect 4604 1160 4606 1162
rect 4634 1160 4636 1162
rect 4664 1160 4666 1162
rect 4694 1160 4696 1162
rect 4724 1160 4726 1162
rect 4754 1160 4756 1162
rect 4784 1160 4786 1162
rect 4814 1160 4816 1162
rect 4844 1160 4846 1162
rect 4874 1160 4876 1162
rect 4904 1160 4906 1162
rect 4934 1160 4936 1162
rect 5084 1160 5086 1162
rect 5114 1160 5116 1162
rect 5144 1160 5146 1162
rect 5174 1160 5176 1162
rect 5204 1160 5206 1162
rect 5234 1160 5236 1162
rect 5264 1160 5266 1162
rect 5294 1160 5296 1162
rect 5324 1160 5326 1162
rect 5354 1160 5356 1162
rect 5384 1160 5386 1162
rect 5414 1160 5416 1162
rect 5444 1160 5446 1162
rect 5474 1160 5476 1162
rect 5504 1160 5506 1162
rect 5534 1160 5536 1162
rect 5684 1160 5686 1162
rect 5714 1160 5716 1162
rect 5744 1160 5746 1162
rect 5774 1160 5776 1162
rect 5804 1160 5806 1162
rect 5834 1160 5836 1162
rect 5864 1160 5866 1162
rect 5894 1160 5896 1162
rect 5924 1160 5926 1162
rect 5954 1160 5956 1162
rect 5984 1160 5986 1162
rect 6014 1160 6016 1162
rect 6044 1160 6046 1162
rect 6074 1160 6076 1162
rect 6104 1160 6106 1162
rect 6134 1160 6136 1162
rect 3250 1159 3252 1160
rect 3748 1159 3750 1160
rect 3850 1159 3852 1160
rect 4348 1159 4350 1160
rect 4476 1158 4478 1160
rect 4482 1158 4484 1160
rect 4506 1158 4508 1160
rect 4512 1158 4514 1160
rect 4536 1158 4538 1160
rect 4542 1158 4544 1160
rect 4566 1158 4568 1160
rect 4572 1158 4574 1160
rect 4596 1158 4598 1160
rect 4602 1158 4604 1160
rect 4626 1158 4628 1160
rect 4632 1158 4634 1160
rect 4656 1158 4658 1160
rect 4662 1158 4664 1160
rect 4686 1158 4688 1160
rect 4692 1158 4694 1160
rect 4716 1158 4718 1160
rect 4722 1158 4724 1160
rect 4746 1158 4748 1160
rect 4752 1158 4754 1160
rect 4776 1158 4778 1160
rect 4782 1158 4784 1160
rect 4806 1158 4808 1160
rect 4812 1158 4814 1160
rect 4836 1158 4838 1160
rect 4842 1158 4844 1160
rect 4866 1158 4868 1160
rect 4872 1158 4874 1160
rect 4896 1158 4898 1160
rect 4902 1158 4904 1160
rect 4926 1158 4928 1160
rect 4932 1158 4934 1160
rect 5076 1158 5078 1160
rect 5082 1158 5084 1160
rect 5106 1158 5108 1160
rect 5112 1158 5114 1160
rect 5136 1158 5138 1160
rect 5142 1158 5144 1160
rect 5166 1158 5168 1160
rect 5172 1158 5174 1160
rect 5196 1158 5198 1160
rect 5202 1158 5204 1160
rect 5226 1158 5228 1160
rect 5232 1158 5234 1160
rect 5256 1158 5258 1160
rect 5262 1158 5264 1160
rect 5286 1158 5288 1160
rect 5292 1158 5294 1160
rect 5316 1158 5318 1160
rect 5322 1158 5324 1160
rect 5346 1158 5348 1160
rect 5352 1158 5354 1160
rect 5376 1158 5378 1160
rect 5382 1158 5384 1160
rect 5406 1158 5408 1160
rect 5412 1158 5414 1160
rect 5436 1158 5438 1160
rect 5442 1158 5444 1160
rect 5466 1158 5468 1160
rect 5472 1158 5474 1160
rect 5496 1158 5498 1160
rect 5502 1158 5504 1160
rect 5526 1158 5528 1160
rect 5532 1158 5534 1160
rect 5676 1158 5678 1160
rect 5682 1158 5684 1160
rect 5706 1158 5708 1160
rect 5712 1158 5714 1160
rect 5736 1158 5738 1160
rect 5742 1158 5744 1160
rect 5766 1158 5768 1160
rect 5772 1158 5774 1160
rect 5796 1158 5798 1160
rect 5802 1158 5804 1160
rect 5826 1158 5828 1160
rect 5832 1158 5834 1160
rect 5856 1158 5858 1160
rect 5862 1158 5864 1160
rect 5886 1158 5888 1160
rect 5892 1158 5894 1160
rect 5916 1158 5918 1160
rect 5922 1158 5924 1160
rect 5946 1158 5948 1160
rect 5952 1158 5954 1160
rect 5976 1158 5978 1160
rect 5982 1158 5984 1160
rect 6006 1158 6008 1160
rect 6012 1158 6014 1160
rect 6036 1158 6038 1160
rect 6042 1158 6044 1160
rect 6066 1158 6068 1160
rect 6072 1158 6074 1160
rect 6096 1158 6098 1160
rect 6102 1158 6104 1160
rect 6126 1158 6128 1160
rect 6132 1158 6134 1160
rect 6250 1159 6252 1160
rect 6748 1159 6750 1160
rect 3248 1157 3250 1158
rect 3750 1157 3752 1158
rect 3848 1157 3850 1158
rect 4350 1157 4352 1158
rect 4474 1156 4476 1158
rect 4504 1156 4506 1158
rect 4534 1156 4536 1158
rect 4564 1156 4566 1158
rect 4594 1156 4596 1158
rect 4624 1156 4626 1158
rect 4654 1156 4656 1158
rect 4684 1156 4686 1158
rect 4714 1156 4716 1158
rect 4744 1156 4746 1158
rect 4774 1156 4776 1158
rect 4804 1156 4806 1158
rect 4834 1156 4836 1158
rect 4864 1156 4866 1158
rect 4894 1156 4896 1158
rect 4924 1156 4926 1158
rect 5074 1156 5076 1158
rect 5104 1156 5106 1158
rect 5134 1156 5136 1158
rect 5164 1156 5166 1158
rect 5194 1156 5196 1158
rect 5224 1156 5226 1158
rect 5254 1156 5256 1158
rect 5284 1156 5286 1158
rect 5314 1156 5316 1158
rect 5344 1156 5346 1158
rect 5374 1156 5376 1158
rect 5404 1156 5406 1158
rect 5434 1156 5436 1158
rect 5464 1156 5466 1158
rect 5494 1156 5496 1158
rect 5524 1156 5526 1158
rect 5674 1156 5676 1158
rect 5704 1156 5706 1158
rect 5734 1156 5736 1158
rect 5764 1156 5766 1158
rect 5794 1156 5796 1158
rect 5824 1156 5826 1158
rect 5854 1156 5856 1158
rect 5884 1156 5886 1158
rect 5914 1156 5916 1158
rect 5944 1156 5946 1158
rect 5974 1156 5976 1158
rect 6004 1156 6006 1158
rect 6034 1156 6036 1158
rect 6064 1156 6066 1158
rect 6094 1156 6096 1158
rect 6124 1156 6126 1158
rect 6248 1157 6250 1158
rect 6750 1157 6752 1158
rect 4474 1150 4476 1152
rect 4504 1150 4506 1152
rect 4534 1150 4536 1152
rect 4564 1150 4566 1152
rect 4594 1150 4596 1152
rect 4624 1150 4626 1152
rect 4654 1150 4656 1152
rect 4684 1150 4686 1152
rect 4714 1150 4716 1152
rect 4744 1150 4746 1152
rect 4774 1150 4776 1152
rect 4804 1150 4806 1152
rect 4834 1150 4836 1152
rect 4864 1150 4866 1152
rect 4894 1150 4896 1152
rect 4924 1150 4926 1152
rect 5074 1150 5076 1152
rect 5104 1150 5106 1152
rect 5134 1150 5136 1152
rect 5164 1150 5166 1152
rect 5194 1150 5196 1152
rect 5224 1150 5226 1152
rect 5254 1150 5256 1152
rect 5284 1150 5286 1152
rect 5314 1150 5316 1152
rect 5344 1150 5346 1152
rect 5374 1150 5376 1152
rect 5404 1150 5406 1152
rect 5434 1150 5436 1152
rect 5464 1150 5466 1152
rect 5494 1150 5496 1152
rect 5524 1150 5526 1152
rect 5674 1150 5676 1152
rect 5704 1150 5706 1152
rect 5734 1150 5736 1152
rect 5764 1150 5766 1152
rect 5794 1150 5796 1152
rect 5824 1150 5826 1152
rect 5854 1150 5856 1152
rect 5884 1150 5886 1152
rect 5914 1150 5916 1152
rect 5944 1150 5946 1152
rect 5974 1150 5976 1152
rect 6004 1150 6006 1152
rect 6034 1150 6036 1152
rect 6064 1150 6066 1152
rect 6094 1150 6096 1152
rect 6124 1150 6126 1152
rect 4476 1148 4478 1150
rect 4482 1148 4484 1150
rect 4506 1148 4508 1150
rect 4512 1148 4514 1150
rect 4536 1148 4538 1150
rect 4542 1148 4544 1150
rect 4566 1148 4568 1150
rect 4572 1148 4574 1150
rect 4596 1148 4598 1150
rect 4602 1148 4604 1150
rect 4626 1148 4628 1150
rect 4632 1148 4634 1150
rect 4656 1148 4658 1150
rect 4662 1148 4664 1150
rect 4686 1148 4688 1150
rect 4692 1148 4694 1150
rect 4716 1148 4718 1150
rect 4722 1148 4724 1150
rect 4746 1148 4748 1150
rect 4752 1148 4754 1150
rect 4776 1148 4778 1150
rect 4782 1148 4784 1150
rect 4806 1148 4808 1150
rect 4812 1148 4814 1150
rect 4836 1148 4838 1150
rect 4842 1148 4844 1150
rect 4866 1148 4868 1150
rect 4872 1148 4874 1150
rect 4896 1148 4898 1150
rect 4902 1148 4904 1150
rect 4926 1148 4928 1150
rect 4932 1148 4934 1150
rect 5076 1148 5078 1150
rect 5082 1148 5084 1150
rect 5106 1148 5108 1150
rect 5112 1148 5114 1150
rect 5136 1148 5138 1150
rect 5142 1148 5144 1150
rect 5166 1148 5168 1150
rect 5172 1148 5174 1150
rect 5196 1148 5198 1150
rect 5202 1148 5204 1150
rect 5226 1148 5228 1150
rect 5232 1148 5234 1150
rect 5256 1148 5258 1150
rect 5262 1148 5264 1150
rect 5286 1148 5288 1150
rect 5292 1148 5294 1150
rect 5316 1148 5318 1150
rect 5322 1148 5324 1150
rect 5346 1148 5348 1150
rect 5352 1148 5354 1150
rect 5376 1148 5378 1150
rect 5382 1148 5384 1150
rect 5406 1148 5408 1150
rect 5412 1148 5414 1150
rect 5436 1148 5438 1150
rect 5442 1148 5444 1150
rect 5466 1148 5468 1150
rect 5472 1148 5474 1150
rect 5496 1148 5498 1150
rect 5502 1148 5504 1150
rect 5526 1148 5528 1150
rect 5532 1148 5534 1150
rect 5676 1148 5678 1150
rect 5682 1148 5684 1150
rect 5706 1148 5708 1150
rect 5712 1148 5714 1150
rect 5736 1148 5738 1150
rect 5742 1148 5744 1150
rect 5766 1148 5768 1150
rect 5772 1148 5774 1150
rect 5796 1148 5798 1150
rect 5802 1148 5804 1150
rect 5826 1148 5828 1150
rect 5832 1148 5834 1150
rect 5856 1148 5858 1150
rect 5862 1148 5864 1150
rect 5886 1148 5888 1150
rect 5892 1148 5894 1150
rect 5916 1148 5918 1150
rect 5922 1148 5924 1150
rect 5946 1148 5948 1150
rect 5952 1148 5954 1150
rect 5976 1148 5978 1150
rect 5982 1148 5984 1150
rect 6006 1148 6008 1150
rect 6012 1148 6014 1150
rect 6036 1148 6038 1150
rect 6042 1148 6044 1150
rect 6066 1148 6068 1150
rect 6072 1148 6074 1150
rect 6096 1148 6098 1150
rect 6102 1148 6104 1150
rect 6126 1148 6128 1150
rect 6132 1148 6134 1150
rect 4484 1146 4486 1148
rect 4514 1146 4516 1148
rect 4544 1146 4546 1148
rect 4574 1146 4576 1148
rect 4604 1146 4606 1148
rect 4634 1146 4636 1148
rect 4664 1146 4666 1148
rect 4694 1146 4696 1148
rect 4724 1146 4726 1148
rect 4754 1146 4756 1148
rect 4784 1146 4786 1148
rect 4814 1146 4816 1148
rect 4844 1146 4846 1148
rect 4874 1146 4876 1148
rect 4904 1146 4906 1148
rect 4934 1146 4936 1148
rect 5084 1146 5086 1148
rect 5114 1146 5116 1148
rect 5144 1146 5146 1148
rect 5174 1146 5176 1148
rect 5204 1146 5206 1148
rect 5234 1146 5236 1148
rect 5264 1146 5266 1148
rect 5294 1146 5296 1148
rect 5324 1146 5326 1148
rect 5354 1146 5356 1148
rect 5384 1146 5386 1148
rect 5414 1146 5416 1148
rect 5444 1146 5446 1148
rect 5474 1146 5476 1148
rect 5504 1146 5506 1148
rect 5534 1146 5536 1148
rect 5684 1146 5686 1148
rect 5714 1146 5716 1148
rect 5744 1146 5746 1148
rect 5774 1146 5776 1148
rect 5804 1146 5806 1148
rect 5834 1146 5836 1148
rect 5864 1146 5866 1148
rect 5894 1146 5896 1148
rect 5924 1146 5926 1148
rect 5954 1146 5956 1148
rect 5984 1146 5986 1148
rect 6014 1146 6016 1148
rect 6044 1146 6046 1148
rect 6074 1146 6076 1148
rect 6104 1146 6106 1148
rect 6134 1146 6136 1148
rect 4484 1140 4486 1142
rect 4514 1140 4516 1142
rect 4544 1140 4546 1142
rect 4574 1140 4576 1142
rect 4604 1140 4606 1142
rect 4634 1140 4636 1142
rect 4664 1140 4666 1142
rect 4694 1140 4696 1142
rect 4724 1140 4726 1142
rect 4754 1140 4756 1142
rect 4784 1140 4786 1142
rect 4814 1140 4816 1142
rect 4844 1140 4846 1142
rect 4874 1140 4876 1142
rect 4904 1140 4906 1142
rect 4934 1140 4936 1142
rect 5084 1140 5086 1142
rect 5114 1140 5116 1142
rect 5144 1140 5146 1142
rect 5174 1140 5176 1142
rect 5204 1140 5206 1142
rect 5234 1140 5236 1142
rect 5264 1140 5266 1142
rect 5294 1140 5296 1142
rect 5324 1140 5326 1142
rect 5354 1140 5356 1142
rect 5384 1140 5386 1142
rect 5414 1140 5416 1142
rect 5444 1140 5446 1142
rect 5474 1140 5476 1142
rect 5504 1140 5506 1142
rect 5534 1140 5536 1142
rect 5684 1140 5686 1142
rect 5714 1140 5716 1142
rect 5744 1140 5746 1142
rect 5774 1140 5776 1142
rect 5804 1140 5806 1142
rect 5834 1140 5836 1142
rect 5864 1140 5866 1142
rect 5894 1140 5896 1142
rect 5924 1140 5926 1142
rect 5954 1140 5956 1142
rect 5984 1140 5986 1142
rect 6014 1140 6016 1142
rect 6044 1140 6046 1142
rect 6074 1140 6076 1142
rect 6104 1140 6106 1142
rect 6134 1140 6136 1142
rect 3250 1139 3252 1140
rect 3748 1139 3750 1140
rect 3850 1139 3852 1140
rect 4348 1139 4350 1140
rect 4476 1138 4478 1140
rect 4482 1138 4484 1140
rect 4506 1138 4508 1140
rect 4512 1138 4514 1140
rect 4536 1138 4538 1140
rect 4542 1138 4544 1140
rect 4566 1138 4568 1140
rect 4572 1138 4574 1140
rect 4596 1138 4598 1140
rect 4602 1138 4604 1140
rect 4626 1138 4628 1140
rect 4632 1138 4634 1140
rect 4656 1138 4658 1140
rect 4662 1138 4664 1140
rect 4686 1138 4688 1140
rect 4692 1138 4694 1140
rect 4716 1138 4718 1140
rect 4722 1138 4724 1140
rect 4746 1138 4748 1140
rect 4752 1138 4754 1140
rect 4776 1138 4778 1140
rect 4782 1138 4784 1140
rect 4806 1138 4808 1140
rect 4812 1138 4814 1140
rect 4836 1138 4838 1140
rect 4842 1138 4844 1140
rect 4866 1138 4868 1140
rect 4872 1138 4874 1140
rect 4896 1138 4898 1140
rect 4902 1138 4904 1140
rect 4926 1138 4928 1140
rect 4932 1138 4934 1140
rect 5076 1138 5078 1140
rect 5082 1138 5084 1140
rect 5106 1138 5108 1140
rect 5112 1138 5114 1140
rect 5136 1138 5138 1140
rect 5142 1138 5144 1140
rect 5166 1138 5168 1140
rect 5172 1138 5174 1140
rect 5196 1138 5198 1140
rect 5202 1138 5204 1140
rect 5226 1138 5228 1140
rect 5232 1138 5234 1140
rect 5256 1138 5258 1140
rect 5262 1138 5264 1140
rect 5286 1138 5288 1140
rect 5292 1138 5294 1140
rect 5316 1138 5318 1140
rect 5322 1138 5324 1140
rect 5346 1138 5348 1140
rect 5352 1138 5354 1140
rect 5376 1138 5378 1140
rect 5382 1138 5384 1140
rect 5406 1138 5408 1140
rect 5412 1138 5414 1140
rect 5436 1138 5438 1140
rect 5442 1138 5444 1140
rect 5466 1138 5468 1140
rect 5472 1138 5474 1140
rect 5496 1138 5498 1140
rect 5502 1138 5504 1140
rect 5526 1138 5528 1140
rect 5532 1138 5534 1140
rect 5676 1138 5678 1140
rect 5682 1138 5684 1140
rect 5706 1138 5708 1140
rect 5712 1138 5714 1140
rect 5736 1138 5738 1140
rect 5742 1138 5744 1140
rect 5766 1138 5768 1140
rect 5772 1138 5774 1140
rect 5796 1138 5798 1140
rect 5802 1138 5804 1140
rect 5826 1138 5828 1140
rect 5832 1138 5834 1140
rect 5856 1138 5858 1140
rect 5862 1138 5864 1140
rect 5886 1138 5888 1140
rect 5892 1138 5894 1140
rect 5916 1138 5918 1140
rect 5922 1138 5924 1140
rect 5946 1138 5948 1140
rect 5952 1138 5954 1140
rect 5976 1138 5978 1140
rect 5982 1138 5984 1140
rect 6006 1138 6008 1140
rect 6012 1138 6014 1140
rect 6036 1138 6038 1140
rect 6042 1138 6044 1140
rect 6066 1138 6068 1140
rect 6072 1138 6074 1140
rect 6096 1138 6098 1140
rect 6102 1138 6104 1140
rect 6126 1138 6128 1140
rect 6132 1138 6134 1140
rect 6250 1139 6252 1140
rect 6748 1139 6750 1140
rect 3248 1137 3250 1138
rect 3750 1137 3752 1138
rect 3848 1137 3850 1138
rect 4350 1137 4352 1138
rect 4474 1136 4476 1138
rect 4504 1136 4506 1138
rect 4534 1136 4536 1138
rect 4564 1136 4566 1138
rect 4594 1136 4596 1138
rect 4624 1136 4626 1138
rect 4654 1136 4656 1138
rect 4684 1136 4686 1138
rect 4714 1136 4716 1138
rect 4744 1136 4746 1138
rect 4774 1136 4776 1138
rect 4804 1136 4806 1138
rect 4834 1136 4836 1138
rect 4864 1136 4866 1138
rect 4894 1136 4896 1138
rect 4924 1136 4926 1138
rect 5074 1136 5076 1138
rect 5104 1136 5106 1138
rect 5134 1136 5136 1138
rect 5164 1136 5166 1138
rect 5194 1136 5196 1138
rect 5224 1136 5226 1138
rect 5254 1136 5256 1138
rect 5284 1136 5286 1138
rect 5314 1136 5316 1138
rect 5344 1136 5346 1138
rect 5374 1136 5376 1138
rect 5404 1136 5406 1138
rect 5434 1136 5436 1138
rect 5464 1136 5466 1138
rect 5494 1136 5496 1138
rect 5524 1136 5526 1138
rect 5674 1136 5676 1138
rect 5704 1136 5706 1138
rect 5734 1136 5736 1138
rect 5764 1136 5766 1138
rect 5794 1136 5796 1138
rect 5824 1136 5826 1138
rect 5854 1136 5856 1138
rect 5884 1136 5886 1138
rect 5914 1136 5916 1138
rect 5944 1136 5946 1138
rect 5974 1136 5976 1138
rect 6004 1136 6006 1138
rect 6034 1136 6036 1138
rect 6064 1136 6066 1138
rect 6094 1136 6096 1138
rect 6124 1136 6126 1138
rect 6248 1137 6250 1138
rect 6750 1137 6752 1138
rect 4474 1130 4476 1132
rect 4504 1130 4506 1132
rect 4534 1130 4536 1132
rect 4564 1130 4566 1132
rect 4594 1130 4596 1132
rect 4624 1130 4626 1132
rect 4654 1130 4656 1132
rect 4684 1130 4686 1132
rect 4714 1130 4716 1132
rect 4744 1130 4746 1132
rect 4774 1130 4776 1132
rect 4804 1130 4806 1132
rect 4834 1130 4836 1132
rect 4864 1130 4866 1132
rect 4894 1130 4896 1132
rect 4924 1130 4926 1132
rect 5074 1130 5076 1132
rect 5104 1130 5106 1132
rect 5134 1130 5136 1132
rect 5164 1130 5166 1132
rect 5194 1130 5196 1132
rect 5224 1130 5226 1132
rect 5254 1130 5256 1132
rect 5284 1130 5286 1132
rect 5314 1130 5316 1132
rect 5344 1130 5346 1132
rect 5374 1130 5376 1132
rect 5404 1130 5406 1132
rect 5434 1130 5436 1132
rect 5464 1130 5466 1132
rect 5494 1130 5496 1132
rect 5524 1130 5526 1132
rect 5674 1130 5676 1132
rect 5704 1130 5706 1132
rect 5734 1130 5736 1132
rect 5764 1130 5766 1132
rect 5794 1130 5796 1132
rect 5824 1130 5826 1132
rect 5854 1130 5856 1132
rect 5884 1130 5886 1132
rect 5914 1130 5916 1132
rect 5944 1130 5946 1132
rect 5974 1130 5976 1132
rect 6004 1130 6006 1132
rect 6034 1130 6036 1132
rect 6064 1130 6066 1132
rect 6094 1130 6096 1132
rect 6124 1130 6126 1132
rect 4476 1128 4478 1130
rect 4482 1128 4484 1130
rect 4506 1128 4508 1130
rect 4512 1128 4514 1130
rect 4536 1128 4538 1130
rect 4542 1128 4544 1130
rect 4566 1128 4568 1130
rect 4572 1128 4574 1130
rect 4596 1128 4598 1130
rect 4602 1128 4604 1130
rect 4626 1128 4628 1130
rect 4632 1128 4634 1130
rect 4656 1128 4658 1130
rect 4662 1128 4664 1130
rect 4686 1128 4688 1130
rect 4692 1128 4694 1130
rect 4716 1128 4718 1130
rect 4722 1128 4724 1130
rect 4746 1128 4748 1130
rect 4752 1128 4754 1130
rect 4776 1128 4778 1130
rect 4782 1128 4784 1130
rect 4806 1128 4808 1130
rect 4812 1128 4814 1130
rect 4836 1128 4838 1130
rect 4842 1128 4844 1130
rect 4866 1128 4868 1130
rect 4872 1128 4874 1130
rect 4896 1128 4898 1130
rect 4902 1128 4904 1130
rect 4926 1128 4928 1130
rect 4932 1128 4934 1130
rect 5076 1128 5078 1130
rect 5082 1128 5084 1130
rect 5106 1128 5108 1130
rect 5112 1128 5114 1130
rect 5136 1128 5138 1130
rect 5142 1128 5144 1130
rect 5166 1128 5168 1130
rect 5172 1128 5174 1130
rect 5196 1128 5198 1130
rect 5202 1128 5204 1130
rect 5226 1128 5228 1130
rect 5232 1128 5234 1130
rect 5256 1128 5258 1130
rect 5262 1128 5264 1130
rect 5286 1128 5288 1130
rect 5292 1128 5294 1130
rect 5316 1128 5318 1130
rect 5322 1128 5324 1130
rect 5346 1128 5348 1130
rect 5352 1128 5354 1130
rect 5376 1128 5378 1130
rect 5382 1128 5384 1130
rect 5406 1128 5408 1130
rect 5412 1128 5414 1130
rect 5436 1128 5438 1130
rect 5442 1128 5444 1130
rect 5466 1128 5468 1130
rect 5472 1128 5474 1130
rect 5496 1128 5498 1130
rect 5502 1128 5504 1130
rect 5526 1128 5528 1130
rect 5532 1128 5534 1130
rect 5676 1128 5678 1130
rect 5682 1128 5684 1130
rect 5706 1128 5708 1130
rect 5712 1128 5714 1130
rect 5736 1128 5738 1130
rect 5742 1128 5744 1130
rect 5766 1128 5768 1130
rect 5772 1128 5774 1130
rect 5796 1128 5798 1130
rect 5802 1128 5804 1130
rect 5826 1128 5828 1130
rect 5832 1128 5834 1130
rect 5856 1128 5858 1130
rect 5862 1128 5864 1130
rect 5886 1128 5888 1130
rect 5892 1128 5894 1130
rect 5916 1128 5918 1130
rect 5922 1128 5924 1130
rect 5946 1128 5948 1130
rect 5952 1128 5954 1130
rect 5976 1128 5978 1130
rect 5982 1128 5984 1130
rect 6006 1128 6008 1130
rect 6012 1128 6014 1130
rect 6036 1128 6038 1130
rect 6042 1128 6044 1130
rect 6066 1128 6068 1130
rect 6072 1128 6074 1130
rect 6096 1128 6098 1130
rect 6102 1128 6104 1130
rect 6126 1128 6128 1130
rect 6132 1128 6134 1130
rect 4484 1126 4486 1128
rect 4514 1126 4516 1128
rect 4544 1126 4546 1128
rect 4574 1126 4576 1128
rect 4604 1126 4606 1128
rect 4634 1126 4636 1128
rect 4664 1126 4666 1128
rect 4694 1126 4696 1128
rect 4724 1126 4726 1128
rect 4754 1126 4756 1128
rect 4784 1126 4786 1128
rect 4814 1126 4816 1128
rect 4844 1126 4846 1128
rect 4874 1126 4876 1128
rect 4904 1126 4906 1128
rect 4934 1126 4936 1128
rect 5084 1126 5086 1128
rect 5114 1126 5116 1128
rect 5144 1126 5146 1128
rect 5174 1126 5176 1128
rect 5204 1126 5206 1128
rect 5234 1126 5236 1128
rect 5264 1126 5266 1128
rect 5294 1126 5296 1128
rect 5324 1126 5326 1128
rect 5354 1126 5356 1128
rect 5384 1126 5386 1128
rect 5414 1126 5416 1128
rect 5444 1126 5446 1128
rect 5474 1126 5476 1128
rect 5504 1126 5506 1128
rect 5534 1126 5536 1128
rect 5684 1126 5686 1128
rect 5714 1126 5716 1128
rect 5744 1126 5746 1128
rect 5774 1126 5776 1128
rect 5804 1126 5806 1128
rect 5834 1126 5836 1128
rect 5864 1126 5866 1128
rect 5894 1126 5896 1128
rect 5924 1126 5926 1128
rect 5954 1126 5956 1128
rect 5984 1126 5986 1128
rect 6014 1126 6016 1128
rect 6044 1126 6046 1128
rect 6074 1126 6076 1128
rect 6104 1126 6106 1128
rect 6134 1126 6136 1128
rect 4484 1120 4486 1122
rect 4904 1120 4906 1122
rect 4934 1120 4936 1122
rect 5084 1120 5086 1122
rect 5504 1120 5506 1122
rect 5534 1120 5536 1122
rect 5684 1120 5686 1122
rect 6104 1120 6106 1122
rect 6134 1120 6136 1122
rect 3250 1119 3252 1120
rect 3748 1119 3750 1120
rect 3850 1119 3852 1120
rect 4348 1119 4350 1120
rect 4486 1118 4488 1120
rect 4906 1118 4908 1120
rect 4932 1118 4934 1120
rect 5086 1118 5088 1120
rect 5506 1118 5508 1120
rect 5532 1118 5534 1120
rect 5686 1118 5688 1120
rect 6106 1118 6108 1120
rect 6132 1118 6134 1120
rect 6250 1119 6252 1120
rect 6748 1119 6750 1120
rect 3248 1117 3250 1118
rect 3750 1117 3752 1118
rect 3848 1117 3850 1118
rect 4350 1117 4352 1118
rect 6248 1117 6250 1118
rect 6750 1117 6752 1118
rect 3296 1114 3298 1116
rect 3702 1114 3704 1116
rect 3896 1114 3898 1116
rect 4302 1114 4304 1116
rect 6296 1114 6298 1116
rect 6702 1114 6704 1116
rect 3294 1112 3296 1114
rect 3704 1112 3706 1114
rect 3894 1112 3896 1114
rect 4304 1112 4306 1114
rect 6294 1112 6296 1114
rect 6704 1112 6706 1114
rect 4486 1108 4488 1110
rect 4906 1108 4908 1110
rect 4932 1108 4934 1110
rect 5086 1108 5088 1110
rect 5506 1108 5508 1110
rect 5532 1108 5534 1110
rect 5686 1108 5688 1110
rect 6106 1108 6108 1110
rect 6132 1108 6134 1110
rect 2102 1105 2104 1107
rect 2702 1105 2704 1107
rect 4484 1106 4486 1108
rect 4904 1106 4906 1108
rect 4934 1106 4936 1108
rect 5084 1106 5086 1108
rect 5504 1106 5506 1108
rect 5534 1106 5536 1108
rect 5684 1106 5686 1108
rect 6104 1106 6106 1108
rect 6134 1106 6136 1108
rect 6902 1105 6904 1107
rect 2100 1103 2102 1105
rect 2700 1103 2702 1105
rect 6900 1103 6902 1105
rect 4484 1100 4486 1102
rect 4514 1100 4516 1102
rect 4544 1100 4546 1102
rect 4574 1100 4576 1102
rect 4604 1100 4606 1102
rect 4634 1100 4636 1102
rect 4664 1100 4666 1102
rect 4694 1100 4696 1102
rect 4724 1100 4726 1102
rect 4754 1100 4756 1102
rect 4784 1100 4786 1102
rect 4814 1100 4816 1102
rect 4844 1100 4846 1102
rect 4874 1100 4876 1102
rect 4904 1100 4906 1102
rect 4934 1100 4936 1102
rect 5084 1100 5086 1102
rect 5114 1100 5116 1102
rect 5144 1100 5146 1102
rect 5174 1100 5176 1102
rect 5204 1100 5206 1102
rect 5234 1100 5236 1102
rect 5264 1100 5266 1102
rect 5294 1100 5296 1102
rect 5324 1100 5326 1102
rect 5354 1100 5356 1102
rect 5384 1100 5386 1102
rect 5414 1100 5416 1102
rect 5444 1100 5446 1102
rect 5474 1100 5476 1102
rect 5504 1100 5506 1102
rect 5534 1100 5536 1102
rect 5684 1100 5686 1102
rect 5714 1100 5716 1102
rect 5744 1100 5746 1102
rect 5774 1100 5776 1102
rect 5804 1100 5806 1102
rect 5834 1100 5836 1102
rect 5864 1100 5866 1102
rect 5894 1100 5896 1102
rect 5924 1100 5926 1102
rect 5954 1100 5956 1102
rect 5984 1100 5986 1102
rect 6014 1100 6016 1102
rect 6044 1100 6046 1102
rect 6074 1100 6076 1102
rect 6104 1100 6106 1102
rect 6134 1100 6136 1102
rect 3250 1099 3252 1100
rect 3748 1099 3750 1100
rect 3850 1099 3852 1100
rect 4348 1099 4350 1100
rect 4476 1098 4478 1100
rect 4482 1098 4484 1100
rect 4506 1098 4508 1100
rect 4512 1098 4514 1100
rect 4536 1098 4538 1100
rect 4542 1098 4544 1100
rect 4566 1098 4568 1100
rect 4572 1098 4574 1100
rect 4596 1098 4598 1100
rect 4602 1098 4604 1100
rect 4626 1098 4628 1100
rect 4632 1098 4634 1100
rect 4656 1098 4658 1100
rect 4662 1098 4664 1100
rect 4686 1098 4688 1100
rect 4692 1098 4694 1100
rect 4716 1098 4718 1100
rect 4722 1098 4724 1100
rect 4746 1098 4748 1100
rect 4752 1098 4754 1100
rect 4776 1098 4778 1100
rect 4782 1098 4784 1100
rect 4806 1098 4808 1100
rect 4812 1098 4814 1100
rect 4836 1098 4838 1100
rect 4842 1098 4844 1100
rect 4866 1098 4868 1100
rect 4872 1098 4874 1100
rect 4896 1098 4898 1100
rect 4902 1098 4904 1100
rect 4926 1098 4928 1100
rect 4932 1098 4934 1100
rect 5076 1098 5078 1100
rect 5082 1098 5084 1100
rect 5106 1098 5108 1100
rect 5112 1098 5114 1100
rect 5136 1098 5138 1100
rect 5142 1098 5144 1100
rect 5166 1098 5168 1100
rect 5172 1098 5174 1100
rect 5196 1098 5198 1100
rect 5202 1098 5204 1100
rect 5226 1098 5228 1100
rect 5232 1098 5234 1100
rect 5256 1098 5258 1100
rect 5262 1098 5264 1100
rect 5286 1098 5288 1100
rect 5292 1098 5294 1100
rect 5316 1098 5318 1100
rect 5322 1098 5324 1100
rect 5346 1098 5348 1100
rect 5352 1098 5354 1100
rect 5376 1098 5378 1100
rect 5382 1098 5384 1100
rect 5406 1098 5408 1100
rect 5412 1098 5414 1100
rect 5436 1098 5438 1100
rect 5442 1098 5444 1100
rect 5466 1098 5468 1100
rect 5472 1098 5474 1100
rect 5496 1098 5498 1100
rect 5502 1098 5504 1100
rect 5526 1098 5528 1100
rect 5532 1098 5534 1100
rect 5676 1098 5678 1100
rect 5682 1098 5684 1100
rect 5706 1098 5708 1100
rect 5712 1098 5714 1100
rect 5736 1098 5738 1100
rect 5742 1098 5744 1100
rect 5766 1098 5768 1100
rect 5772 1098 5774 1100
rect 5796 1098 5798 1100
rect 5802 1098 5804 1100
rect 5826 1098 5828 1100
rect 5832 1098 5834 1100
rect 5856 1098 5858 1100
rect 5862 1098 5864 1100
rect 5886 1098 5888 1100
rect 5892 1098 5894 1100
rect 5916 1098 5918 1100
rect 5922 1098 5924 1100
rect 5946 1098 5948 1100
rect 5952 1098 5954 1100
rect 5976 1098 5978 1100
rect 5982 1098 5984 1100
rect 6006 1098 6008 1100
rect 6012 1098 6014 1100
rect 6036 1098 6038 1100
rect 6042 1098 6044 1100
rect 6066 1098 6068 1100
rect 6072 1098 6074 1100
rect 6096 1098 6098 1100
rect 6102 1098 6104 1100
rect 6126 1098 6128 1100
rect 6132 1098 6134 1100
rect 6250 1099 6252 1100
rect 6748 1099 6750 1100
rect 3248 1097 3250 1098
rect 3750 1097 3752 1098
rect 3848 1097 3850 1098
rect 4350 1097 4352 1098
rect 4474 1096 4476 1098
rect 4504 1096 4506 1098
rect 4534 1096 4536 1098
rect 4564 1096 4566 1098
rect 4594 1096 4596 1098
rect 4624 1096 4626 1098
rect 4654 1096 4656 1098
rect 4684 1096 4686 1098
rect 4714 1096 4716 1098
rect 4744 1096 4746 1098
rect 4774 1096 4776 1098
rect 4804 1096 4806 1098
rect 4834 1096 4836 1098
rect 4864 1096 4866 1098
rect 4894 1096 4896 1098
rect 4924 1096 4926 1098
rect 5074 1096 5076 1098
rect 5104 1096 5106 1098
rect 5134 1096 5136 1098
rect 5164 1096 5166 1098
rect 5194 1096 5196 1098
rect 5224 1096 5226 1098
rect 5254 1096 5256 1098
rect 5284 1096 5286 1098
rect 5314 1096 5316 1098
rect 5344 1096 5346 1098
rect 5374 1096 5376 1098
rect 5404 1096 5406 1098
rect 5434 1096 5436 1098
rect 5464 1096 5466 1098
rect 5494 1096 5496 1098
rect 5524 1096 5526 1098
rect 5674 1096 5676 1098
rect 5704 1096 5706 1098
rect 5734 1096 5736 1098
rect 5764 1096 5766 1098
rect 5794 1096 5796 1098
rect 5824 1096 5826 1098
rect 5854 1096 5856 1098
rect 5884 1096 5886 1098
rect 5914 1096 5916 1098
rect 5944 1096 5946 1098
rect 5974 1096 5976 1098
rect 6004 1096 6006 1098
rect 6034 1096 6036 1098
rect 6064 1096 6066 1098
rect 6094 1096 6096 1098
rect 6124 1096 6126 1098
rect 6248 1097 6250 1098
rect 6750 1097 6752 1098
rect 4474 1090 4476 1092
rect 4504 1090 4506 1092
rect 4534 1090 4536 1092
rect 4564 1090 4566 1092
rect 4594 1090 4596 1092
rect 4624 1090 4626 1092
rect 4654 1090 4656 1092
rect 4684 1090 4686 1092
rect 4714 1090 4716 1092
rect 4744 1090 4746 1092
rect 4774 1090 4776 1092
rect 4804 1090 4806 1092
rect 4834 1090 4836 1092
rect 4864 1090 4866 1092
rect 4894 1090 4896 1092
rect 4924 1090 4926 1092
rect 5074 1090 5076 1092
rect 5104 1090 5106 1092
rect 5134 1090 5136 1092
rect 5164 1090 5166 1092
rect 5194 1090 5196 1092
rect 5224 1090 5226 1092
rect 5254 1090 5256 1092
rect 5284 1090 5286 1092
rect 5314 1090 5316 1092
rect 5344 1090 5346 1092
rect 5374 1090 5376 1092
rect 5404 1090 5406 1092
rect 5434 1090 5436 1092
rect 5464 1090 5466 1092
rect 5494 1090 5496 1092
rect 5524 1090 5526 1092
rect 5674 1090 5676 1092
rect 5704 1090 5706 1092
rect 5734 1090 5736 1092
rect 5764 1090 5766 1092
rect 5794 1090 5796 1092
rect 5824 1090 5826 1092
rect 5854 1090 5856 1092
rect 5884 1090 5886 1092
rect 5914 1090 5916 1092
rect 5944 1090 5946 1092
rect 5974 1090 5976 1092
rect 6004 1090 6006 1092
rect 6034 1090 6036 1092
rect 6064 1090 6066 1092
rect 6094 1090 6096 1092
rect 6124 1090 6126 1092
rect 4476 1088 4478 1090
rect 4482 1088 4484 1090
rect 4506 1088 4508 1090
rect 4512 1088 4514 1090
rect 4536 1088 4538 1090
rect 4542 1088 4544 1090
rect 4566 1088 4568 1090
rect 4572 1088 4574 1090
rect 4596 1088 4598 1090
rect 4602 1088 4604 1090
rect 4626 1088 4628 1090
rect 4632 1088 4634 1090
rect 4656 1088 4658 1090
rect 4662 1088 4664 1090
rect 4686 1088 4688 1090
rect 4692 1088 4694 1090
rect 4716 1088 4718 1090
rect 4722 1088 4724 1090
rect 4746 1088 4748 1090
rect 4752 1088 4754 1090
rect 4776 1088 4778 1090
rect 4782 1088 4784 1090
rect 4806 1088 4808 1090
rect 4812 1088 4814 1090
rect 4836 1088 4838 1090
rect 4842 1088 4844 1090
rect 4866 1088 4868 1090
rect 4872 1088 4874 1090
rect 4896 1088 4898 1090
rect 4902 1088 4904 1090
rect 4926 1088 4928 1090
rect 4932 1088 4934 1090
rect 5076 1088 5078 1090
rect 5082 1088 5084 1090
rect 5106 1088 5108 1090
rect 5112 1088 5114 1090
rect 5136 1088 5138 1090
rect 5142 1088 5144 1090
rect 5166 1088 5168 1090
rect 5172 1088 5174 1090
rect 5196 1088 5198 1090
rect 5202 1088 5204 1090
rect 5226 1088 5228 1090
rect 5232 1088 5234 1090
rect 5256 1088 5258 1090
rect 5262 1088 5264 1090
rect 5286 1088 5288 1090
rect 5292 1088 5294 1090
rect 5316 1088 5318 1090
rect 5322 1088 5324 1090
rect 5346 1088 5348 1090
rect 5352 1088 5354 1090
rect 5376 1088 5378 1090
rect 5382 1088 5384 1090
rect 5406 1088 5408 1090
rect 5412 1088 5414 1090
rect 5436 1088 5438 1090
rect 5442 1088 5444 1090
rect 5466 1088 5468 1090
rect 5472 1088 5474 1090
rect 5496 1088 5498 1090
rect 5502 1088 5504 1090
rect 5526 1088 5528 1090
rect 5532 1088 5534 1090
rect 5676 1088 5678 1090
rect 5682 1088 5684 1090
rect 5706 1088 5708 1090
rect 5712 1088 5714 1090
rect 5736 1088 5738 1090
rect 5742 1088 5744 1090
rect 5766 1088 5768 1090
rect 5772 1088 5774 1090
rect 5796 1088 5798 1090
rect 5802 1088 5804 1090
rect 5826 1088 5828 1090
rect 5832 1088 5834 1090
rect 5856 1088 5858 1090
rect 5862 1088 5864 1090
rect 5886 1088 5888 1090
rect 5892 1088 5894 1090
rect 5916 1088 5918 1090
rect 5922 1088 5924 1090
rect 5946 1088 5948 1090
rect 5952 1088 5954 1090
rect 5976 1088 5978 1090
rect 5982 1088 5984 1090
rect 6006 1088 6008 1090
rect 6012 1088 6014 1090
rect 6036 1088 6038 1090
rect 6042 1088 6044 1090
rect 6066 1088 6068 1090
rect 6072 1088 6074 1090
rect 6096 1088 6098 1090
rect 6102 1088 6104 1090
rect 6126 1088 6128 1090
rect 6132 1088 6134 1090
rect 4484 1086 4486 1088
rect 4514 1086 4516 1088
rect 4544 1086 4546 1088
rect 4574 1086 4576 1088
rect 4604 1086 4606 1088
rect 4634 1086 4636 1088
rect 4664 1086 4666 1088
rect 4694 1086 4696 1088
rect 4724 1086 4726 1088
rect 4754 1086 4756 1088
rect 4784 1086 4786 1088
rect 4814 1086 4816 1088
rect 4844 1086 4846 1088
rect 4874 1086 4876 1088
rect 4904 1086 4906 1088
rect 4934 1086 4936 1088
rect 5084 1086 5086 1088
rect 5114 1086 5116 1088
rect 5144 1086 5146 1088
rect 5174 1086 5176 1088
rect 5204 1086 5206 1088
rect 5234 1086 5236 1088
rect 5264 1086 5266 1088
rect 5294 1086 5296 1088
rect 5324 1086 5326 1088
rect 5354 1086 5356 1088
rect 5384 1086 5386 1088
rect 5414 1086 5416 1088
rect 5444 1086 5446 1088
rect 5474 1086 5476 1088
rect 5504 1086 5506 1088
rect 5534 1086 5536 1088
rect 5684 1086 5686 1088
rect 5714 1086 5716 1088
rect 5744 1086 5746 1088
rect 5774 1086 5776 1088
rect 5804 1086 5806 1088
rect 5834 1086 5836 1088
rect 5864 1086 5866 1088
rect 5894 1086 5896 1088
rect 5924 1086 5926 1088
rect 5954 1086 5956 1088
rect 5984 1086 5986 1088
rect 6014 1086 6016 1088
rect 6044 1086 6046 1088
rect 6074 1086 6076 1088
rect 6104 1086 6106 1088
rect 6134 1086 6136 1088
rect 4484 1080 4486 1082
rect 4514 1080 4516 1082
rect 4544 1080 4546 1082
rect 4574 1080 4576 1082
rect 4604 1080 4606 1082
rect 4634 1080 4636 1082
rect 4664 1080 4666 1082
rect 4694 1080 4696 1082
rect 4724 1080 4726 1082
rect 4754 1080 4756 1082
rect 4784 1080 4786 1082
rect 4814 1080 4816 1082
rect 4844 1080 4846 1082
rect 4874 1080 4876 1082
rect 4904 1080 4906 1082
rect 4934 1080 4936 1082
rect 5084 1080 5086 1082
rect 5114 1080 5116 1082
rect 5144 1080 5146 1082
rect 5174 1080 5176 1082
rect 5204 1080 5206 1082
rect 5234 1080 5236 1082
rect 5264 1080 5266 1082
rect 5294 1080 5296 1082
rect 5324 1080 5326 1082
rect 5354 1080 5356 1082
rect 5384 1080 5386 1082
rect 5414 1080 5416 1082
rect 5444 1080 5446 1082
rect 5474 1080 5476 1082
rect 5504 1080 5506 1082
rect 5534 1080 5536 1082
rect 5684 1080 5686 1082
rect 5714 1080 5716 1082
rect 5744 1080 5746 1082
rect 5774 1080 5776 1082
rect 5804 1080 5806 1082
rect 5834 1080 5836 1082
rect 5864 1080 5866 1082
rect 5894 1080 5896 1082
rect 5924 1080 5926 1082
rect 5954 1080 5956 1082
rect 5984 1080 5986 1082
rect 6014 1080 6016 1082
rect 6044 1080 6046 1082
rect 6074 1080 6076 1082
rect 6104 1080 6106 1082
rect 6134 1080 6136 1082
rect 3250 1079 3252 1080
rect 3748 1079 3750 1080
rect 3850 1079 3852 1080
rect 4348 1079 4350 1080
rect 4476 1078 4478 1080
rect 4482 1078 4484 1080
rect 4506 1078 4508 1080
rect 4512 1078 4514 1080
rect 4536 1078 4538 1080
rect 4542 1078 4544 1080
rect 4566 1078 4568 1080
rect 4572 1078 4574 1080
rect 4596 1078 4598 1080
rect 4602 1078 4604 1080
rect 4626 1078 4628 1080
rect 4632 1078 4634 1080
rect 4656 1078 4658 1080
rect 4662 1078 4664 1080
rect 4686 1078 4688 1080
rect 4692 1078 4694 1080
rect 4716 1078 4718 1080
rect 4722 1078 4724 1080
rect 4746 1078 4748 1080
rect 4752 1078 4754 1080
rect 4776 1078 4778 1080
rect 4782 1078 4784 1080
rect 4806 1078 4808 1080
rect 4812 1078 4814 1080
rect 4836 1078 4838 1080
rect 4842 1078 4844 1080
rect 4866 1078 4868 1080
rect 4872 1078 4874 1080
rect 4896 1078 4898 1080
rect 4902 1078 4904 1080
rect 4926 1078 4928 1080
rect 4932 1078 4934 1080
rect 5076 1078 5078 1080
rect 5082 1078 5084 1080
rect 5106 1078 5108 1080
rect 5112 1078 5114 1080
rect 5136 1078 5138 1080
rect 5142 1078 5144 1080
rect 5166 1078 5168 1080
rect 5172 1078 5174 1080
rect 5196 1078 5198 1080
rect 5202 1078 5204 1080
rect 5226 1078 5228 1080
rect 5232 1078 5234 1080
rect 5256 1078 5258 1080
rect 5262 1078 5264 1080
rect 5286 1078 5288 1080
rect 5292 1078 5294 1080
rect 5316 1078 5318 1080
rect 5322 1078 5324 1080
rect 5346 1078 5348 1080
rect 5352 1078 5354 1080
rect 5376 1078 5378 1080
rect 5382 1078 5384 1080
rect 5406 1078 5408 1080
rect 5412 1078 5414 1080
rect 5436 1078 5438 1080
rect 5442 1078 5444 1080
rect 5466 1078 5468 1080
rect 5472 1078 5474 1080
rect 5496 1078 5498 1080
rect 5502 1078 5504 1080
rect 5526 1078 5528 1080
rect 5532 1078 5534 1080
rect 5676 1078 5678 1080
rect 5682 1078 5684 1080
rect 5706 1078 5708 1080
rect 5712 1078 5714 1080
rect 5736 1078 5738 1080
rect 5742 1078 5744 1080
rect 5766 1078 5768 1080
rect 5772 1078 5774 1080
rect 5796 1078 5798 1080
rect 5802 1078 5804 1080
rect 5826 1078 5828 1080
rect 5832 1078 5834 1080
rect 5856 1078 5858 1080
rect 5862 1078 5864 1080
rect 5886 1078 5888 1080
rect 5892 1078 5894 1080
rect 5916 1078 5918 1080
rect 5922 1078 5924 1080
rect 5946 1078 5948 1080
rect 5952 1078 5954 1080
rect 5976 1078 5978 1080
rect 5982 1078 5984 1080
rect 6006 1078 6008 1080
rect 6012 1078 6014 1080
rect 6036 1078 6038 1080
rect 6042 1078 6044 1080
rect 6066 1078 6068 1080
rect 6072 1078 6074 1080
rect 6096 1078 6098 1080
rect 6102 1078 6104 1080
rect 6126 1078 6128 1080
rect 6132 1078 6134 1080
rect 6250 1079 6252 1080
rect 6748 1079 6750 1080
rect 3248 1077 3250 1078
rect 3750 1077 3752 1078
rect 3848 1077 3850 1078
rect 4350 1077 4352 1078
rect 4474 1076 4476 1078
rect 4504 1076 4506 1078
rect 4534 1076 4536 1078
rect 4564 1076 4566 1078
rect 4594 1076 4596 1078
rect 4624 1076 4626 1078
rect 4654 1076 4656 1078
rect 4684 1076 4686 1078
rect 4714 1076 4716 1078
rect 4744 1076 4746 1078
rect 4774 1076 4776 1078
rect 4804 1076 4806 1078
rect 4834 1076 4836 1078
rect 4864 1076 4866 1078
rect 4894 1076 4896 1078
rect 4924 1076 4926 1078
rect 5074 1076 5076 1078
rect 5104 1076 5106 1078
rect 5134 1076 5136 1078
rect 5164 1076 5166 1078
rect 5194 1076 5196 1078
rect 5224 1076 5226 1078
rect 5254 1076 5256 1078
rect 5284 1076 5286 1078
rect 5314 1076 5316 1078
rect 5344 1076 5346 1078
rect 5374 1076 5376 1078
rect 5404 1076 5406 1078
rect 5434 1076 5436 1078
rect 5464 1076 5466 1078
rect 5494 1076 5496 1078
rect 5524 1076 5526 1078
rect 5674 1076 5676 1078
rect 5704 1076 5706 1078
rect 5734 1076 5736 1078
rect 5764 1076 5766 1078
rect 5794 1076 5796 1078
rect 5824 1076 5826 1078
rect 5854 1076 5856 1078
rect 5884 1076 5886 1078
rect 5914 1076 5916 1078
rect 5944 1076 5946 1078
rect 5974 1076 5976 1078
rect 6004 1076 6006 1078
rect 6034 1076 6036 1078
rect 6064 1076 6066 1078
rect 6094 1076 6096 1078
rect 6124 1076 6126 1078
rect 6248 1077 6250 1078
rect 6750 1077 6752 1078
rect 4474 1070 4476 1072
rect 4504 1070 4506 1072
rect 4534 1070 4536 1072
rect 4564 1070 4566 1072
rect 4594 1070 4596 1072
rect 4624 1070 4626 1072
rect 4654 1070 4656 1072
rect 4684 1070 4686 1072
rect 4714 1070 4716 1072
rect 4744 1070 4746 1072
rect 4774 1070 4776 1072
rect 4804 1070 4806 1072
rect 4834 1070 4836 1072
rect 4864 1070 4866 1072
rect 4894 1070 4896 1072
rect 4924 1070 4926 1072
rect 5074 1070 5076 1072
rect 5104 1070 5106 1072
rect 5134 1070 5136 1072
rect 5164 1070 5166 1072
rect 5194 1070 5196 1072
rect 5224 1070 5226 1072
rect 5254 1070 5256 1072
rect 5284 1070 5286 1072
rect 5314 1070 5316 1072
rect 5344 1070 5346 1072
rect 5374 1070 5376 1072
rect 5404 1070 5406 1072
rect 5434 1070 5436 1072
rect 5464 1070 5466 1072
rect 5494 1070 5496 1072
rect 5524 1070 5526 1072
rect 5674 1070 5676 1072
rect 5704 1070 5706 1072
rect 5734 1070 5736 1072
rect 5764 1070 5766 1072
rect 5794 1070 5796 1072
rect 5824 1070 5826 1072
rect 5854 1070 5856 1072
rect 5884 1070 5886 1072
rect 5914 1070 5916 1072
rect 5944 1070 5946 1072
rect 5974 1070 5976 1072
rect 6004 1070 6006 1072
rect 6034 1070 6036 1072
rect 6064 1070 6066 1072
rect 6094 1070 6096 1072
rect 6124 1070 6126 1072
rect 4476 1068 4478 1070
rect 4482 1068 4484 1070
rect 4506 1068 4508 1070
rect 4512 1068 4514 1070
rect 4536 1068 4538 1070
rect 4542 1068 4544 1070
rect 4566 1068 4568 1070
rect 4572 1068 4574 1070
rect 4596 1068 4598 1070
rect 4602 1068 4604 1070
rect 4626 1068 4628 1070
rect 4632 1068 4634 1070
rect 4656 1068 4658 1070
rect 4662 1068 4664 1070
rect 4686 1068 4688 1070
rect 4692 1068 4694 1070
rect 4716 1068 4718 1070
rect 4722 1068 4724 1070
rect 4746 1068 4748 1070
rect 4752 1068 4754 1070
rect 4776 1068 4778 1070
rect 4782 1068 4784 1070
rect 4806 1068 4808 1070
rect 4812 1068 4814 1070
rect 4836 1068 4838 1070
rect 4842 1068 4844 1070
rect 4866 1068 4868 1070
rect 4872 1068 4874 1070
rect 4896 1068 4898 1070
rect 4902 1068 4904 1070
rect 4926 1068 4928 1070
rect 4932 1068 4934 1070
rect 5076 1068 5078 1070
rect 5082 1068 5084 1070
rect 5106 1068 5108 1070
rect 5112 1068 5114 1070
rect 5136 1068 5138 1070
rect 5142 1068 5144 1070
rect 5166 1068 5168 1070
rect 5172 1068 5174 1070
rect 5196 1068 5198 1070
rect 5202 1068 5204 1070
rect 5226 1068 5228 1070
rect 5232 1068 5234 1070
rect 5256 1068 5258 1070
rect 5262 1068 5264 1070
rect 5286 1068 5288 1070
rect 5292 1068 5294 1070
rect 5316 1068 5318 1070
rect 5322 1068 5324 1070
rect 5346 1068 5348 1070
rect 5352 1068 5354 1070
rect 5376 1068 5378 1070
rect 5382 1068 5384 1070
rect 5406 1068 5408 1070
rect 5412 1068 5414 1070
rect 5436 1068 5438 1070
rect 5442 1068 5444 1070
rect 5466 1068 5468 1070
rect 5472 1068 5474 1070
rect 5496 1068 5498 1070
rect 5502 1068 5504 1070
rect 5526 1068 5528 1070
rect 5532 1068 5534 1070
rect 5676 1068 5678 1070
rect 5682 1068 5684 1070
rect 5706 1068 5708 1070
rect 5712 1068 5714 1070
rect 5736 1068 5738 1070
rect 5742 1068 5744 1070
rect 5766 1068 5768 1070
rect 5772 1068 5774 1070
rect 5796 1068 5798 1070
rect 5802 1068 5804 1070
rect 5826 1068 5828 1070
rect 5832 1068 5834 1070
rect 5856 1068 5858 1070
rect 5862 1068 5864 1070
rect 5886 1068 5888 1070
rect 5892 1068 5894 1070
rect 5916 1068 5918 1070
rect 5922 1068 5924 1070
rect 5946 1068 5948 1070
rect 5952 1068 5954 1070
rect 5976 1068 5978 1070
rect 5982 1068 5984 1070
rect 6006 1068 6008 1070
rect 6012 1068 6014 1070
rect 6036 1068 6038 1070
rect 6042 1068 6044 1070
rect 6066 1068 6068 1070
rect 6072 1068 6074 1070
rect 6096 1068 6098 1070
rect 6102 1068 6104 1070
rect 6126 1068 6128 1070
rect 6132 1068 6134 1070
rect 4484 1066 4486 1068
rect 4514 1066 4516 1068
rect 4544 1066 4546 1068
rect 4574 1066 4576 1068
rect 4604 1066 4606 1068
rect 4634 1066 4636 1068
rect 4664 1066 4666 1068
rect 4694 1066 4696 1068
rect 4724 1066 4726 1068
rect 4754 1066 4756 1068
rect 4784 1066 4786 1068
rect 4814 1066 4816 1068
rect 4844 1066 4846 1068
rect 4874 1066 4876 1068
rect 4904 1066 4906 1068
rect 4934 1066 4936 1068
rect 5084 1066 5086 1068
rect 5114 1066 5116 1068
rect 5144 1066 5146 1068
rect 5174 1066 5176 1068
rect 5204 1066 5206 1068
rect 5234 1066 5236 1068
rect 5264 1066 5266 1068
rect 5294 1066 5296 1068
rect 5324 1066 5326 1068
rect 5354 1066 5356 1068
rect 5384 1066 5386 1068
rect 5414 1066 5416 1068
rect 5444 1066 5446 1068
rect 5474 1066 5476 1068
rect 5504 1066 5506 1068
rect 5534 1066 5536 1068
rect 5684 1066 5686 1068
rect 5714 1066 5716 1068
rect 5744 1066 5746 1068
rect 5774 1066 5776 1068
rect 5804 1066 5806 1068
rect 5834 1066 5836 1068
rect 5864 1066 5866 1068
rect 5894 1066 5896 1068
rect 5924 1066 5926 1068
rect 5954 1066 5956 1068
rect 5984 1066 5986 1068
rect 6014 1066 6016 1068
rect 6044 1066 6046 1068
rect 6074 1066 6076 1068
rect 6104 1066 6106 1068
rect 6134 1066 6136 1068
rect 4484 1060 4486 1062
rect 4514 1060 4516 1062
rect 4544 1060 4546 1062
rect 4574 1060 4576 1062
rect 4604 1060 4606 1062
rect 4634 1060 4636 1062
rect 4664 1060 4666 1062
rect 4694 1060 4696 1062
rect 4724 1060 4726 1062
rect 4754 1060 4756 1062
rect 4784 1060 4786 1062
rect 4814 1060 4816 1062
rect 4844 1060 4846 1062
rect 4874 1060 4876 1062
rect 4904 1060 4906 1062
rect 4934 1060 4936 1062
rect 5084 1060 5086 1062
rect 5114 1060 5116 1062
rect 5144 1060 5146 1062
rect 5174 1060 5176 1062
rect 5204 1060 5206 1062
rect 5234 1060 5236 1062
rect 5264 1060 5266 1062
rect 5294 1060 5296 1062
rect 5324 1060 5326 1062
rect 5354 1060 5356 1062
rect 5384 1060 5386 1062
rect 5414 1060 5416 1062
rect 5444 1060 5446 1062
rect 5474 1060 5476 1062
rect 5504 1060 5506 1062
rect 5534 1060 5536 1062
rect 5684 1060 5686 1062
rect 5714 1060 5716 1062
rect 5744 1060 5746 1062
rect 5774 1060 5776 1062
rect 5804 1060 5806 1062
rect 5834 1060 5836 1062
rect 5864 1060 5866 1062
rect 5894 1060 5896 1062
rect 5924 1060 5926 1062
rect 5954 1060 5956 1062
rect 5984 1060 5986 1062
rect 6014 1060 6016 1062
rect 6044 1060 6046 1062
rect 6074 1060 6076 1062
rect 6104 1060 6106 1062
rect 6134 1060 6136 1062
rect 3250 1059 3252 1060
rect 3748 1059 3750 1060
rect 3850 1059 3852 1060
rect 4348 1059 4350 1060
rect 4476 1058 4478 1060
rect 4482 1058 4484 1060
rect 4506 1058 4508 1060
rect 4512 1058 4514 1060
rect 4536 1058 4538 1060
rect 4542 1058 4544 1060
rect 4566 1058 4568 1060
rect 4572 1058 4574 1060
rect 4596 1058 4598 1060
rect 4602 1058 4604 1060
rect 4626 1058 4628 1060
rect 4632 1058 4634 1060
rect 4656 1058 4658 1060
rect 4662 1058 4664 1060
rect 4686 1058 4688 1060
rect 4692 1058 4694 1060
rect 4716 1058 4718 1060
rect 4722 1058 4724 1060
rect 4746 1058 4748 1060
rect 4752 1058 4754 1060
rect 4776 1058 4778 1060
rect 4782 1058 4784 1060
rect 4806 1058 4808 1060
rect 4812 1058 4814 1060
rect 4836 1058 4838 1060
rect 4842 1058 4844 1060
rect 4866 1058 4868 1060
rect 4872 1058 4874 1060
rect 4896 1058 4898 1060
rect 4902 1058 4904 1060
rect 4926 1058 4928 1060
rect 4932 1058 4934 1060
rect 5076 1058 5078 1060
rect 5082 1058 5084 1060
rect 5106 1058 5108 1060
rect 5112 1058 5114 1060
rect 5136 1058 5138 1060
rect 5142 1058 5144 1060
rect 5166 1058 5168 1060
rect 5172 1058 5174 1060
rect 5196 1058 5198 1060
rect 5202 1058 5204 1060
rect 5226 1058 5228 1060
rect 5232 1058 5234 1060
rect 5256 1058 5258 1060
rect 5262 1058 5264 1060
rect 5286 1058 5288 1060
rect 5292 1058 5294 1060
rect 5316 1058 5318 1060
rect 5322 1058 5324 1060
rect 5346 1058 5348 1060
rect 5352 1058 5354 1060
rect 5376 1058 5378 1060
rect 5382 1058 5384 1060
rect 5406 1058 5408 1060
rect 5412 1058 5414 1060
rect 5436 1058 5438 1060
rect 5442 1058 5444 1060
rect 5466 1058 5468 1060
rect 5472 1058 5474 1060
rect 5496 1058 5498 1060
rect 5502 1058 5504 1060
rect 5526 1058 5528 1060
rect 5532 1058 5534 1060
rect 5676 1058 5678 1060
rect 5682 1058 5684 1060
rect 5706 1058 5708 1060
rect 5712 1058 5714 1060
rect 5736 1058 5738 1060
rect 5742 1058 5744 1060
rect 5766 1058 5768 1060
rect 5772 1058 5774 1060
rect 5796 1058 5798 1060
rect 5802 1058 5804 1060
rect 5826 1058 5828 1060
rect 5832 1058 5834 1060
rect 5856 1058 5858 1060
rect 5862 1058 5864 1060
rect 5886 1058 5888 1060
rect 5892 1058 5894 1060
rect 5916 1058 5918 1060
rect 5922 1058 5924 1060
rect 5946 1058 5948 1060
rect 5952 1058 5954 1060
rect 5976 1058 5978 1060
rect 5982 1058 5984 1060
rect 6006 1058 6008 1060
rect 6012 1058 6014 1060
rect 6036 1058 6038 1060
rect 6042 1058 6044 1060
rect 6066 1058 6068 1060
rect 6072 1058 6074 1060
rect 6096 1058 6098 1060
rect 6102 1058 6104 1060
rect 6126 1058 6128 1060
rect 6132 1058 6134 1060
rect 6250 1059 6252 1060
rect 6748 1059 6750 1060
rect 3248 1057 3250 1058
rect 3750 1057 3752 1058
rect 3848 1057 3850 1058
rect 4350 1057 4352 1058
rect 4474 1056 4476 1058
rect 4504 1056 4506 1058
rect 4534 1056 4536 1058
rect 4564 1056 4566 1058
rect 4594 1056 4596 1058
rect 4624 1056 4626 1058
rect 4654 1056 4656 1058
rect 4684 1056 4686 1058
rect 4714 1056 4716 1058
rect 4744 1056 4746 1058
rect 4774 1056 4776 1058
rect 4804 1056 4806 1058
rect 4834 1056 4836 1058
rect 4864 1056 4866 1058
rect 4894 1056 4896 1058
rect 4924 1056 4926 1058
rect 5074 1056 5076 1058
rect 5104 1056 5106 1058
rect 5134 1056 5136 1058
rect 5164 1056 5166 1058
rect 5194 1056 5196 1058
rect 5224 1056 5226 1058
rect 5254 1056 5256 1058
rect 5284 1056 5286 1058
rect 5314 1056 5316 1058
rect 5344 1056 5346 1058
rect 5374 1056 5376 1058
rect 5404 1056 5406 1058
rect 5434 1056 5436 1058
rect 5464 1056 5466 1058
rect 5494 1056 5496 1058
rect 5524 1056 5526 1058
rect 5674 1056 5676 1058
rect 5704 1056 5706 1058
rect 5734 1056 5736 1058
rect 5764 1056 5766 1058
rect 5794 1056 5796 1058
rect 5824 1056 5826 1058
rect 5854 1056 5856 1058
rect 5884 1056 5886 1058
rect 5914 1056 5916 1058
rect 5944 1056 5946 1058
rect 5974 1056 5976 1058
rect 6004 1056 6006 1058
rect 6034 1056 6036 1058
rect 6064 1056 6066 1058
rect 6094 1056 6096 1058
rect 6124 1056 6126 1058
rect 6248 1057 6250 1058
rect 6750 1057 6752 1058
rect 3294 1052 3296 1054
rect 3704 1052 3706 1054
rect 3894 1052 3896 1054
rect 4304 1052 4306 1054
rect 6294 1052 6296 1054
rect 6704 1052 6706 1054
rect 3296 1050 3298 1052
rect 3702 1050 3704 1052
rect 3896 1050 3898 1052
rect 4302 1050 4304 1052
rect 4474 1050 4476 1052
rect 4504 1050 4506 1052
rect 4534 1050 4536 1052
rect 4564 1050 4566 1052
rect 4594 1050 4596 1052
rect 4624 1050 4626 1052
rect 4654 1050 4656 1052
rect 4684 1050 4686 1052
rect 4714 1050 4716 1052
rect 4744 1050 4746 1052
rect 4774 1050 4776 1052
rect 4804 1050 4806 1052
rect 4834 1050 4836 1052
rect 4864 1050 4866 1052
rect 4894 1050 4896 1052
rect 4924 1050 4926 1052
rect 5074 1050 5076 1052
rect 5104 1050 5106 1052
rect 5134 1050 5136 1052
rect 5164 1050 5166 1052
rect 5194 1050 5196 1052
rect 5224 1050 5226 1052
rect 5254 1050 5256 1052
rect 5284 1050 5286 1052
rect 5314 1050 5316 1052
rect 5344 1050 5346 1052
rect 5374 1050 5376 1052
rect 5404 1050 5406 1052
rect 5434 1050 5436 1052
rect 5464 1050 5466 1052
rect 5494 1050 5496 1052
rect 5524 1050 5526 1052
rect 5674 1050 5676 1052
rect 5704 1050 5706 1052
rect 5734 1050 5736 1052
rect 5764 1050 5766 1052
rect 5794 1050 5796 1052
rect 5824 1050 5826 1052
rect 5854 1050 5856 1052
rect 5884 1050 5886 1052
rect 5914 1050 5916 1052
rect 5944 1050 5946 1052
rect 5974 1050 5976 1052
rect 6004 1050 6006 1052
rect 6034 1050 6036 1052
rect 6064 1050 6066 1052
rect 6094 1050 6096 1052
rect 6124 1050 6126 1052
rect 6296 1050 6298 1052
rect 6702 1050 6704 1052
rect 4476 1048 4478 1050
rect 4482 1048 4484 1050
rect 4506 1048 4508 1050
rect 4512 1048 4514 1050
rect 4536 1048 4538 1050
rect 4542 1048 4544 1050
rect 4566 1048 4568 1050
rect 4572 1048 4574 1050
rect 4596 1048 4598 1050
rect 4602 1048 4604 1050
rect 4626 1048 4628 1050
rect 4632 1048 4634 1050
rect 4656 1048 4658 1050
rect 4662 1048 4664 1050
rect 4686 1048 4688 1050
rect 4692 1048 4694 1050
rect 4716 1048 4718 1050
rect 4722 1048 4724 1050
rect 4746 1048 4748 1050
rect 4752 1048 4754 1050
rect 4776 1048 4778 1050
rect 4782 1048 4784 1050
rect 4806 1048 4808 1050
rect 4812 1048 4814 1050
rect 4836 1048 4838 1050
rect 4842 1048 4844 1050
rect 4866 1048 4868 1050
rect 4872 1048 4874 1050
rect 4896 1048 4898 1050
rect 4902 1048 4904 1050
rect 4926 1048 4928 1050
rect 4932 1048 4934 1050
rect 5076 1048 5078 1050
rect 5082 1048 5084 1050
rect 5106 1048 5108 1050
rect 5112 1048 5114 1050
rect 5136 1048 5138 1050
rect 5142 1048 5144 1050
rect 5166 1048 5168 1050
rect 5172 1048 5174 1050
rect 5196 1048 5198 1050
rect 5202 1048 5204 1050
rect 5226 1048 5228 1050
rect 5232 1048 5234 1050
rect 5256 1048 5258 1050
rect 5262 1048 5264 1050
rect 5286 1048 5288 1050
rect 5292 1048 5294 1050
rect 5316 1048 5318 1050
rect 5322 1048 5324 1050
rect 5346 1048 5348 1050
rect 5352 1048 5354 1050
rect 5376 1048 5378 1050
rect 5382 1048 5384 1050
rect 5406 1048 5408 1050
rect 5412 1048 5414 1050
rect 5436 1048 5438 1050
rect 5442 1048 5444 1050
rect 5466 1048 5468 1050
rect 5472 1048 5474 1050
rect 5496 1048 5498 1050
rect 5502 1048 5504 1050
rect 5526 1048 5528 1050
rect 5532 1048 5534 1050
rect 5676 1048 5678 1050
rect 5682 1048 5684 1050
rect 5706 1048 5708 1050
rect 5712 1048 5714 1050
rect 5736 1048 5738 1050
rect 5742 1048 5744 1050
rect 5766 1048 5768 1050
rect 5772 1048 5774 1050
rect 5796 1048 5798 1050
rect 5802 1048 5804 1050
rect 5826 1048 5828 1050
rect 5832 1048 5834 1050
rect 5856 1048 5858 1050
rect 5862 1048 5864 1050
rect 5886 1048 5888 1050
rect 5892 1048 5894 1050
rect 5916 1048 5918 1050
rect 5922 1048 5924 1050
rect 5946 1048 5948 1050
rect 5952 1048 5954 1050
rect 5976 1048 5978 1050
rect 5982 1048 5984 1050
rect 6006 1048 6008 1050
rect 6012 1048 6014 1050
rect 6036 1048 6038 1050
rect 6042 1048 6044 1050
rect 6066 1048 6068 1050
rect 6072 1048 6074 1050
rect 6096 1048 6098 1050
rect 6102 1048 6104 1050
rect 6126 1048 6128 1050
rect 6132 1048 6134 1050
rect 4484 1046 4486 1048
rect 4514 1046 4516 1048
rect 4544 1046 4546 1048
rect 4574 1046 4576 1048
rect 4604 1046 4606 1048
rect 4634 1046 4636 1048
rect 4664 1046 4666 1048
rect 4694 1046 4696 1048
rect 4724 1046 4726 1048
rect 4754 1046 4756 1048
rect 4784 1046 4786 1048
rect 4814 1046 4816 1048
rect 4844 1046 4846 1048
rect 4874 1046 4876 1048
rect 4904 1046 4906 1048
rect 4934 1046 4936 1048
rect 5084 1046 5086 1048
rect 5114 1046 5116 1048
rect 5144 1046 5146 1048
rect 5174 1046 5176 1048
rect 5204 1046 5206 1048
rect 5234 1046 5236 1048
rect 5264 1046 5266 1048
rect 5294 1046 5296 1048
rect 5324 1046 5326 1048
rect 5354 1046 5356 1048
rect 5384 1046 5386 1048
rect 5414 1046 5416 1048
rect 5444 1046 5446 1048
rect 5474 1046 5476 1048
rect 5504 1046 5506 1048
rect 5534 1046 5536 1048
rect 5684 1046 5686 1048
rect 5714 1046 5716 1048
rect 5744 1046 5746 1048
rect 5774 1046 5776 1048
rect 5804 1046 5806 1048
rect 5834 1046 5836 1048
rect 5864 1046 5866 1048
rect 5894 1046 5896 1048
rect 5924 1046 5926 1048
rect 5954 1046 5956 1048
rect 5984 1046 5986 1048
rect 6014 1046 6016 1048
rect 6044 1046 6046 1048
rect 6074 1046 6076 1048
rect 6104 1046 6106 1048
rect 6134 1046 6136 1048
rect 4484 1040 4486 1042
rect 4904 1040 4906 1042
rect 4934 1040 4936 1042
rect 5084 1040 5086 1042
rect 5504 1040 5506 1042
rect 5534 1040 5536 1042
rect 5684 1040 5686 1042
rect 6104 1040 6106 1042
rect 6134 1040 6136 1042
rect 3250 1039 3252 1040
rect 3748 1039 3750 1040
rect 3850 1039 3852 1040
rect 4348 1039 4350 1040
rect 4476 1038 4478 1040
rect 4482 1038 4484 1040
rect 4906 1038 4908 1040
rect 4932 1038 4934 1040
rect 5076 1038 5078 1040
rect 5082 1038 5084 1040
rect 5506 1038 5508 1040
rect 5532 1038 5534 1040
rect 5676 1038 5678 1040
rect 5682 1038 5684 1040
rect 6106 1038 6108 1040
rect 6132 1038 6134 1040
rect 6250 1039 6252 1040
rect 6748 1039 6750 1040
rect 3248 1037 3250 1038
rect 3750 1037 3752 1038
rect 3848 1037 3850 1038
rect 4350 1037 4352 1038
rect 4474 1036 4476 1038
rect 5074 1036 5076 1038
rect 5674 1036 5676 1038
rect 6248 1037 6250 1038
rect 6750 1037 6752 1038
rect 4474 1030 4476 1032
rect 5074 1030 5076 1032
rect 5674 1030 5676 1032
rect 4476 1028 4478 1030
rect 4482 1028 4484 1030
rect 4906 1028 4908 1030
rect 4932 1028 4934 1030
rect 5076 1028 5078 1030
rect 5082 1028 5084 1030
rect 5506 1028 5508 1030
rect 5532 1028 5534 1030
rect 5676 1028 5678 1030
rect 5682 1028 5684 1030
rect 6106 1028 6108 1030
rect 6132 1028 6134 1030
rect 4484 1026 4486 1028
rect 4904 1026 4906 1028
rect 4934 1026 4936 1028
rect 5084 1026 5086 1028
rect 5504 1026 5506 1028
rect 5534 1026 5536 1028
rect 5684 1026 5686 1028
rect 6104 1026 6106 1028
rect 6134 1026 6136 1028
rect 4484 1020 4486 1022
rect 4514 1020 4516 1022
rect 4544 1020 4546 1022
rect 4574 1020 4576 1022
rect 4604 1020 4606 1022
rect 4634 1020 4636 1022
rect 4664 1020 4666 1022
rect 4694 1020 4696 1022
rect 4724 1020 4726 1022
rect 4754 1020 4756 1022
rect 4784 1020 4786 1022
rect 4814 1020 4816 1022
rect 4844 1020 4846 1022
rect 4874 1020 4876 1022
rect 4904 1020 4906 1022
rect 4934 1020 4936 1022
rect 5084 1020 5086 1022
rect 5114 1020 5116 1022
rect 5144 1020 5146 1022
rect 5174 1020 5176 1022
rect 5204 1020 5206 1022
rect 5234 1020 5236 1022
rect 5264 1020 5266 1022
rect 5294 1020 5296 1022
rect 5324 1020 5326 1022
rect 5354 1020 5356 1022
rect 5384 1020 5386 1022
rect 5414 1020 5416 1022
rect 5444 1020 5446 1022
rect 5474 1020 5476 1022
rect 5504 1020 5506 1022
rect 5534 1020 5536 1022
rect 5684 1020 5686 1022
rect 5714 1020 5716 1022
rect 5744 1020 5746 1022
rect 5774 1020 5776 1022
rect 5804 1020 5806 1022
rect 5834 1020 5836 1022
rect 5864 1020 5866 1022
rect 5894 1020 5896 1022
rect 5924 1020 5926 1022
rect 5954 1020 5956 1022
rect 5984 1020 5986 1022
rect 6014 1020 6016 1022
rect 6044 1020 6046 1022
rect 6074 1020 6076 1022
rect 6104 1020 6106 1022
rect 6134 1020 6136 1022
rect 3250 1019 3252 1020
rect 3748 1019 3750 1020
rect 3850 1019 3852 1020
rect 4348 1019 4350 1020
rect 4476 1018 4478 1020
rect 4482 1018 4484 1020
rect 4506 1018 4508 1020
rect 4512 1018 4514 1020
rect 4536 1018 4538 1020
rect 4542 1018 4544 1020
rect 4566 1018 4568 1020
rect 4572 1018 4574 1020
rect 4596 1018 4598 1020
rect 4602 1018 4604 1020
rect 4626 1018 4628 1020
rect 4632 1018 4634 1020
rect 4656 1018 4658 1020
rect 4662 1018 4664 1020
rect 4686 1018 4688 1020
rect 4692 1018 4694 1020
rect 4716 1018 4718 1020
rect 4722 1018 4724 1020
rect 4746 1018 4748 1020
rect 4752 1018 4754 1020
rect 4776 1018 4778 1020
rect 4782 1018 4784 1020
rect 4806 1018 4808 1020
rect 4812 1018 4814 1020
rect 4836 1018 4838 1020
rect 4842 1018 4844 1020
rect 4866 1018 4868 1020
rect 4872 1018 4874 1020
rect 4896 1018 4898 1020
rect 4902 1018 4904 1020
rect 4926 1018 4928 1020
rect 4932 1018 4934 1020
rect 5076 1018 5078 1020
rect 5082 1018 5084 1020
rect 5106 1018 5108 1020
rect 5112 1018 5114 1020
rect 5136 1018 5138 1020
rect 5142 1018 5144 1020
rect 5166 1018 5168 1020
rect 5172 1018 5174 1020
rect 5196 1018 5198 1020
rect 5202 1018 5204 1020
rect 5226 1018 5228 1020
rect 5232 1018 5234 1020
rect 5256 1018 5258 1020
rect 5262 1018 5264 1020
rect 5286 1018 5288 1020
rect 5292 1018 5294 1020
rect 5316 1018 5318 1020
rect 5322 1018 5324 1020
rect 5346 1018 5348 1020
rect 5352 1018 5354 1020
rect 5376 1018 5378 1020
rect 5382 1018 5384 1020
rect 5406 1018 5408 1020
rect 5412 1018 5414 1020
rect 5436 1018 5438 1020
rect 5442 1018 5444 1020
rect 5466 1018 5468 1020
rect 5472 1018 5474 1020
rect 5496 1018 5498 1020
rect 5502 1018 5504 1020
rect 5526 1018 5528 1020
rect 5532 1018 5534 1020
rect 5676 1018 5678 1020
rect 5682 1018 5684 1020
rect 5706 1018 5708 1020
rect 5712 1018 5714 1020
rect 5736 1018 5738 1020
rect 5742 1018 5744 1020
rect 5766 1018 5768 1020
rect 5772 1018 5774 1020
rect 5796 1018 5798 1020
rect 5802 1018 5804 1020
rect 5826 1018 5828 1020
rect 5832 1018 5834 1020
rect 5856 1018 5858 1020
rect 5862 1018 5864 1020
rect 5886 1018 5888 1020
rect 5892 1018 5894 1020
rect 5916 1018 5918 1020
rect 5922 1018 5924 1020
rect 5946 1018 5948 1020
rect 5952 1018 5954 1020
rect 5976 1018 5978 1020
rect 5982 1018 5984 1020
rect 6006 1018 6008 1020
rect 6012 1018 6014 1020
rect 6036 1018 6038 1020
rect 6042 1018 6044 1020
rect 6066 1018 6068 1020
rect 6072 1018 6074 1020
rect 6096 1018 6098 1020
rect 6102 1018 6104 1020
rect 6126 1018 6128 1020
rect 6132 1018 6134 1020
rect 6250 1019 6252 1020
rect 6748 1019 6750 1020
rect 3248 1017 3250 1018
rect 3750 1017 3752 1018
rect 3848 1017 3850 1018
rect 4350 1017 4352 1018
rect 4474 1016 4476 1018
rect 4504 1016 4506 1018
rect 4534 1016 4536 1018
rect 4564 1016 4566 1018
rect 4594 1016 4596 1018
rect 4624 1016 4626 1018
rect 4654 1016 4656 1018
rect 4684 1016 4686 1018
rect 4714 1016 4716 1018
rect 4744 1016 4746 1018
rect 4774 1016 4776 1018
rect 4804 1016 4806 1018
rect 4834 1016 4836 1018
rect 4864 1016 4866 1018
rect 4894 1016 4896 1018
rect 4924 1016 4926 1018
rect 5074 1016 5076 1018
rect 5104 1016 5106 1018
rect 5134 1016 5136 1018
rect 5164 1016 5166 1018
rect 5194 1016 5196 1018
rect 5224 1016 5226 1018
rect 5254 1016 5256 1018
rect 5284 1016 5286 1018
rect 5314 1016 5316 1018
rect 5344 1016 5346 1018
rect 5374 1016 5376 1018
rect 5404 1016 5406 1018
rect 5434 1016 5436 1018
rect 5464 1016 5466 1018
rect 5494 1016 5496 1018
rect 5524 1016 5526 1018
rect 5674 1016 5676 1018
rect 5704 1016 5706 1018
rect 5734 1016 5736 1018
rect 5764 1016 5766 1018
rect 5794 1016 5796 1018
rect 5824 1016 5826 1018
rect 5854 1016 5856 1018
rect 5884 1016 5886 1018
rect 5914 1016 5916 1018
rect 5944 1016 5946 1018
rect 5974 1016 5976 1018
rect 6004 1016 6006 1018
rect 6034 1016 6036 1018
rect 6064 1016 6066 1018
rect 6094 1016 6096 1018
rect 6124 1016 6126 1018
rect 6248 1017 6250 1018
rect 6750 1017 6752 1018
rect 4474 1010 4476 1012
rect 4504 1010 4506 1012
rect 4534 1010 4536 1012
rect 4564 1010 4566 1012
rect 4594 1010 4596 1012
rect 4624 1010 4626 1012
rect 4654 1010 4656 1012
rect 4684 1010 4686 1012
rect 4714 1010 4716 1012
rect 4744 1010 4746 1012
rect 4774 1010 4776 1012
rect 4804 1010 4806 1012
rect 4834 1010 4836 1012
rect 4864 1010 4866 1012
rect 4894 1010 4896 1012
rect 4924 1010 4926 1012
rect 5074 1010 5076 1012
rect 5104 1010 5106 1012
rect 5134 1010 5136 1012
rect 5164 1010 5166 1012
rect 5194 1010 5196 1012
rect 5224 1010 5226 1012
rect 5254 1010 5256 1012
rect 5284 1010 5286 1012
rect 5314 1010 5316 1012
rect 5344 1010 5346 1012
rect 5374 1010 5376 1012
rect 5404 1010 5406 1012
rect 5434 1010 5436 1012
rect 5464 1010 5466 1012
rect 5494 1010 5496 1012
rect 5524 1010 5526 1012
rect 5674 1010 5676 1012
rect 5704 1010 5706 1012
rect 5734 1010 5736 1012
rect 5764 1010 5766 1012
rect 5794 1010 5796 1012
rect 5824 1010 5826 1012
rect 5854 1010 5856 1012
rect 5884 1010 5886 1012
rect 5914 1010 5916 1012
rect 5944 1010 5946 1012
rect 5974 1010 5976 1012
rect 6004 1010 6006 1012
rect 6034 1010 6036 1012
rect 6064 1010 6066 1012
rect 6094 1010 6096 1012
rect 6124 1010 6126 1012
rect 4476 1008 4478 1010
rect 4482 1008 4484 1010
rect 4506 1008 4508 1010
rect 4512 1008 4514 1010
rect 4536 1008 4538 1010
rect 4542 1008 4544 1010
rect 4566 1008 4568 1010
rect 4572 1008 4574 1010
rect 4596 1008 4598 1010
rect 4602 1008 4604 1010
rect 4626 1008 4628 1010
rect 4632 1008 4634 1010
rect 4656 1008 4658 1010
rect 4662 1008 4664 1010
rect 4686 1008 4688 1010
rect 4692 1008 4694 1010
rect 4716 1008 4718 1010
rect 4722 1008 4724 1010
rect 4746 1008 4748 1010
rect 4752 1008 4754 1010
rect 4776 1008 4778 1010
rect 4782 1008 4784 1010
rect 4806 1008 4808 1010
rect 4812 1008 4814 1010
rect 4836 1008 4838 1010
rect 4842 1008 4844 1010
rect 4866 1008 4868 1010
rect 4872 1008 4874 1010
rect 4896 1008 4898 1010
rect 4902 1008 4904 1010
rect 4926 1008 4928 1010
rect 4932 1008 4934 1010
rect 5076 1008 5078 1010
rect 5082 1008 5084 1010
rect 5106 1008 5108 1010
rect 5112 1008 5114 1010
rect 5136 1008 5138 1010
rect 5142 1008 5144 1010
rect 5166 1008 5168 1010
rect 5172 1008 5174 1010
rect 5196 1008 5198 1010
rect 5202 1008 5204 1010
rect 5226 1008 5228 1010
rect 5232 1008 5234 1010
rect 5256 1008 5258 1010
rect 5262 1008 5264 1010
rect 5286 1008 5288 1010
rect 5292 1008 5294 1010
rect 5316 1008 5318 1010
rect 5322 1008 5324 1010
rect 5346 1008 5348 1010
rect 5352 1008 5354 1010
rect 5376 1008 5378 1010
rect 5382 1008 5384 1010
rect 5406 1008 5408 1010
rect 5412 1008 5414 1010
rect 5436 1008 5438 1010
rect 5442 1008 5444 1010
rect 5466 1008 5468 1010
rect 5472 1008 5474 1010
rect 5496 1008 5498 1010
rect 5502 1008 5504 1010
rect 5526 1008 5528 1010
rect 5532 1008 5534 1010
rect 5676 1008 5678 1010
rect 5682 1008 5684 1010
rect 5706 1008 5708 1010
rect 5712 1008 5714 1010
rect 5736 1008 5738 1010
rect 5742 1008 5744 1010
rect 5766 1008 5768 1010
rect 5772 1008 5774 1010
rect 5796 1008 5798 1010
rect 5802 1008 5804 1010
rect 5826 1008 5828 1010
rect 5832 1008 5834 1010
rect 5856 1008 5858 1010
rect 5862 1008 5864 1010
rect 5886 1008 5888 1010
rect 5892 1008 5894 1010
rect 5916 1008 5918 1010
rect 5922 1008 5924 1010
rect 5946 1008 5948 1010
rect 5952 1008 5954 1010
rect 5976 1008 5978 1010
rect 5982 1008 5984 1010
rect 6006 1008 6008 1010
rect 6012 1008 6014 1010
rect 6036 1008 6038 1010
rect 6042 1008 6044 1010
rect 6066 1008 6068 1010
rect 6072 1008 6074 1010
rect 6096 1008 6098 1010
rect 6102 1008 6104 1010
rect 6126 1008 6128 1010
rect 6132 1008 6134 1010
rect 4484 1006 4486 1008
rect 4514 1006 4516 1008
rect 4544 1006 4546 1008
rect 4574 1006 4576 1008
rect 4604 1006 4606 1008
rect 4634 1006 4636 1008
rect 4664 1006 4666 1008
rect 4694 1006 4696 1008
rect 4724 1006 4726 1008
rect 4754 1006 4756 1008
rect 4784 1006 4786 1008
rect 4814 1006 4816 1008
rect 4844 1006 4846 1008
rect 4874 1006 4876 1008
rect 4904 1006 4906 1008
rect 4934 1006 4936 1008
rect 5084 1006 5086 1008
rect 5114 1006 5116 1008
rect 5144 1006 5146 1008
rect 5174 1006 5176 1008
rect 5204 1006 5206 1008
rect 5234 1006 5236 1008
rect 5264 1006 5266 1008
rect 5294 1006 5296 1008
rect 5324 1006 5326 1008
rect 5354 1006 5356 1008
rect 5384 1006 5386 1008
rect 5414 1006 5416 1008
rect 5444 1006 5446 1008
rect 5474 1006 5476 1008
rect 5504 1006 5506 1008
rect 5534 1006 5536 1008
rect 5684 1006 5686 1008
rect 5714 1006 5716 1008
rect 5744 1006 5746 1008
rect 5774 1006 5776 1008
rect 5804 1006 5806 1008
rect 5834 1006 5836 1008
rect 5864 1006 5866 1008
rect 5894 1006 5896 1008
rect 5924 1006 5926 1008
rect 5954 1006 5956 1008
rect 5984 1006 5986 1008
rect 6014 1006 6016 1008
rect 6044 1006 6046 1008
rect 6074 1006 6076 1008
rect 6104 1006 6106 1008
rect 6134 1006 6136 1008
rect 4484 1000 4486 1002
rect 4514 1000 4516 1002
rect 4544 1000 4546 1002
rect 4574 1000 4576 1002
rect 4604 1000 4606 1002
rect 4634 1000 4636 1002
rect 4664 1000 4666 1002
rect 4694 1000 4696 1002
rect 4724 1000 4726 1002
rect 4754 1000 4756 1002
rect 4784 1000 4786 1002
rect 4814 1000 4816 1002
rect 4844 1000 4846 1002
rect 4874 1000 4876 1002
rect 4904 1000 4906 1002
rect 4934 1000 4936 1002
rect 5084 1000 5086 1002
rect 5114 1000 5116 1002
rect 5144 1000 5146 1002
rect 5174 1000 5176 1002
rect 5204 1000 5206 1002
rect 5234 1000 5236 1002
rect 5264 1000 5266 1002
rect 5294 1000 5296 1002
rect 5324 1000 5326 1002
rect 5354 1000 5356 1002
rect 5384 1000 5386 1002
rect 5414 1000 5416 1002
rect 5444 1000 5446 1002
rect 5474 1000 5476 1002
rect 5504 1000 5506 1002
rect 5534 1000 5536 1002
rect 5684 1000 5686 1002
rect 5714 1000 5716 1002
rect 5744 1000 5746 1002
rect 5774 1000 5776 1002
rect 5804 1000 5806 1002
rect 5834 1000 5836 1002
rect 5864 1000 5866 1002
rect 5894 1000 5896 1002
rect 5924 1000 5926 1002
rect 5954 1000 5956 1002
rect 5984 1000 5986 1002
rect 6014 1000 6016 1002
rect 6044 1000 6046 1002
rect 6074 1000 6076 1002
rect 6104 1000 6106 1002
rect 6134 1000 6136 1002
rect 3250 999 3252 1000
rect 3748 999 3750 1000
rect 3850 999 3852 1000
rect 4348 999 4350 1000
rect 4476 998 4478 1000
rect 4482 998 4484 1000
rect 4506 998 4508 1000
rect 4512 998 4514 1000
rect 4536 998 4538 1000
rect 4542 998 4544 1000
rect 4566 998 4568 1000
rect 4572 998 4574 1000
rect 4596 998 4598 1000
rect 4602 998 4604 1000
rect 4626 998 4628 1000
rect 4632 998 4634 1000
rect 4656 998 4658 1000
rect 4662 998 4664 1000
rect 4686 998 4688 1000
rect 4692 998 4694 1000
rect 4716 998 4718 1000
rect 4722 998 4724 1000
rect 4746 998 4748 1000
rect 4752 998 4754 1000
rect 4776 998 4778 1000
rect 4782 998 4784 1000
rect 4806 998 4808 1000
rect 4812 998 4814 1000
rect 4836 998 4838 1000
rect 4842 998 4844 1000
rect 4866 998 4868 1000
rect 4872 998 4874 1000
rect 4896 998 4898 1000
rect 4902 998 4904 1000
rect 4926 998 4928 1000
rect 4932 998 4934 1000
rect 5076 998 5078 1000
rect 5082 998 5084 1000
rect 5106 998 5108 1000
rect 5112 998 5114 1000
rect 5136 998 5138 1000
rect 5142 998 5144 1000
rect 5166 998 5168 1000
rect 5172 998 5174 1000
rect 5196 998 5198 1000
rect 5202 998 5204 1000
rect 5226 998 5228 1000
rect 5232 998 5234 1000
rect 5256 998 5258 1000
rect 5262 998 5264 1000
rect 5286 998 5288 1000
rect 5292 998 5294 1000
rect 5316 998 5318 1000
rect 5322 998 5324 1000
rect 5346 998 5348 1000
rect 5352 998 5354 1000
rect 5376 998 5378 1000
rect 5382 998 5384 1000
rect 5406 998 5408 1000
rect 5412 998 5414 1000
rect 5436 998 5438 1000
rect 5442 998 5444 1000
rect 5466 998 5468 1000
rect 5472 998 5474 1000
rect 5496 998 5498 1000
rect 5502 998 5504 1000
rect 5526 998 5528 1000
rect 5532 998 5534 1000
rect 5676 998 5678 1000
rect 5682 998 5684 1000
rect 5706 998 5708 1000
rect 5712 998 5714 1000
rect 5736 998 5738 1000
rect 5742 998 5744 1000
rect 5766 998 5768 1000
rect 5772 998 5774 1000
rect 5796 998 5798 1000
rect 5802 998 5804 1000
rect 5826 998 5828 1000
rect 5832 998 5834 1000
rect 5856 998 5858 1000
rect 5862 998 5864 1000
rect 5886 998 5888 1000
rect 5892 998 5894 1000
rect 5916 998 5918 1000
rect 5922 998 5924 1000
rect 5946 998 5948 1000
rect 5952 998 5954 1000
rect 5976 998 5978 1000
rect 5982 998 5984 1000
rect 6006 998 6008 1000
rect 6012 998 6014 1000
rect 6036 998 6038 1000
rect 6042 998 6044 1000
rect 6066 998 6068 1000
rect 6072 998 6074 1000
rect 6096 998 6098 1000
rect 6102 998 6104 1000
rect 6126 998 6128 1000
rect 6132 998 6134 1000
rect 6250 999 6252 1000
rect 6748 999 6750 1000
rect 3248 997 3250 998
rect 3750 997 3752 998
rect 3848 997 3850 998
rect 4350 997 4352 998
rect 4474 996 4476 998
rect 4504 996 4506 998
rect 4534 996 4536 998
rect 4564 996 4566 998
rect 4594 996 4596 998
rect 4624 996 4626 998
rect 4654 996 4656 998
rect 4684 996 4686 998
rect 4714 996 4716 998
rect 4744 996 4746 998
rect 4774 996 4776 998
rect 4804 996 4806 998
rect 4834 996 4836 998
rect 4864 996 4866 998
rect 4894 996 4896 998
rect 4924 996 4926 998
rect 5074 996 5076 998
rect 5104 996 5106 998
rect 5134 996 5136 998
rect 5164 996 5166 998
rect 5194 996 5196 998
rect 5224 996 5226 998
rect 5254 996 5256 998
rect 5284 996 5286 998
rect 5314 996 5316 998
rect 5344 996 5346 998
rect 5374 996 5376 998
rect 5404 996 5406 998
rect 5434 996 5436 998
rect 5464 996 5466 998
rect 5494 996 5496 998
rect 5524 996 5526 998
rect 5674 996 5676 998
rect 5704 996 5706 998
rect 5734 996 5736 998
rect 5764 996 5766 998
rect 5794 996 5796 998
rect 5824 996 5826 998
rect 5854 996 5856 998
rect 5884 996 5886 998
rect 5914 996 5916 998
rect 5944 996 5946 998
rect 5974 996 5976 998
rect 6004 996 6006 998
rect 6034 996 6036 998
rect 6064 996 6066 998
rect 6094 996 6096 998
rect 6124 996 6126 998
rect 6248 997 6250 998
rect 6750 997 6752 998
rect 4474 990 4476 992
rect 4504 990 4506 992
rect 4534 990 4536 992
rect 4564 990 4566 992
rect 4594 990 4596 992
rect 4624 990 4626 992
rect 4654 990 4656 992
rect 4684 990 4686 992
rect 4714 990 4716 992
rect 4744 990 4746 992
rect 4774 990 4776 992
rect 4804 990 4806 992
rect 4834 990 4836 992
rect 4864 990 4866 992
rect 4894 990 4896 992
rect 4924 990 4926 992
rect 5074 990 5076 992
rect 5104 990 5106 992
rect 5134 990 5136 992
rect 5164 990 5166 992
rect 5194 990 5196 992
rect 5224 990 5226 992
rect 5254 990 5256 992
rect 5284 990 5286 992
rect 5314 990 5316 992
rect 5344 990 5346 992
rect 5374 990 5376 992
rect 5404 990 5406 992
rect 5434 990 5436 992
rect 5464 990 5466 992
rect 5494 990 5496 992
rect 5524 990 5526 992
rect 5674 990 5676 992
rect 5704 990 5706 992
rect 5734 990 5736 992
rect 5764 990 5766 992
rect 5794 990 5796 992
rect 5824 990 5826 992
rect 5854 990 5856 992
rect 5884 990 5886 992
rect 5914 990 5916 992
rect 5944 990 5946 992
rect 5974 990 5976 992
rect 6004 990 6006 992
rect 6034 990 6036 992
rect 6064 990 6066 992
rect 6094 990 6096 992
rect 6124 990 6126 992
rect 4476 988 4478 990
rect 4482 988 4484 990
rect 4506 988 4508 990
rect 4512 988 4514 990
rect 4536 988 4538 990
rect 4542 988 4544 990
rect 4566 988 4568 990
rect 4572 988 4574 990
rect 4596 988 4598 990
rect 4602 988 4604 990
rect 4626 988 4628 990
rect 4632 988 4634 990
rect 4656 988 4658 990
rect 4662 988 4664 990
rect 4686 988 4688 990
rect 4692 988 4694 990
rect 4716 988 4718 990
rect 4722 988 4724 990
rect 4746 988 4748 990
rect 4752 988 4754 990
rect 4776 988 4778 990
rect 4782 988 4784 990
rect 4806 988 4808 990
rect 4812 988 4814 990
rect 4836 988 4838 990
rect 4842 988 4844 990
rect 4866 988 4868 990
rect 4872 988 4874 990
rect 4896 988 4898 990
rect 4902 988 4904 990
rect 4926 988 4928 990
rect 4932 988 4934 990
rect 5076 988 5078 990
rect 5082 988 5084 990
rect 5106 988 5108 990
rect 5112 988 5114 990
rect 5136 988 5138 990
rect 5142 988 5144 990
rect 5166 988 5168 990
rect 5172 988 5174 990
rect 5196 988 5198 990
rect 5202 988 5204 990
rect 5226 988 5228 990
rect 5232 988 5234 990
rect 5256 988 5258 990
rect 5262 988 5264 990
rect 5286 988 5288 990
rect 5292 988 5294 990
rect 5316 988 5318 990
rect 5322 988 5324 990
rect 5346 988 5348 990
rect 5352 988 5354 990
rect 5376 988 5378 990
rect 5382 988 5384 990
rect 5406 988 5408 990
rect 5412 988 5414 990
rect 5436 988 5438 990
rect 5442 988 5444 990
rect 5466 988 5468 990
rect 5472 988 5474 990
rect 5496 988 5498 990
rect 5502 988 5504 990
rect 5526 988 5528 990
rect 5532 988 5534 990
rect 5676 988 5678 990
rect 5682 988 5684 990
rect 5706 988 5708 990
rect 5712 988 5714 990
rect 5736 988 5738 990
rect 5742 988 5744 990
rect 5766 988 5768 990
rect 5772 988 5774 990
rect 5796 988 5798 990
rect 5802 988 5804 990
rect 5826 988 5828 990
rect 5832 988 5834 990
rect 5856 988 5858 990
rect 5862 988 5864 990
rect 5886 988 5888 990
rect 5892 988 5894 990
rect 5916 988 5918 990
rect 5922 988 5924 990
rect 5946 988 5948 990
rect 5952 988 5954 990
rect 5976 988 5978 990
rect 5982 988 5984 990
rect 6006 988 6008 990
rect 6012 988 6014 990
rect 6036 988 6038 990
rect 6042 988 6044 990
rect 6066 988 6068 990
rect 6072 988 6074 990
rect 6096 988 6098 990
rect 6102 988 6104 990
rect 6126 988 6128 990
rect 6132 988 6134 990
rect 4484 986 4486 988
rect 4514 986 4516 988
rect 4544 986 4546 988
rect 4574 986 4576 988
rect 4604 986 4606 988
rect 4634 986 4636 988
rect 4664 986 4666 988
rect 4694 986 4696 988
rect 4724 986 4726 988
rect 4754 986 4756 988
rect 4784 986 4786 988
rect 4814 986 4816 988
rect 4844 986 4846 988
rect 4874 986 4876 988
rect 4904 986 4906 988
rect 4934 986 4936 988
rect 5084 986 5086 988
rect 5114 986 5116 988
rect 5144 986 5146 988
rect 5174 986 5176 988
rect 5204 986 5206 988
rect 5234 986 5236 988
rect 5264 986 5266 988
rect 5294 986 5296 988
rect 5324 986 5326 988
rect 5354 986 5356 988
rect 5384 986 5386 988
rect 5414 986 5416 988
rect 5444 986 5446 988
rect 5474 986 5476 988
rect 5504 986 5506 988
rect 5534 986 5536 988
rect 5684 986 5686 988
rect 5714 986 5716 988
rect 5744 986 5746 988
rect 5774 986 5776 988
rect 5804 986 5806 988
rect 5834 986 5836 988
rect 5864 986 5866 988
rect 5894 986 5896 988
rect 5924 986 5926 988
rect 5954 986 5956 988
rect 5984 986 5986 988
rect 6014 986 6016 988
rect 6044 986 6046 988
rect 6074 986 6076 988
rect 6104 986 6106 988
rect 6134 986 6136 988
rect 3296 984 3298 986
rect 3702 984 3704 986
rect 3896 984 3898 986
rect 4302 984 4304 986
rect 6296 984 6298 986
rect 6702 984 6704 986
rect 3294 982 3296 984
rect 3704 982 3706 984
rect 3894 982 3896 984
rect 4304 982 4306 984
rect 6294 982 6296 984
rect 6704 982 6706 984
rect 4484 980 4486 982
rect 4514 980 4516 982
rect 4544 980 4546 982
rect 4574 980 4576 982
rect 4604 980 4606 982
rect 4634 980 4636 982
rect 4664 980 4666 982
rect 4694 980 4696 982
rect 4724 980 4726 982
rect 4754 980 4756 982
rect 4784 980 4786 982
rect 4814 980 4816 982
rect 4844 980 4846 982
rect 4874 980 4876 982
rect 4904 980 4906 982
rect 4934 980 4936 982
rect 5084 980 5086 982
rect 5114 980 5116 982
rect 5144 980 5146 982
rect 5174 980 5176 982
rect 5204 980 5206 982
rect 5234 980 5236 982
rect 5264 980 5266 982
rect 5294 980 5296 982
rect 5324 980 5326 982
rect 5354 980 5356 982
rect 5384 980 5386 982
rect 5414 980 5416 982
rect 5444 980 5446 982
rect 5474 980 5476 982
rect 5504 980 5506 982
rect 5534 980 5536 982
rect 5684 980 5686 982
rect 5714 980 5716 982
rect 5744 980 5746 982
rect 5774 980 5776 982
rect 5804 980 5806 982
rect 5834 980 5836 982
rect 5864 980 5866 982
rect 5894 980 5896 982
rect 5924 980 5926 982
rect 5954 980 5956 982
rect 5984 980 5986 982
rect 6014 980 6016 982
rect 6044 980 6046 982
rect 6074 980 6076 982
rect 6104 980 6106 982
rect 6134 980 6136 982
rect 3250 979 3252 980
rect 3748 979 3750 980
rect 3850 979 3852 980
rect 4348 979 4350 980
rect 4476 978 4478 980
rect 4482 978 4484 980
rect 4506 978 4508 980
rect 4512 978 4514 980
rect 4536 978 4538 980
rect 4542 978 4544 980
rect 4566 978 4568 980
rect 4572 978 4574 980
rect 4596 978 4598 980
rect 4602 978 4604 980
rect 4626 978 4628 980
rect 4632 978 4634 980
rect 4656 978 4658 980
rect 4662 978 4664 980
rect 4686 978 4688 980
rect 4692 978 4694 980
rect 4716 978 4718 980
rect 4722 978 4724 980
rect 4746 978 4748 980
rect 4752 978 4754 980
rect 4776 978 4778 980
rect 4782 978 4784 980
rect 4806 978 4808 980
rect 4812 978 4814 980
rect 4836 978 4838 980
rect 4842 978 4844 980
rect 4866 978 4868 980
rect 4872 978 4874 980
rect 4896 978 4898 980
rect 4902 978 4904 980
rect 4926 978 4928 980
rect 4932 978 4934 980
rect 5076 978 5078 980
rect 5082 978 5084 980
rect 5106 978 5108 980
rect 5112 978 5114 980
rect 5136 978 5138 980
rect 5142 978 5144 980
rect 5166 978 5168 980
rect 5172 978 5174 980
rect 5196 978 5198 980
rect 5202 978 5204 980
rect 5226 978 5228 980
rect 5232 978 5234 980
rect 5256 978 5258 980
rect 5262 978 5264 980
rect 5286 978 5288 980
rect 5292 978 5294 980
rect 5316 978 5318 980
rect 5322 978 5324 980
rect 5346 978 5348 980
rect 5352 978 5354 980
rect 5376 978 5378 980
rect 5382 978 5384 980
rect 5406 978 5408 980
rect 5412 978 5414 980
rect 5436 978 5438 980
rect 5442 978 5444 980
rect 5466 978 5468 980
rect 5472 978 5474 980
rect 5496 978 5498 980
rect 5502 978 5504 980
rect 5526 978 5528 980
rect 5532 978 5534 980
rect 5676 978 5678 980
rect 5682 978 5684 980
rect 5706 978 5708 980
rect 5712 978 5714 980
rect 5736 978 5738 980
rect 5742 978 5744 980
rect 5766 978 5768 980
rect 5772 978 5774 980
rect 5796 978 5798 980
rect 5802 978 5804 980
rect 5826 978 5828 980
rect 5832 978 5834 980
rect 5856 978 5858 980
rect 5862 978 5864 980
rect 5886 978 5888 980
rect 5892 978 5894 980
rect 5916 978 5918 980
rect 5922 978 5924 980
rect 5946 978 5948 980
rect 5952 978 5954 980
rect 5976 978 5978 980
rect 5982 978 5984 980
rect 6006 978 6008 980
rect 6012 978 6014 980
rect 6036 978 6038 980
rect 6042 978 6044 980
rect 6066 978 6068 980
rect 6072 978 6074 980
rect 6096 978 6098 980
rect 6102 978 6104 980
rect 6126 978 6128 980
rect 6132 978 6134 980
rect 6250 979 6252 980
rect 6748 979 6750 980
rect 3248 977 3250 978
rect 3750 977 3752 978
rect 3848 977 3850 978
rect 4350 977 4352 978
rect 4474 976 4476 978
rect 4504 976 4506 978
rect 4534 976 4536 978
rect 4564 976 4566 978
rect 4594 976 4596 978
rect 4624 976 4626 978
rect 4654 976 4656 978
rect 4684 976 4686 978
rect 4714 976 4716 978
rect 4744 976 4746 978
rect 4774 976 4776 978
rect 4804 976 4806 978
rect 4834 976 4836 978
rect 4864 976 4866 978
rect 4894 976 4896 978
rect 4924 976 4926 978
rect 5074 976 5076 978
rect 5104 976 5106 978
rect 5134 976 5136 978
rect 5164 976 5166 978
rect 5194 976 5196 978
rect 5224 976 5226 978
rect 5254 976 5256 978
rect 5284 976 5286 978
rect 5314 976 5316 978
rect 5344 976 5346 978
rect 5374 976 5376 978
rect 5404 976 5406 978
rect 5434 976 5436 978
rect 5464 976 5466 978
rect 5494 976 5496 978
rect 5524 976 5526 978
rect 5674 976 5676 978
rect 5704 976 5706 978
rect 5734 976 5736 978
rect 5764 976 5766 978
rect 5794 976 5796 978
rect 5824 976 5826 978
rect 5854 976 5856 978
rect 5884 976 5886 978
rect 5914 976 5916 978
rect 5944 976 5946 978
rect 5974 976 5976 978
rect 6004 976 6006 978
rect 6034 976 6036 978
rect 6064 976 6066 978
rect 6094 976 6096 978
rect 6124 976 6126 978
rect 6248 977 6250 978
rect 6750 977 6752 978
rect 3250 959 3252 960
rect 3748 959 3750 960
rect 3850 959 3852 960
rect 4348 959 4350 960
rect 6250 959 6252 960
rect 6748 959 6750 960
rect 3248 957 3250 958
rect 3750 957 3752 958
rect 3848 957 3850 958
rect 4350 957 4352 958
rect 6248 957 6250 958
rect 6750 957 6752 958
rect 4474 950 4476 952
rect 4504 950 4506 952
rect 4534 950 4536 952
rect 4564 950 4566 952
rect 4594 950 4596 952
rect 4624 950 4626 952
rect 4654 950 4656 952
rect 4684 950 4686 952
rect 4714 950 4716 952
rect 4744 950 4746 952
rect 4774 950 4776 952
rect 4804 950 4806 952
rect 4834 950 4836 952
rect 4864 950 4866 952
rect 4894 950 4896 952
rect 4924 950 4926 952
rect 5074 950 5076 952
rect 5104 950 5106 952
rect 5134 950 5136 952
rect 5164 950 5166 952
rect 5194 950 5196 952
rect 5224 950 5226 952
rect 5254 950 5256 952
rect 5284 950 5286 952
rect 5314 950 5316 952
rect 5344 950 5346 952
rect 5374 950 5376 952
rect 5404 950 5406 952
rect 5434 950 5436 952
rect 5464 950 5466 952
rect 5494 950 5496 952
rect 5524 950 5526 952
rect 5674 950 5676 952
rect 5704 950 5706 952
rect 5734 950 5736 952
rect 5764 950 5766 952
rect 5794 950 5796 952
rect 5824 950 5826 952
rect 5854 950 5856 952
rect 5884 950 5886 952
rect 5914 950 5916 952
rect 5944 950 5946 952
rect 5974 950 5976 952
rect 6004 950 6006 952
rect 6034 950 6036 952
rect 6064 950 6066 952
rect 6094 950 6096 952
rect 6124 950 6126 952
rect 4476 948 4478 950
rect 4482 948 4484 950
rect 4506 948 4508 950
rect 4512 948 4514 950
rect 4536 948 4538 950
rect 4542 948 4544 950
rect 4566 948 4568 950
rect 4572 948 4574 950
rect 4596 948 4598 950
rect 4602 948 4604 950
rect 4626 948 4628 950
rect 4632 948 4634 950
rect 4656 948 4658 950
rect 4662 948 4664 950
rect 4686 948 4688 950
rect 4692 948 4694 950
rect 4716 948 4718 950
rect 4722 948 4724 950
rect 4746 948 4748 950
rect 4752 948 4754 950
rect 4776 948 4778 950
rect 4782 948 4784 950
rect 4806 948 4808 950
rect 4812 948 4814 950
rect 4836 948 4838 950
rect 4842 948 4844 950
rect 4866 948 4868 950
rect 4872 948 4874 950
rect 4896 948 4898 950
rect 4902 948 4904 950
rect 4926 948 4928 950
rect 4932 948 4934 950
rect 5076 948 5078 950
rect 5082 948 5084 950
rect 5106 948 5108 950
rect 5112 948 5114 950
rect 5136 948 5138 950
rect 5142 948 5144 950
rect 5166 948 5168 950
rect 5172 948 5174 950
rect 5196 948 5198 950
rect 5202 948 5204 950
rect 5226 948 5228 950
rect 5232 948 5234 950
rect 5256 948 5258 950
rect 5262 948 5264 950
rect 5286 948 5288 950
rect 5292 948 5294 950
rect 5316 948 5318 950
rect 5322 948 5324 950
rect 5346 948 5348 950
rect 5352 948 5354 950
rect 5376 948 5378 950
rect 5382 948 5384 950
rect 5406 948 5408 950
rect 5412 948 5414 950
rect 5436 948 5438 950
rect 5442 948 5444 950
rect 5466 948 5468 950
rect 5472 948 5474 950
rect 5496 948 5498 950
rect 5502 948 5504 950
rect 5526 948 5528 950
rect 5532 948 5534 950
rect 5676 948 5678 950
rect 5682 948 5684 950
rect 5706 948 5708 950
rect 5712 948 5714 950
rect 5736 948 5738 950
rect 5742 948 5744 950
rect 5766 948 5768 950
rect 5772 948 5774 950
rect 5796 948 5798 950
rect 5802 948 5804 950
rect 5826 948 5828 950
rect 5832 948 5834 950
rect 5856 948 5858 950
rect 5862 948 5864 950
rect 5886 948 5888 950
rect 5892 948 5894 950
rect 5916 948 5918 950
rect 5922 948 5924 950
rect 5946 948 5948 950
rect 5952 948 5954 950
rect 5976 948 5978 950
rect 5982 948 5984 950
rect 6006 948 6008 950
rect 6012 948 6014 950
rect 6036 948 6038 950
rect 6042 948 6044 950
rect 6066 948 6068 950
rect 6072 948 6074 950
rect 6096 948 6098 950
rect 6102 948 6104 950
rect 6126 948 6128 950
rect 6132 948 6134 950
rect 4484 946 4486 948
rect 4514 946 4516 948
rect 4544 946 4546 948
rect 4574 946 4576 948
rect 4604 946 4606 948
rect 4634 946 4636 948
rect 4664 946 4666 948
rect 4694 946 4696 948
rect 4724 946 4726 948
rect 4754 946 4756 948
rect 4784 946 4786 948
rect 4814 946 4816 948
rect 4844 946 4846 948
rect 4874 946 4876 948
rect 4904 946 4906 948
rect 4934 946 4936 948
rect 5084 946 5086 948
rect 5114 946 5116 948
rect 5144 946 5146 948
rect 5174 946 5176 948
rect 5204 946 5206 948
rect 5234 946 5236 948
rect 5264 946 5266 948
rect 5294 946 5296 948
rect 5324 946 5326 948
rect 5354 946 5356 948
rect 5384 946 5386 948
rect 5414 946 5416 948
rect 5444 946 5446 948
rect 5474 946 5476 948
rect 5504 946 5506 948
rect 5534 946 5536 948
rect 5684 946 5686 948
rect 5714 946 5716 948
rect 5744 946 5746 948
rect 5774 946 5776 948
rect 5804 946 5806 948
rect 5834 946 5836 948
rect 5864 946 5866 948
rect 5894 946 5896 948
rect 5924 946 5926 948
rect 5954 946 5956 948
rect 5984 946 5986 948
rect 6014 946 6016 948
rect 6044 946 6046 948
rect 6074 946 6076 948
rect 6104 946 6106 948
rect 6134 946 6136 948
rect 4484 940 4486 942
rect 4514 940 4516 942
rect 4544 940 4546 942
rect 4574 940 4576 942
rect 4604 940 4606 942
rect 4634 940 4636 942
rect 4664 940 4666 942
rect 4694 940 4696 942
rect 4724 940 4726 942
rect 4754 940 4756 942
rect 4784 940 4786 942
rect 4814 940 4816 942
rect 4844 940 4846 942
rect 4874 940 4876 942
rect 4904 940 4906 942
rect 4934 940 4936 942
rect 5084 940 5086 942
rect 5114 940 5116 942
rect 5144 940 5146 942
rect 5174 940 5176 942
rect 5204 940 5206 942
rect 5234 940 5236 942
rect 5264 940 5266 942
rect 5294 940 5296 942
rect 5324 940 5326 942
rect 5354 940 5356 942
rect 5384 940 5386 942
rect 5414 940 5416 942
rect 5444 940 5446 942
rect 5474 940 5476 942
rect 5504 940 5506 942
rect 5534 940 5536 942
rect 5684 940 5686 942
rect 5714 940 5716 942
rect 5744 940 5746 942
rect 5774 940 5776 942
rect 5804 940 5806 942
rect 5834 940 5836 942
rect 5864 940 5866 942
rect 5894 940 5896 942
rect 5924 940 5926 942
rect 5954 940 5956 942
rect 5984 940 5986 942
rect 6014 940 6016 942
rect 6044 940 6046 942
rect 6074 940 6076 942
rect 6104 940 6106 942
rect 6134 940 6136 942
rect 3250 939 3252 940
rect 3748 939 3750 940
rect 3850 939 3852 940
rect 4348 939 4350 940
rect 4476 938 4478 940
rect 4482 938 4484 940
rect 4506 938 4508 940
rect 4512 938 4514 940
rect 4536 938 4538 940
rect 4542 938 4544 940
rect 4566 938 4568 940
rect 4572 938 4574 940
rect 4596 938 4598 940
rect 4602 938 4604 940
rect 4626 938 4628 940
rect 4632 938 4634 940
rect 4656 938 4658 940
rect 4662 938 4664 940
rect 4686 938 4688 940
rect 4692 938 4694 940
rect 4716 938 4718 940
rect 4722 938 4724 940
rect 4746 938 4748 940
rect 4752 938 4754 940
rect 4776 938 4778 940
rect 4782 938 4784 940
rect 4806 938 4808 940
rect 4812 938 4814 940
rect 4836 938 4838 940
rect 4842 938 4844 940
rect 4866 938 4868 940
rect 4872 938 4874 940
rect 4896 938 4898 940
rect 4902 938 4904 940
rect 4926 938 4928 940
rect 4932 938 4934 940
rect 5076 938 5078 940
rect 5082 938 5084 940
rect 5106 938 5108 940
rect 5112 938 5114 940
rect 5136 938 5138 940
rect 5142 938 5144 940
rect 5166 938 5168 940
rect 5172 938 5174 940
rect 5196 938 5198 940
rect 5202 938 5204 940
rect 5226 938 5228 940
rect 5232 938 5234 940
rect 5256 938 5258 940
rect 5262 938 5264 940
rect 5286 938 5288 940
rect 5292 938 5294 940
rect 5316 938 5318 940
rect 5322 938 5324 940
rect 5346 938 5348 940
rect 5352 938 5354 940
rect 5376 938 5378 940
rect 5382 938 5384 940
rect 5406 938 5408 940
rect 5412 938 5414 940
rect 5436 938 5438 940
rect 5442 938 5444 940
rect 5466 938 5468 940
rect 5472 938 5474 940
rect 5496 938 5498 940
rect 5502 938 5504 940
rect 5526 938 5528 940
rect 5532 938 5534 940
rect 5676 938 5678 940
rect 5682 938 5684 940
rect 5706 938 5708 940
rect 5712 938 5714 940
rect 5736 938 5738 940
rect 5742 938 5744 940
rect 5766 938 5768 940
rect 5772 938 5774 940
rect 5796 938 5798 940
rect 5802 938 5804 940
rect 5826 938 5828 940
rect 5832 938 5834 940
rect 5856 938 5858 940
rect 5862 938 5864 940
rect 5886 938 5888 940
rect 5892 938 5894 940
rect 5916 938 5918 940
rect 5922 938 5924 940
rect 5946 938 5948 940
rect 5952 938 5954 940
rect 5976 938 5978 940
rect 5982 938 5984 940
rect 6006 938 6008 940
rect 6012 938 6014 940
rect 6036 938 6038 940
rect 6042 938 6044 940
rect 6066 938 6068 940
rect 6072 938 6074 940
rect 6096 938 6098 940
rect 6102 938 6104 940
rect 6126 938 6128 940
rect 6132 938 6134 940
rect 6250 939 6252 940
rect 6748 939 6750 940
rect 3248 937 3250 938
rect 3750 937 3752 938
rect 3848 937 3850 938
rect 4350 937 4352 938
rect 4474 936 4476 938
rect 4504 936 4506 938
rect 4534 936 4536 938
rect 4564 936 4566 938
rect 4594 936 4596 938
rect 4624 936 4626 938
rect 4654 936 4656 938
rect 4684 936 4686 938
rect 4714 936 4716 938
rect 4744 936 4746 938
rect 4774 936 4776 938
rect 4804 936 4806 938
rect 4834 936 4836 938
rect 4864 936 4866 938
rect 4894 936 4896 938
rect 4924 936 4926 938
rect 5074 936 5076 938
rect 5104 936 5106 938
rect 5134 936 5136 938
rect 5164 936 5166 938
rect 5194 936 5196 938
rect 5224 936 5226 938
rect 5254 936 5256 938
rect 5284 936 5286 938
rect 5314 936 5316 938
rect 5344 936 5346 938
rect 5374 936 5376 938
rect 5404 936 5406 938
rect 5434 936 5436 938
rect 5464 936 5466 938
rect 5494 936 5496 938
rect 5524 936 5526 938
rect 5674 936 5676 938
rect 5704 936 5706 938
rect 5734 936 5736 938
rect 5764 936 5766 938
rect 5794 936 5796 938
rect 5824 936 5826 938
rect 5854 936 5856 938
rect 5884 936 5886 938
rect 5914 936 5916 938
rect 5944 936 5946 938
rect 5974 936 5976 938
rect 6004 936 6006 938
rect 6034 936 6036 938
rect 6064 936 6066 938
rect 6094 936 6096 938
rect 6124 936 6126 938
rect 6248 937 6250 938
rect 6750 937 6752 938
rect 4474 930 4476 932
rect 4504 930 4506 932
rect 4534 930 4536 932
rect 4564 930 4566 932
rect 4594 930 4596 932
rect 4624 930 4626 932
rect 4654 930 4656 932
rect 4684 930 4686 932
rect 4714 930 4716 932
rect 4744 930 4746 932
rect 4774 930 4776 932
rect 4804 930 4806 932
rect 4834 930 4836 932
rect 4864 930 4866 932
rect 4894 930 4896 932
rect 4924 930 4926 932
rect 5074 930 5076 932
rect 5104 930 5106 932
rect 5134 930 5136 932
rect 5164 930 5166 932
rect 5194 930 5196 932
rect 5224 930 5226 932
rect 5254 930 5256 932
rect 5284 930 5286 932
rect 5314 930 5316 932
rect 5344 930 5346 932
rect 5374 930 5376 932
rect 5404 930 5406 932
rect 5434 930 5436 932
rect 5464 930 5466 932
rect 5494 930 5496 932
rect 5524 930 5526 932
rect 5674 930 5676 932
rect 5704 930 5706 932
rect 5734 930 5736 932
rect 5764 930 5766 932
rect 5794 930 5796 932
rect 5824 930 5826 932
rect 5854 930 5856 932
rect 5884 930 5886 932
rect 5914 930 5916 932
rect 5944 930 5946 932
rect 5974 930 5976 932
rect 6004 930 6006 932
rect 6034 930 6036 932
rect 6064 930 6066 932
rect 6094 930 6096 932
rect 6124 930 6126 932
rect 4476 928 4478 930
rect 4482 928 4484 930
rect 4506 928 4508 930
rect 4512 928 4514 930
rect 4536 928 4538 930
rect 4542 928 4544 930
rect 4566 928 4568 930
rect 4572 928 4574 930
rect 4596 928 4598 930
rect 4602 928 4604 930
rect 4626 928 4628 930
rect 4632 928 4634 930
rect 4656 928 4658 930
rect 4662 928 4664 930
rect 4686 928 4688 930
rect 4692 928 4694 930
rect 4716 928 4718 930
rect 4722 928 4724 930
rect 4746 928 4748 930
rect 4752 928 4754 930
rect 4776 928 4778 930
rect 4782 928 4784 930
rect 4806 928 4808 930
rect 4812 928 4814 930
rect 4836 928 4838 930
rect 4842 928 4844 930
rect 4866 928 4868 930
rect 4872 928 4874 930
rect 4896 928 4898 930
rect 4902 928 4904 930
rect 4926 928 4928 930
rect 4932 928 4934 930
rect 5076 928 5078 930
rect 5082 928 5084 930
rect 5106 928 5108 930
rect 5112 928 5114 930
rect 5136 928 5138 930
rect 5142 928 5144 930
rect 5166 928 5168 930
rect 5172 928 5174 930
rect 5196 928 5198 930
rect 5202 928 5204 930
rect 5226 928 5228 930
rect 5232 928 5234 930
rect 5256 928 5258 930
rect 5262 928 5264 930
rect 5286 928 5288 930
rect 5292 928 5294 930
rect 5316 928 5318 930
rect 5322 928 5324 930
rect 5346 928 5348 930
rect 5352 928 5354 930
rect 5376 928 5378 930
rect 5382 928 5384 930
rect 5406 928 5408 930
rect 5412 928 5414 930
rect 5436 928 5438 930
rect 5442 928 5444 930
rect 5466 928 5468 930
rect 5472 928 5474 930
rect 5496 928 5498 930
rect 5502 928 5504 930
rect 5526 928 5528 930
rect 5532 928 5534 930
rect 5676 928 5678 930
rect 5682 928 5684 930
rect 5706 928 5708 930
rect 5712 928 5714 930
rect 5736 928 5738 930
rect 5742 928 5744 930
rect 5766 928 5768 930
rect 5772 928 5774 930
rect 5796 928 5798 930
rect 5802 928 5804 930
rect 5826 928 5828 930
rect 5832 928 5834 930
rect 5856 928 5858 930
rect 5862 928 5864 930
rect 5886 928 5888 930
rect 5892 928 5894 930
rect 5916 928 5918 930
rect 5922 928 5924 930
rect 5946 928 5948 930
rect 5952 928 5954 930
rect 5976 928 5978 930
rect 5982 928 5984 930
rect 6006 928 6008 930
rect 6012 928 6014 930
rect 6036 928 6038 930
rect 6042 928 6044 930
rect 6066 928 6068 930
rect 6072 928 6074 930
rect 6096 928 6098 930
rect 6102 928 6104 930
rect 6126 928 6128 930
rect 6132 928 6134 930
rect 4484 926 4486 928
rect 4514 926 4516 928
rect 4544 926 4546 928
rect 4574 926 4576 928
rect 4604 926 4606 928
rect 4634 926 4636 928
rect 4664 926 4666 928
rect 4694 926 4696 928
rect 4724 926 4726 928
rect 4754 926 4756 928
rect 4784 926 4786 928
rect 4814 926 4816 928
rect 4844 926 4846 928
rect 4874 926 4876 928
rect 4904 926 4906 928
rect 4934 926 4936 928
rect 5084 926 5086 928
rect 5114 926 5116 928
rect 5144 926 5146 928
rect 5174 926 5176 928
rect 5204 926 5206 928
rect 5234 926 5236 928
rect 5264 926 5266 928
rect 5294 926 5296 928
rect 5324 926 5326 928
rect 5354 926 5356 928
rect 5384 926 5386 928
rect 5414 926 5416 928
rect 5444 926 5446 928
rect 5474 926 5476 928
rect 5504 926 5506 928
rect 5534 926 5536 928
rect 5684 926 5686 928
rect 5714 926 5716 928
rect 5744 926 5746 928
rect 5774 926 5776 928
rect 5804 926 5806 928
rect 5834 926 5836 928
rect 5864 926 5866 928
rect 5894 926 5896 928
rect 5924 926 5926 928
rect 5954 926 5956 928
rect 5984 926 5986 928
rect 6014 926 6016 928
rect 6044 926 6046 928
rect 6074 926 6076 928
rect 6104 926 6106 928
rect 6134 926 6136 928
rect 3294 922 3296 924
rect 3704 922 3706 924
rect 3894 922 3896 924
rect 4304 922 4306 924
rect 6294 922 6296 924
rect 6704 922 6706 924
rect 3296 920 3298 922
rect 3702 920 3704 922
rect 3896 920 3898 922
rect 4302 920 4304 922
rect 4484 920 4486 922
rect 4514 920 4516 922
rect 4544 920 4546 922
rect 4574 920 4576 922
rect 4604 920 4606 922
rect 4634 920 4636 922
rect 4664 920 4666 922
rect 4694 920 4696 922
rect 4724 920 4726 922
rect 4754 920 4756 922
rect 4784 920 4786 922
rect 4814 920 4816 922
rect 4844 920 4846 922
rect 4874 920 4876 922
rect 4904 920 4906 922
rect 4934 920 4936 922
rect 5084 920 5086 922
rect 5114 920 5116 922
rect 5144 920 5146 922
rect 5174 920 5176 922
rect 5204 920 5206 922
rect 5234 920 5236 922
rect 5264 920 5266 922
rect 5294 920 5296 922
rect 5324 920 5326 922
rect 5354 920 5356 922
rect 5384 920 5386 922
rect 5414 920 5416 922
rect 5444 920 5446 922
rect 5474 920 5476 922
rect 5504 920 5506 922
rect 5534 920 5536 922
rect 5684 920 5686 922
rect 5714 920 5716 922
rect 5744 920 5746 922
rect 5774 920 5776 922
rect 5804 920 5806 922
rect 5834 920 5836 922
rect 5864 920 5866 922
rect 5894 920 5896 922
rect 5924 920 5926 922
rect 5954 920 5956 922
rect 5984 920 5986 922
rect 6014 920 6016 922
rect 6044 920 6046 922
rect 6074 920 6076 922
rect 6104 920 6106 922
rect 6134 920 6136 922
rect 6296 920 6298 922
rect 6702 920 6704 922
rect 3250 919 3252 920
rect 3748 919 3750 920
rect 3850 919 3852 920
rect 4348 919 4350 920
rect 4476 918 4478 920
rect 4482 918 4484 920
rect 4506 918 4508 920
rect 4512 918 4514 920
rect 4536 918 4538 920
rect 4542 918 4544 920
rect 4566 918 4568 920
rect 4572 918 4574 920
rect 4596 918 4598 920
rect 4602 918 4604 920
rect 4626 918 4628 920
rect 4632 918 4634 920
rect 4656 918 4658 920
rect 4662 918 4664 920
rect 4686 918 4688 920
rect 4692 918 4694 920
rect 4716 918 4718 920
rect 4722 918 4724 920
rect 4746 918 4748 920
rect 4752 918 4754 920
rect 4776 918 4778 920
rect 4782 918 4784 920
rect 4806 918 4808 920
rect 4812 918 4814 920
rect 4836 918 4838 920
rect 4842 918 4844 920
rect 4866 918 4868 920
rect 4872 918 4874 920
rect 4896 918 4898 920
rect 4902 918 4904 920
rect 4926 918 4928 920
rect 4932 918 4934 920
rect 5076 918 5078 920
rect 5082 918 5084 920
rect 5106 918 5108 920
rect 5112 918 5114 920
rect 5136 918 5138 920
rect 5142 918 5144 920
rect 5166 918 5168 920
rect 5172 918 5174 920
rect 5196 918 5198 920
rect 5202 918 5204 920
rect 5226 918 5228 920
rect 5232 918 5234 920
rect 5256 918 5258 920
rect 5262 918 5264 920
rect 5286 918 5288 920
rect 5292 918 5294 920
rect 5316 918 5318 920
rect 5322 918 5324 920
rect 5346 918 5348 920
rect 5352 918 5354 920
rect 5376 918 5378 920
rect 5382 918 5384 920
rect 5406 918 5408 920
rect 5412 918 5414 920
rect 5436 918 5438 920
rect 5442 918 5444 920
rect 5466 918 5468 920
rect 5472 918 5474 920
rect 5496 918 5498 920
rect 5502 918 5504 920
rect 5526 918 5528 920
rect 5532 918 5534 920
rect 5676 918 5678 920
rect 5682 918 5684 920
rect 5706 918 5708 920
rect 5712 918 5714 920
rect 5736 918 5738 920
rect 5742 918 5744 920
rect 5766 918 5768 920
rect 5772 918 5774 920
rect 5796 918 5798 920
rect 5802 918 5804 920
rect 5826 918 5828 920
rect 5832 918 5834 920
rect 5856 918 5858 920
rect 5862 918 5864 920
rect 5886 918 5888 920
rect 5892 918 5894 920
rect 5916 918 5918 920
rect 5922 918 5924 920
rect 5946 918 5948 920
rect 5952 918 5954 920
rect 5976 918 5978 920
rect 5982 918 5984 920
rect 6006 918 6008 920
rect 6012 918 6014 920
rect 6036 918 6038 920
rect 6042 918 6044 920
rect 6066 918 6068 920
rect 6072 918 6074 920
rect 6096 918 6098 920
rect 6102 918 6104 920
rect 6126 918 6128 920
rect 6132 918 6134 920
rect 6250 919 6252 920
rect 6748 919 6750 920
rect 3248 917 3250 918
rect 3750 917 3752 918
rect 3848 917 3850 918
rect 4350 917 4352 918
rect 4474 916 4476 918
rect 4504 916 4506 918
rect 4534 916 4536 918
rect 4564 916 4566 918
rect 4594 916 4596 918
rect 4624 916 4626 918
rect 4654 916 4656 918
rect 4684 916 4686 918
rect 4714 916 4716 918
rect 4744 916 4746 918
rect 4774 916 4776 918
rect 4804 916 4806 918
rect 4834 916 4836 918
rect 4864 916 4866 918
rect 4894 916 4896 918
rect 4924 916 4926 918
rect 5074 916 5076 918
rect 5104 916 5106 918
rect 5134 916 5136 918
rect 5164 916 5166 918
rect 5194 916 5196 918
rect 5224 916 5226 918
rect 5254 916 5256 918
rect 5284 916 5286 918
rect 5314 916 5316 918
rect 5344 916 5346 918
rect 5374 916 5376 918
rect 5404 916 5406 918
rect 5434 916 5436 918
rect 5464 916 5466 918
rect 5494 916 5496 918
rect 5524 916 5526 918
rect 5674 916 5676 918
rect 5704 916 5706 918
rect 5734 916 5736 918
rect 5764 916 5766 918
rect 5794 916 5796 918
rect 5824 916 5826 918
rect 5854 916 5856 918
rect 5884 916 5886 918
rect 5914 916 5916 918
rect 5944 916 5946 918
rect 5974 916 5976 918
rect 6004 916 6006 918
rect 6034 916 6036 918
rect 6064 916 6066 918
rect 6094 916 6096 918
rect 6124 916 6126 918
rect 6248 917 6250 918
rect 6750 917 6752 918
rect 4474 910 4476 912
rect 4504 910 4506 912
rect 4534 910 4536 912
rect 4564 910 4566 912
rect 4594 910 4596 912
rect 4624 910 4626 912
rect 4654 910 4656 912
rect 4684 910 4686 912
rect 4714 910 4716 912
rect 4744 910 4746 912
rect 4774 910 4776 912
rect 4804 910 4806 912
rect 4834 910 4836 912
rect 4864 910 4866 912
rect 4894 910 4896 912
rect 4924 910 4926 912
rect 5074 910 5076 912
rect 5104 910 5106 912
rect 5134 910 5136 912
rect 5164 910 5166 912
rect 5194 910 5196 912
rect 5224 910 5226 912
rect 5254 910 5256 912
rect 5284 910 5286 912
rect 5314 910 5316 912
rect 5344 910 5346 912
rect 5374 910 5376 912
rect 5404 910 5406 912
rect 5434 910 5436 912
rect 5464 910 5466 912
rect 5494 910 5496 912
rect 5524 910 5526 912
rect 5674 910 5676 912
rect 5704 910 5706 912
rect 5734 910 5736 912
rect 5764 910 5766 912
rect 5794 910 5796 912
rect 5824 910 5826 912
rect 5854 910 5856 912
rect 5884 910 5886 912
rect 5914 910 5916 912
rect 5944 910 5946 912
rect 5974 910 5976 912
rect 6004 910 6006 912
rect 6034 910 6036 912
rect 6064 910 6066 912
rect 6094 910 6096 912
rect 6124 910 6126 912
rect 4476 908 4478 910
rect 4482 908 4484 910
rect 4506 908 4508 910
rect 4512 908 4514 910
rect 4536 908 4538 910
rect 4542 908 4544 910
rect 4566 908 4568 910
rect 4572 908 4574 910
rect 4596 908 4598 910
rect 4602 908 4604 910
rect 4626 908 4628 910
rect 4632 908 4634 910
rect 4656 908 4658 910
rect 4662 908 4664 910
rect 4686 908 4688 910
rect 4692 908 4694 910
rect 4716 908 4718 910
rect 4722 908 4724 910
rect 4746 908 4748 910
rect 4752 908 4754 910
rect 4776 908 4778 910
rect 4782 908 4784 910
rect 4806 908 4808 910
rect 4812 908 4814 910
rect 4836 908 4838 910
rect 4842 908 4844 910
rect 4866 908 4868 910
rect 4872 908 4874 910
rect 4896 908 4898 910
rect 4902 908 4904 910
rect 4926 908 4928 910
rect 4932 908 4934 910
rect 5076 908 5078 910
rect 5082 908 5084 910
rect 5106 908 5108 910
rect 5112 908 5114 910
rect 5136 908 5138 910
rect 5142 908 5144 910
rect 5166 908 5168 910
rect 5172 908 5174 910
rect 5196 908 5198 910
rect 5202 908 5204 910
rect 5226 908 5228 910
rect 5232 908 5234 910
rect 5256 908 5258 910
rect 5262 908 5264 910
rect 5286 908 5288 910
rect 5292 908 5294 910
rect 5316 908 5318 910
rect 5322 908 5324 910
rect 5346 908 5348 910
rect 5352 908 5354 910
rect 5376 908 5378 910
rect 5382 908 5384 910
rect 5406 908 5408 910
rect 5412 908 5414 910
rect 5436 908 5438 910
rect 5442 908 5444 910
rect 5466 908 5468 910
rect 5472 908 5474 910
rect 5496 908 5498 910
rect 5502 908 5504 910
rect 5526 908 5528 910
rect 5532 908 5534 910
rect 5676 908 5678 910
rect 5682 908 5684 910
rect 5706 908 5708 910
rect 5712 908 5714 910
rect 5736 908 5738 910
rect 5742 908 5744 910
rect 5766 908 5768 910
rect 5772 908 5774 910
rect 5796 908 5798 910
rect 5802 908 5804 910
rect 5826 908 5828 910
rect 5832 908 5834 910
rect 5856 908 5858 910
rect 5862 908 5864 910
rect 5886 908 5888 910
rect 5892 908 5894 910
rect 5916 908 5918 910
rect 5922 908 5924 910
rect 5946 908 5948 910
rect 5952 908 5954 910
rect 5976 908 5978 910
rect 5982 908 5984 910
rect 6006 908 6008 910
rect 6012 908 6014 910
rect 6036 908 6038 910
rect 6042 908 6044 910
rect 6066 908 6068 910
rect 6072 908 6074 910
rect 6096 908 6098 910
rect 6102 908 6104 910
rect 6126 908 6128 910
rect 6132 908 6134 910
rect 4484 906 4486 908
rect 4514 906 4516 908
rect 4544 906 4546 908
rect 4574 906 4576 908
rect 4604 906 4606 908
rect 4634 906 4636 908
rect 4664 906 4666 908
rect 4694 906 4696 908
rect 4724 906 4726 908
rect 4754 906 4756 908
rect 4784 906 4786 908
rect 4814 906 4816 908
rect 4844 906 4846 908
rect 4874 906 4876 908
rect 4904 906 4906 908
rect 4934 906 4936 908
rect 5084 906 5086 908
rect 5114 906 5116 908
rect 5144 906 5146 908
rect 5174 906 5176 908
rect 5204 906 5206 908
rect 5234 906 5236 908
rect 5264 906 5266 908
rect 5294 906 5296 908
rect 5324 906 5326 908
rect 5354 906 5356 908
rect 5384 906 5386 908
rect 5414 906 5416 908
rect 5444 906 5446 908
rect 5474 906 5476 908
rect 5504 906 5506 908
rect 5534 906 5536 908
rect 5684 906 5686 908
rect 5714 906 5716 908
rect 5744 906 5746 908
rect 5774 906 5776 908
rect 5804 906 5806 908
rect 5834 906 5836 908
rect 5864 906 5866 908
rect 5894 906 5896 908
rect 5924 906 5926 908
rect 5954 906 5956 908
rect 5984 906 5986 908
rect 6014 906 6016 908
rect 6044 906 6046 908
rect 6074 906 6076 908
rect 6104 906 6106 908
rect 6134 906 6136 908
rect 4484 900 4486 902
rect 4514 900 4516 902
rect 4544 900 4546 902
rect 4574 900 4576 902
rect 4604 900 4606 902
rect 4634 900 4636 902
rect 4664 900 4666 902
rect 4694 900 4696 902
rect 4724 900 4726 902
rect 4754 900 4756 902
rect 4784 900 4786 902
rect 4814 900 4816 902
rect 4844 900 4846 902
rect 4874 900 4876 902
rect 4904 900 4906 902
rect 4934 900 4936 902
rect 5084 900 5086 902
rect 5114 900 5116 902
rect 5144 900 5146 902
rect 5174 900 5176 902
rect 5204 900 5206 902
rect 5234 900 5236 902
rect 5264 900 5266 902
rect 5294 900 5296 902
rect 5324 900 5326 902
rect 5354 900 5356 902
rect 5384 900 5386 902
rect 5414 900 5416 902
rect 5444 900 5446 902
rect 5474 900 5476 902
rect 5504 900 5506 902
rect 5534 900 5536 902
rect 5684 900 5686 902
rect 5714 900 5716 902
rect 5744 900 5746 902
rect 5774 900 5776 902
rect 5804 900 5806 902
rect 5834 900 5836 902
rect 5864 900 5866 902
rect 5894 900 5896 902
rect 5924 900 5926 902
rect 5954 900 5956 902
rect 5984 900 5986 902
rect 6014 900 6016 902
rect 6044 900 6046 902
rect 6074 900 6076 902
rect 6104 900 6106 902
rect 6134 900 6136 902
rect 3250 899 3252 900
rect 3748 899 3750 900
rect 3850 899 3852 900
rect 4348 899 4350 900
rect 4476 898 4478 900
rect 4482 898 4484 900
rect 4506 898 4508 900
rect 4512 898 4514 900
rect 4536 898 4538 900
rect 4542 898 4544 900
rect 4566 898 4568 900
rect 4572 898 4574 900
rect 4596 898 4598 900
rect 4602 898 4604 900
rect 4626 898 4628 900
rect 4632 898 4634 900
rect 4656 898 4658 900
rect 4662 898 4664 900
rect 4686 898 4688 900
rect 4692 898 4694 900
rect 4716 898 4718 900
rect 4722 898 4724 900
rect 4746 898 4748 900
rect 4752 898 4754 900
rect 4776 898 4778 900
rect 4782 898 4784 900
rect 4806 898 4808 900
rect 4812 898 4814 900
rect 4836 898 4838 900
rect 4842 898 4844 900
rect 4866 898 4868 900
rect 4872 898 4874 900
rect 4896 898 4898 900
rect 4902 898 4904 900
rect 4926 898 4928 900
rect 4932 898 4934 900
rect 5076 898 5078 900
rect 5082 898 5084 900
rect 5106 898 5108 900
rect 5112 898 5114 900
rect 5136 898 5138 900
rect 5142 898 5144 900
rect 5166 898 5168 900
rect 5172 898 5174 900
rect 5196 898 5198 900
rect 5202 898 5204 900
rect 5226 898 5228 900
rect 5232 898 5234 900
rect 5256 898 5258 900
rect 5262 898 5264 900
rect 5286 898 5288 900
rect 5292 898 5294 900
rect 5316 898 5318 900
rect 5322 898 5324 900
rect 5346 898 5348 900
rect 5352 898 5354 900
rect 5376 898 5378 900
rect 5382 898 5384 900
rect 5406 898 5408 900
rect 5412 898 5414 900
rect 5436 898 5438 900
rect 5442 898 5444 900
rect 5466 898 5468 900
rect 5472 898 5474 900
rect 5496 898 5498 900
rect 5502 898 5504 900
rect 5526 898 5528 900
rect 5532 898 5534 900
rect 5676 898 5678 900
rect 5682 898 5684 900
rect 5706 898 5708 900
rect 5712 898 5714 900
rect 5736 898 5738 900
rect 5742 898 5744 900
rect 5766 898 5768 900
rect 5772 898 5774 900
rect 5796 898 5798 900
rect 5802 898 5804 900
rect 5826 898 5828 900
rect 5832 898 5834 900
rect 5856 898 5858 900
rect 5862 898 5864 900
rect 5886 898 5888 900
rect 5892 898 5894 900
rect 5916 898 5918 900
rect 5922 898 5924 900
rect 5946 898 5948 900
rect 5952 898 5954 900
rect 5976 898 5978 900
rect 5982 898 5984 900
rect 6006 898 6008 900
rect 6012 898 6014 900
rect 6036 898 6038 900
rect 6042 898 6044 900
rect 6066 898 6068 900
rect 6072 898 6074 900
rect 6096 898 6098 900
rect 6102 898 6104 900
rect 6126 898 6128 900
rect 6132 898 6134 900
rect 6250 899 6252 900
rect 6748 899 6750 900
rect 3248 897 3250 898
rect 3750 897 3752 898
rect 3848 897 3850 898
rect 4350 897 4352 898
rect 4094 895 4096 897
rect 4104 895 4106 897
rect 4474 896 4476 898
rect 4504 896 4506 898
rect 4534 896 4536 898
rect 4564 896 4566 898
rect 4594 896 4596 898
rect 4624 896 4626 898
rect 4654 896 4656 898
rect 4684 896 4686 898
rect 4714 896 4716 898
rect 4744 896 4746 898
rect 4774 896 4776 898
rect 4804 896 4806 898
rect 4834 896 4836 898
rect 4864 896 4866 898
rect 4894 896 4896 898
rect 4924 896 4926 898
rect 5074 896 5076 898
rect 5104 896 5106 898
rect 5134 896 5136 898
rect 5164 896 5166 898
rect 5194 896 5196 898
rect 5224 896 5226 898
rect 5254 896 5256 898
rect 5284 896 5286 898
rect 5314 896 5316 898
rect 5344 896 5346 898
rect 5374 896 5376 898
rect 5404 896 5406 898
rect 5434 896 5436 898
rect 5464 896 5466 898
rect 5494 896 5496 898
rect 5524 896 5526 898
rect 5674 896 5676 898
rect 5704 896 5706 898
rect 5734 896 5736 898
rect 5764 896 5766 898
rect 5794 896 5796 898
rect 5824 896 5826 898
rect 5854 896 5856 898
rect 5884 896 5886 898
rect 5914 896 5916 898
rect 5944 896 5946 898
rect 5974 896 5976 898
rect 6004 896 6006 898
rect 6034 896 6036 898
rect 6064 896 6066 898
rect 6094 896 6096 898
rect 6124 896 6126 898
rect 6248 897 6250 898
rect 6750 897 6752 898
rect 4092 893 4094 895
rect 4106 893 4108 895
rect 4474 890 4476 892
rect 4504 890 4506 892
rect 4534 890 4536 892
rect 4564 890 4566 892
rect 4594 890 4596 892
rect 4624 890 4626 892
rect 4654 890 4656 892
rect 4684 890 4686 892
rect 4714 890 4716 892
rect 4744 890 4746 892
rect 4774 890 4776 892
rect 4804 890 4806 892
rect 4834 890 4836 892
rect 4864 890 4866 892
rect 4894 890 4896 892
rect 4924 890 4926 892
rect 5074 890 5076 892
rect 5104 890 5106 892
rect 5134 890 5136 892
rect 5164 890 5166 892
rect 5194 890 5196 892
rect 5224 890 5226 892
rect 5254 890 5256 892
rect 5284 890 5286 892
rect 5314 890 5316 892
rect 5344 890 5346 892
rect 5374 890 5376 892
rect 5404 890 5406 892
rect 5434 890 5436 892
rect 5464 890 5466 892
rect 5494 890 5496 892
rect 5524 890 5526 892
rect 5674 890 5676 892
rect 5704 890 5706 892
rect 5734 890 5736 892
rect 5764 890 5766 892
rect 5794 890 5796 892
rect 5824 890 5826 892
rect 5854 890 5856 892
rect 5884 890 5886 892
rect 5914 890 5916 892
rect 5944 890 5946 892
rect 5974 890 5976 892
rect 6004 890 6006 892
rect 6034 890 6036 892
rect 6064 890 6066 892
rect 6094 890 6096 892
rect 6124 890 6126 892
rect 4476 888 4478 890
rect 4482 888 4484 890
rect 4506 888 4508 890
rect 4512 888 4514 890
rect 4536 888 4538 890
rect 4542 888 4544 890
rect 4566 888 4568 890
rect 4572 888 4574 890
rect 4596 888 4598 890
rect 4602 888 4604 890
rect 4626 888 4628 890
rect 4632 888 4634 890
rect 4656 888 4658 890
rect 4662 888 4664 890
rect 4686 888 4688 890
rect 4692 888 4694 890
rect 4716 888 4718 890
rect 4722 888 4724 890
rect 4746 888 4748 890
rect 4752 888 4754 890
rect 4776 888 4778 890
rect 4782 888 4784 890
rect 4806 888 4808 890
rect 4812 888 4814 890
rect 4836 888 4838 890
rect 4842 888 4844 890
rect 4866 888 4868 890
rect 4872 888 4874 890
rect 4896 888 4898 890
rect 4902 888 4904 890
rect 4926 888 4928 890
rect 4932 888 4934 890
rect 5076 888 5078 890
rect 5082 888 5084 890
rect 5106 888 5108 890
rect 5112 888 5114 890
rect 5136 888 5138 890
rect 5142 888 5144 890
rect 5166 888 5168 890
rect 5172 888 5174 890
rect 5196 888 5198 890
rect 5202 888 5204 890
rect 5226 888 5228 890
rect 5232 888 5234 890
rect 5256 888 5258 890
rect 5262 888 5264 890
rect 5286 888 5288 890
rect 5292 888 5294 890
rect 5316 888 5318 890
rect 5322 888 5324 890
rect 5346 888 5348 890
rect 5352 888 5354 890
rect 5376 888 5378 890
rect 5382 888 5384 890
rect 5406 888 5408 890
rect 5412 888 5414 890
rect 5436 888 5438 890
rect 5442 888 5444 890
rect 5466 888 5468 890
rect 5472 888 5474 890
rect 5496 888 5498 890
rect 5502 888 5504 890
rect 5526 888 5528 890
rect 5532 888 5534 890
rect 5676 888 5678 890
rect 5682 888 5684 890
rect 5706 888 5708 890
rect 5712 888 5714 890
rect 5736 888 5738 890
rect 5742 888 5744 890
rect 5766 888 5768 890
rect 5772 888 5774 890
rect 5796 888 5798 890
rect 5802 888 5804 890
rect 5826 888 5828 890
rect 5832 888 5834 890
rect 5856 888 5858 890
rect 5862 888 5864 890
rect 5886 888 5888 890
rect 5892 888 5894 890
rect 5916 888 5918 890
rect 5922 888 5924 890
rect 5946 888 5948 890
rect 5952 888 5954 890
rect 5976 888 5978 890
rect 5982 888 5984 890
rect 6006 888 6008 890
rect 6012 888 6014 890
rect 6036 888 6038 890
rect 6042 888 6044 890
rect 6066 888 6068 890
rect 6072 888 6074 890
rect 6096 888 6098 890
rect 6102 888 6104 890
rect 6126 888 6128 890
rect 6132 888 6134 890
rect 4484 886 4486 888
rect 4514 886 4516 888
rect 4544 886 4546 888
rect 4574 886 4576 888
rect 4604 886 4606 888
rect 4634 886 4636 888
rect 4664 886 4666 888
rect 4694 886 4696 888
rect 4724 886 4726 888
rect 4754 886 4756 888
rect 4784 886 4786 888
rect 4814 886 4816 888
rect 4844 886 4846 888
rect 4874 886 4876 888
rect 4904 886 4906 888
rect 4934 886 4936 888
rect 5084 886 5086 888
rect 5114 886 5116 888
rect 5144 886 5146 888
rect 5174 886 5176 888
rect 5204 886 5206 888
rect 5234 886 5236 888
rect 5264 886 5266 888
rect 5294 886 5296 888
rect 5324 886 5326 888
rect 5354 886 5356 888
rect 5384 886 5386 888
rect 5414 886 5416 888
rect 5444 886 5446 888
rect 5474 886 5476 888
rect 5504 886 5506 888
rect 5534 886 5536 888
rect 5684 886 5686 888
rect 5714 886 5716 888
rect 5744 886 5746 888
rect 5774 886 5776 888
rect 5804 886 5806 888
rect 5834 886 5836 888
rect 5864 886 5866 888
rect 5894 886 5896 888
rect 5924 886 5926 888
rect 5954 886 5956 888
rect 5984 886 5986 888
rect 6014 886 6016 888
rect 6044 886 6046 888
rect 6074 886 6076 888
rect 6104 886 6106 888
rect 6134 886 6136 888
rect 1702 884 1704 886
rect 1732 884 1734 886
rect 1700 882 1702 884
rect 1734 882 1736 884
rect 4456 878 4458 880
rect 4462 878 4464 880
rect 4476 878 4478 880
rect 4492 878 4494 880
rect 4506 878 4508 880
rect 4522 878 4524 880
rect 4536 878 4538 880
rect 4552 878 4554 880
rect 4566 878 4568 880
rect 4582 878 4584 880
rect 4596 878 4598 880
rect 4612 878 4614 880
rect 4626 878 4628 880
rect 4642 878 4644 880
rect 4656 878 4658 880
rect 4672 878 4674 880
rect 4686 878 4688 880
rect 4702 878 4704 880
rect 4716 878 4718 880
rect 4732 878 4734 880
rect 4746 878 4748 880
rect 4762 878 4764 880
rect 4776 878 4778 880
rect 4792 878 4794 880
rect 4806 878 4808 880
rect 4822 878 4824 880
rect 4836 878 4838 880
rect 4852 878 4854 880
rect 4866 878 4868 880
rect 4882 878 4884 880
rect 4896 878 4898 880
rect 4912 878 4914 880
rect 4926 878 4928 880
rect 4942 878 4944 880
rect 5056 878 5058 880
rect 5062 878 5064 880
rect 5076 878 5078 880
rect 5092 878 5094 880
rect 5106 878 5108 880
rect 5122 878 5124 880
rect 5136 878 5138 880
rect 5152 878 5154 880
rect 5166 878 5168 880
rect 5182 878 5184 880
rect 5196 878 5198 880
rect 5212 878 5214 880
rect 5226 878 5228 880
rect 5242 878 5244 880
rect 5256 878 5258 880
rect 5272 878 5274 880
rect 5286 878 5288 880
rect 5302 878 5304 880
rect 5316 878 5318 880
rect 5332 878 5334 880
rect 5346 878 5348 880
rect 5362 878 5364 880
rect 5376 878 5378 880
rect 5392 878 5394 880
rect 5406 878 5408 880
rect 5422 878 5424 880
rect 5436 878 5438 880
rect 5452 878 5454 880
rect 5466 878 5468 880
rect 5482 878 5484 880
rect 5496 878 5498 880
rect 5512 878 5514 880
rect 5526 878 5528 880
rect 5542 878 5544 880
rect 5656 878 5658 880
rect 5662 878 5664 880
rect 5676 878 5678 880
rect 5692 878 5694 880
rect 5706 878 5708 880
rect 5722 878 5724 880
rect 5736 878 5738 880
rect 5752 878 5754 880
rect 5766 878 5768 880
rect 5782 878 5784 880
rect 5796 878 5798 880
rect 5812 878 5814 880
rect 5826 878 5828 880
rect 5842 878 5844 880
rect 5856 878 5858 880
rect 5872 878 5874 880
rect 5886 878 5888 880
rect 5902 878 5904 880
rect 5916 878 5918 880
rect 5932 878 5934 880
rect 5946 878 5948 880
rect 5962 878 5964 880
rect 5976 878 5978 880
rect 5992 878 5994 880
rect 6006 878 6008 880
rect 6022 878 6024 880
rect 6036 878 6038 880
rect 6052 878 6054 880
rect 6066 878 6068 880
rect 6082 878 6084 880
rect 6096 878 6098 880
rect 6112 878 6114 880
rect 6126 878 6128 880
rect 6142 878 6144 880
rect 4454 876 4456 878
rect 4464 876 4466 878
rect 4474 876 4476 878
rect 4494 876 4496 878
rect 4504 876 4506 878
rect 4524 876 4526 878
rect 4534 876 4536 878
rect 4554 876 4556 878
rect 4564 876 4566 878
rect 4584 876 4586 878
rect 4594 876 4596 878
rect 4614 876 4616 878
rect 4624 876 4626 878
rect 4644 876 4646 878
rect 4654 876 4656 878
rect 4674 876 4676 878
rect 4684 876 4686 878
rect 4704 876 4706 878
rect 4714 876 4716 878
rect 4734 876 4736 878
rect 4744 876 4746 878
rect 4764 876 4766 878
rect 4774 876 4776 878
rect 4794 876 4796 878
rect 4804 876 4806 878
rect 4824 876 4826 878
rect 4834 876 4836 878
rect 4854 876 4856 878
rect 4864 876 4866 878
rect 4884 876 4886 878
rect 4894 876 4896 878
rect 4914 876 4916 878
rect 4924 876 4926 878
rect 4944 876 4946 878
rect 5054 876 5056 878
rect 5064 876 5066 878
rect 5074 876 5076 878
rect 5094 876 5096 878
rect 5104 876 5106 878
rect 5124 876 5126 878
rect 5134 876 5136 878
rect 5154 876 5156 878
rect 5164 876 5166 878
rect 5184 876 5186 878
rect 5194 876 5196 878
rect 5214 876 5216 878
rect 5224 876 5226 878
rect 5244 876 5246 878
rect 5254 876 5256 878
rect 5274 876 5276 878
rect 5284 876 5286 878
rect 5304 876 5306 878
rect 5314 876 5316 878
rect 5334 876 5336 878
rect 5344 876 5346 878
rect 5364 876 5366 878
rect 5374 876 5376 878
rect 5394 876 5396 878
rect 5404 876 5406 878
rect 5424 876 5426 878
rect 5434 876 5436 878
rect 5454 876 5456 878
rect 5464 876 5466 878
rect 5484 876 5486 878
rect 5494 876 5496 878
rect 5514 876 5516 878
rect 5524 876 5526 878
rect 5544 876 5546 878
rect 5654 876 5656 878
rect 5664 876 5666 878
rect 5674 876 5676 878
rect 5694 876 5696 878
rect 5704 876 5706 878
rect 5724 876 5726 878
rect 5734 876 5736 878
rect 5754 876 5756 878
rect 5764 876 5766 878
rect 5784 876 5786 878
rect 5794 876 5796 878
rect 5814 876 5816 878
rect 5824 876 5826 878
rect 5844 876 5846 878
rect 5854 876 5856 878
rect 5874 876 5876 878
rect 5884 876 5886 878
rect 5904 876 5906 878
rect 5914 876 5916 878
rect 5934 876 5936 878
rect 5944 876 5946 878
rect 5964 876 5966 878
rect 5974 876 5976 878
rect 5994 876 5996 878
rect 6004 876 6006 878
rect 6024 876 6026 878
rect 6034 876 6036 878
rect 6054 876 6056 878
rect 6064 876 6066 878
rect 6084 876 6086 878
rect 6094 876 6096 878
rect 6114 876 6116 878
rect 6124 876 6126 878
rect 6144 876 6146 878
rect 1692 874 1694 876
rect 1690 872 1692 874
rect 3262 873 3264 875
rect 3736 873 3738 875
rect 3862 873 3864 875
rect 4336 873 4338 875
rect 6262 873 6264 875
rect 6736 873 6738 875
rect 3260 871 3262 873
rect 3738 871 3740 873
rect 3860 871 3862 873
rect 4338 871 4340 873
rect 6260 871 6262 873
rect 6738 871 6740 873
rect 1682 864 1684 866
rect 1680 862 1682 864
rect 1734 862 1736 864
rect 1732 860 1734 862
rect 1672 854 1674 856
rect 1670 852 1672 854
rect 1724 852 1726 854
rect 1722 850 1724 852
rect 1662 844 1664 846
rect 1722 844 1724 846
rect 1732 844 1734 846
rect 1752 844 1754 846
rect 1762 844 1764 846
rect 1782 844 1784 846
rect 1792 844 1794 846
rect 1812 844 1814 846
rect 1822 844 1824 846
rect 1842 844 1844 846
rect 1852 844 1854 846
rect 1872 844 1874 846
rect 1882 844 1884 846
rect 1902 844 1904 846
rect 1912 844 1914 846
rect 1932 844 1934 846
rect 1942 844 1944 846
rect 1962 844 1964 846
rect 1972 844 1974 846
rect 1660 842 1662 844
rect 1714 842 1716 844
rect 1720 842 1722 844
rect 1734 842 1736 844
rect 1750 842 1752 844
rect 1764 842 1766 844
rect 1780 842 1782 844
rect 1794 842 1796 844
rect 1810 842 1812 844
rect 1824 842 1826 844
rect 1840 842 1842 844
rect 1854 842 1856 844
rect 1870 842 1872 844
rect 1884 842 1886 844
rect 1900 842 1902 844
rect 1914 842 1916 844
rect 1930 842 1932 844
rect 1944 842 1946 844
rect 1960 842 1962 844
rect 1974 842 1976 844
rect 1712 840 1714 842
rect 1652 834 1654 836
rect 1742 834 1744 836
rect 1772 834 1774 836
rect 1802 834 1804 836
rect 1832 834 1834 836
rect 1862 834 1864 836
rect 1892 834 1894 836
rect 1922 834 1924 836
rect 1952 834 1954 836
rect 1982 834 1984 836
rect 1650 832 1652 834
rect 1704 832 1706 834
rect 1720 832 1722 834
rect 1744 832 1746 834
rect 1750 832 1752 834
rect 1774 832 1776 834
rect 1780 832 1782 834
rect 1804 832 1806 834
rect 1810 832 1812 834
rect 1834 832 1836 834
rect 1840 832 1842 834
rect 1864 832 1866 834
rect 1870 832 1872 834
rect 1894 832 1896 834
rect 1900 832 1902 834
rect 1924 832 1926 834
rect 1930 832 1932 834
rect 1954 832 1956 834
rect 1960 832 1962 834
rect 1984 832 1986 834
rect 1702 830 1704 832
rect 1722 830 1724 832
rect 1752 830 1754 832
rect 1782 830 1784 832
rect 1812 830 1814 832
rect 1842 830 1844 832
rect 1872 830 1874 832
rect 1902 830 1904 832
rect 1932 830 1934 832
rect 1962 830 1964 832
rect 3232 828 3234 830
rect 3262 828 3264 830
rect 3292 828 3294 830
rect 3322 828 3324 830
rect 3352 828 3354 830
rect 3382 828 3384 830
rect 3616 828 3618 830
rect 3646 828 3648 830
rect 3676 828 3678 830
rect 3706 828 3708 830
rect 3736 828 3738 830
rect 3766 828 3768 830
rect 3832 828 3834 830
rect 3862 828 3864 830
rect 3892 828 3894 830
rect 3922 828 3924 830
rect 3952 828 3954 830
rect 3982 828 3984 830
rect 4216 828 4218 830
rect 4246 828 4248 830
rect 4276 828 4278 830
rect 4306 828 4308 830
rect 4336 828 4338 830
rect 4366 828 4368 830
rect 4432 828 4434 830
rect 4462 828 4464 830
rect 4492 828 4494 830
rect 4522 828 4524 830
rect 4552 828 4554 830
rect 4582 828 4584 830
rect 4612 828 4614 830
rect 4684 828 4686 830
rect 4714 828 4716 830
rect 4786 828 4788 830
rect 4816 828 4818 830
rect 4846 828 4848 830
rect 4876 828 4878 830
rect 4906 828 4908 830
rect 4936 828 4938 830
rect 4966 828 4968 830
rect 5032 828 5034 830
rect 5062 828 5064 830
rect 5092 828 5094 830
rect 5122 828 5124 830
rect 5152 828 5154 830
rect 5182 828 5184 830
rect 5212 828 5214 830
rect 5284 828 5286 830
rect 5314 828 5316 830
rect 5386 828 5388 830
rect 5416 828 5418 830
rect 5446 828 5448 830
rect 5476 828 5478 830
rect 5506 828 5508 830
rect 5536 828 5538 830
rect 5566 828 5568 830
rect 5632 828 5634 830
rect 5662 828 5664 830
rect 5692 828 5694 830
rect 5722 828 5724 830
rect 5752 828 5754 830
rect 6046 828 6048 830
rect 6076 828 6078 830
rect 6106 828 6108 830
rect 6136 828 6138 830
rect 6166 828 6168 830
rect 6232 828 6234 830
rect 6262 828 6264 830
rect 6292 828 6294 830
rect 6322 828 6324 830
rect 6352 828 6354 830
rect 6382 828 6384 830
rect 6412 828 6414 830
rect 6586 828 6588 830
rect 6616 828 6618 830
rect 6646 828 6648 830
rect 6676 828 6678 830
rect 6706 828 6708 830
rect 6736 828 6738 830
rect 6766 828 6768 830
rect 3234 826 3236 828
rect 3240 826 3242 828
rect 3264 826 3266 828
rect 3270 826 3272 828
rect 3294 826 3296 828
rect 3300 826 3302 828
rect 3324 826 3326 828
rect 3330 826 3332 828
rect 3354 826 3356 828
rect 3360 826 3362 828
rect 3384 826 3386 828
rect 3614 826 3616 828
rect 3638 826 3640 828
rect 3644 826 3646 828
rect 3668 826 3670 828
rect 3674 826 3676 828
rect 3698 826 3700 828
rect 3704 826 3706 828
rect 3728 826 3730 828
rect 3734 826 3736 828
rect 3758 826 3760 828
rect 3764 826 3766 828
rect 3834 826 3836 828
rect 3840 826 3842 828
rect 3864 826 3866 828
rect 3870 826 3872 828
rect 3894 826 3896 828
rect 3900 826 3902 828
rect 3924 826 3926 828
rect 3930 826 3932 828
rect 3954 826 3956 828
rect 3960 826 3962 828
rect 3984 826 3986 828
rect 4214 826 4216 828
rect 4238 826 4240 828
rect 4244 826 4246 828
rect 4268 826 4270 828
rect 4274 826 4276 828
rect 4298 826 4300 828
rect 4304 826 4306 828
rect 4328 826 4330 828
rect 4334 826 4336 828
rect 4358 826 4360 828
rect 4364 826 4366 828
rect 4434 826 4436 828
rect 4440 826 4442 828
rect 4464 826 4466 828
rect 4470 826 4472 828
rect 4494 826 4496 828
rect 4500 826 4502 828
rect 4524 826 4526 828
rect 4530 826 4532 828
rect 4554 826 4556 828
rect 4560 826 4562 828
rect 4584 826 4586 828
rect 4590 826 4592 828
rect 4614 826 4616 828
rect 4620 826 4622 828
rect 4686 826 4688 828
rect 4692 826 4694 828
rect 4716 826 4718 828
rect 4722 826 4724 828
rect 4778 826 4780 828
rect 4784 826 4786 828
rect 4808 826 4810 828
rect 4814 826 4816 828
rect 4838 826 4840 828
rect 4844 826 4846 828
rect 4868 826 4870 828
rect 4874 826 4876 828
rect 4898 826 4900 828
rect 4904 826 4906 828
rect 4928 826 4930 828
rect 4934 826 4936 828
rect 4958 826 4960 828
rect 4964 826 4966 828
rect 5034 826 5036 828
rect 5040 826 5042 828
rect 5064 826 5066 828
rect 5070 826 5072 828
rect 5094 826 5096 828
rect 5100 826 5102 828
rect 5124 826 5126 828
rect 5130 826 5132 828
rect 5154 826 5156 828
rect 5160 826 5162 828
rect 5184 826 5186 828
rect 5190 826 5192 828
rect 5214 826 5216 828
rect 5220 826 5222 828
rect 5286 826 5288 828
rect 5292 826 5294 828
rect 5316 826 5318 828
rect 5322 826 5324 828
rect 5378 826 5380 828
rect 5384 826 5386 828
rect 5408 826 5410 828
rect 5414 826 5416 828
rect 5438 826 5440 828
rect 5444 826 5446 828
rect 5468 826 5470 828
rect 5474 826 5476 828
rect 5498 826 5500 828
rect 5504 826 5506 828
rect 5528 826 5530 828
rect 5534 826 5536 828
rect 5558 826 5560 828
rect 5564 826 5566 828
rect 5634 826 5636 828
rect 5640 826 5642 828
rect 5664 826 5666 828
rect 5670 826 5672 828
rect 5694 826 5696 828
rect 5700 826 5702 828
rect 5724 826 5726 828
rect 5730 826 5732 828
rect 5754 826 5756 828
rect 5760 826 5762 828
rect 6038 826 6040 828
rect 6044 826 6046 828
rect 6068 826 6070 828
rect 6074 826 6076 828
rect 6098 826 6100 828
rect 6104 826 6106 828
rect 6128 826 6130 828
rect 6134 826 6136 828
rect 6158 826 6160 828
rect 6164 826 6166 828
rect 6234 826 6236 828
rect 6240 826 6242 828
rect 6264 826 6266 828
rect 6270 826 6272 828
rect 6294 826 6296 828
rect 6300 826 6302 828
rect 6324 826 6326 828
rect 6330 826 6332 828
rect 6354 826 6356 828
rect 6360 826 6362 828
rect 6384 826 6386 828
rect 6390 826 6392 828
rect 6414 826 6416 828
rect 6420 826 6422 828
rect 6578 826 6580 828
rect 6584 826 6586 828
rect 6608 826 6610 828
rect 6614 826 6616 828
rect 6638 826 6640 828
rect 6644 826 6646 828
rect 6668 826 6670 828
rect 6674 826 6676 828
rect 6698 826 6700 828
rect 6704 826 6706 828
rect 6728 826 6730 828
rect 6734 826 6736 828
rect 6758 826 6760 828
rect 6764 826 6766 828
rect 1642 824 1644 826
rect 1722 824 1724 826
rect 1752 824 1754 826
rect 1782 824 1784 826
rect 1812 824 1814 826
rect 1842 824 1844 826
rect 1872 824 1874 826
rect 1902 824 1904 826
rect 1932 824 1934 826
rect 1962 824 1964 826
rect 3242 824 3244 826
rect 3272 824 3274 826
rect 3302 824 3304 826
rect 3332 824 3334 826
rect 3362 824 3364 826
rect 3636 824 3638 826
rect 3666 824 3668 826
rect 3696 824 3698 826
rect 3726 824 3728 826
rect 3756 824 3758 826
rect 3842 824 3844 826
rect 3872 824 3874 826
rect 3902 824 3904 826
rect 3932 824 3934 826
rect 3962 824 3964 826
rect 4236 824 4238 826
rect 4266 824 4268 826
rect 4296 824 4298 826
rect 4326 824 4328 826
rect 4356 824 4358 826
rect 4442 824 4444 826
rect 4472 824 4474 826
rect 4502 824 4504 826
rect 4532 824 4534 826
rect 4562 824 4564 826
rect 4592 824 4594 826
rect 4622 824 4624 826
rect 4694 824 4696 826
rect 4724 824 4726 826
rect 4776 824 4778 826
rect 4806 824 4808 826
rect 4836 824 4838 826
rect 4866 824 4868 826
rect 4896 824 4898 826
rect 4926 824 4928 826
rect 4956 824 4958 826
rect 5042 824 5044 826
rect 5072 824 5074 826
rect 5102 824 5104 826
rect 5132 824 5134 826
rect 5162 824 5164 826
rect 5192 824 5194 826
rect 5222 824 5224 826
rect 5294 824 5296 826
rect 5324 824 5326 826
rect 5376 824 5378 826
rect 5406 824 5408 826
rect 5436 824 5438 826
rect 5466 824 5468 826
rect 5496 824 5498 826
rect 5526 824 5528 826
rect 5556 824 5558 826
rect 5642 824 5644 826
rect 5672 824 5674 826
rect 5702 824 5704 826
rect 5732 824 5734 826
rect 5762 824 5764 826
rect 6036 824 6038 826
rect 6066 824 6068 826
rect 6096 824 6098 826
rect 6126 824 6128 826
rect 6156 824 6158 826
rect 6242 824 6244 826
rect 6272 824 6274 826
rect 6302 824 6304 826
rect 6332 824 6334 826
rect 6362 824 6364 826
rect 6392 824 6394 826
rect 6422 824 6424 826
rect 6576 824 6578 826
rect 6606 824 6608 826
rect 6636 824 6638 826
rect 6666 824 6668 826
rect 6696 824 6698 826
rect 6726 824 6728 826
rect 6756 824 6758 826
rect 1640 822 1642 824
rect 1694 822 1696 824
rect 1720 822 1722 824
rect 1744 822 1746 824
rect 1750 822 1752 824
rect 1774 822 1776 824
rect 1780 822 1782 824
rect 1804 822 1806 824
rect 1810 822 1812 824
rect 1834 822 1836 824
rect 1840 822 1842 824
rect 1864 822 1866 824
rect 1870 822 1872 824
rect 1894 822 1896 824
rect 1900 822 1902 824
rect 1924 822 1926 824
rect 1930 822 1932 824
rect 1954 822 1956 824
rect 1960 822 1962 824
rect 1984 822 1986 824
rect 1692 820 1694 822
rect 1742 820 1744 822
rect 1772 820 1774 822
rect 1802 820 1804 822
rect 1832 820 1834 822
rect 1862 820 1864 822
rect 1892 820 1894 822
rect 1922 820 1924 822
rect 1952 820 1954 822
rect 1982 820 1984 822
rect 3242 818 3244 820
rect 3272 818 3274 820
rect 3302 818 3304 820
rect 3332 818 3334 820
rect 3362 818 3364 820
rect 3636 818 3638 820
rect 3666 818 3668 820
rect 3696 818 3698 820
rect 3726 818 3728 820
rect 3756 818 3758 820
rect 3842 818 3844 820
rect 3872 818 3874 820
rect 3902 818 3904 820
rect 3932 818 3934 820
rect 3962 818 3964 820
rect 4236 818 4238 820
rect 4266 818 4268 820
rect 4296 818 4298 820
rect 4326 818 4328 820
rect 4356 818 4358 820
rect 4442 818 4444 820
rect 4472 818 4474 820
rect 4502 818 4504 820
rect 4532 818 4534 820
rect 4562 818 4564 820
rect 4592 818 4594 820
rect 4622 818 4624 820
rect 4694 818 4696 820
rect 4724 818 4726 820
rect 4776 818 4778 820
rect 4806 818 4808 820
rect 4836 818 4838 820
rect 4866 818 4868 820
rect 4896 818 4898 820
rect 4926 818 4928 820
rect 4956 818 4958 820
rect 5042 818 5044 820
rect 5072 818 5074 820
rect 5102 818 5104 820
rect 5132 818 5134 820
rect 5162 818 5164 820
rect 5192 818 5194 820
rect 5222 818 5224 820
rect 5294 818 5296 820
rect 5324 818 5326 820
rect 5376 818 5378 820
rect 5406 818 5408 820
rect 5436 818 5438 820
rect 5466 818 5468 820
rect 5496 818 5498 820
rect 5526 818 5528 820
rect 5556 818 5558 820
rect 5642 818 5644 820
rect 5672 818 5674 820
rect 5702 818 5704 820
rect 5732 818 5734 820
rect 5762 818 5764 820
rect 6036 818 6038 820
rect 6066 818 6068 820
rect 6096 818 6098 820
rect 6126 818 6128 820
rect 6156 818 6158 820
rect 6242 818 6244 820
rect 6272 818 6274 820
rect 6302 818 6304 820
rect 6332 818 6334 820
rect 6362 818 6364 820
rect 6392 818 6394 820
rect 6422 818 6424 820
rect 6576 818 6578 820
rect 6606 818 6608 820
rect 6636 818 6638 820
rect 6666 818 6668 820
rect 6696 818 6698 820
rect 6726 818 6728 820
rect 6756 818 6758 820
rect 3234 816 3236 818
rect 3240 816 3242 818
rect 3264 816 3266 818
rect 3270 816 3272 818
rect 3294 816 3296 818
rect 3300 816 3302 818
rect 3324 816 3326 818
rect 3330 816 3332 818
rect 3354 816 3356 818
rect 3360 816 3362 818
rect 3384 816 3386 818
rect 3614 816 3616 818
rect 3638 816 3640 818
rect 3644 816 3646 818
rect 3668 816 3670 818
rect 3674 816 3676 818
rect 3698 816 3700 818
rect 3704 816 3706 818
rect 3728 816 3730 818
rect 3734 816 3736 818
rect 3758 816 3760 818
rect 3764 816 3766 818
rect 3834 816 3836 818
rect 3840 816 3842 818
rect 3864 816 3866 818
rect 3870 816 3872 818
rect 3894 816 3896 818
rect 3900 816 3902 818
rect 3924 816 3926 818
rect 3930 816 3932 818
rect 3954 816 3956 818
rect 3960 816 3962 818
rect 3984 816 3986 818
rect 4214 816 4216 818
rect 4238 816 4240 818
rect 4244 816 4246 818
rect 4268 816 4270 818
rect 4274 816 4276 818
rect 4298 816 4300 818
rect 4304 816 4306 818
rect 4328 816 4330 818
rect 4334 816 4336 818
rect 4358 816 4360 818
rect 4364 816 4366 818
rect 4434 816 4436 818
rect 4440 816 4442 818
rect 4464 816 4466 818
rect 4470 816 4472 818
rect 4494 816 4496 818
rect 4500 816 4502 818
rect 4524 816 4526 818
rect 4530 816 4532 818
rect 4554 816 4556 818
rect 4560 816 4562 818
rect 4584 816 4586 818
rect 4590 816 4592 818
rect 4614 816 4616 818
rect 4620 816 4622 818
rect 4686 816 4688 818
rect 4692 816 4694 818
rect 4716 816 4718 818
rect 4722 816 4724 818
rect 4778 816 4780 818
rect 4784 816 4786 818
rect 4808 816 4810 818
rect 4814 816 4816 818
rect 4838 816 4840 818
rect 4844 816 4846 818
rect 4868 816 4870 818
rect 4874 816 4876 818
rect 4898 816 4900 818
rect 4904 816 4906 818
rect 4928 816 4930 818
rect 4934 816 4936 818
rect 4958 816 4960 818
rect 4964 816 4966 818
rect 5034 816 5036 818
rect 5040 816 5042 818
rect 5064 816 5066 818
rect 5070 816 5072 818
rect 5094 816 5096 818
rect 5100 816 5102 818
rect 5124 816 5126 818
rect 5130 816 5132 818
rect 5154 816 5156 818
rect 5160 816 5162 818
rect 5184 816 5186 818
rect 5190 816 5192 818
rect 5214 816 5216 818
rect 5220 816 5222 818
rect 5286 816 5288 818
rect 5292 816 5294 818
rect 5316 816 5318 818
rect 5322 816 5324 818
rect 5378 816 5380 818
rect 5384 816 5386 818
rect 5408 816 5410 818
rect 5414 816 5416 818
rect 5438 816 5440 818
rect 5444 816 5446 818
rect 5468 816 5470 818
rect 5474 816 5476 818
rect 5498 816 5500 818
rect 5504 816 5506 818
rect 5528 816 5530 818
rect 5534 816 5536 818
rect 5558 816 5560 818
rect 5564 816 5566 818
rect 5634 816 5636 818
rect 5640 816 5642 818
rect 5664 816 5666 818
rect 5670 816 5672 818
rect 5694 816 5696 818
rect 5700 816 5702 818
rect 5724 816 5726 818
rect 5730 816 5732 818
rect 5754 816 5756 818
rect 5760 816 5762 818
rect 6038 816 6040 818
rect 6044 816 6046 818
rect 6068 816 6070 818
rect 6074 816 6076 818
rect 6098 816 6100 818
rect 6104 816 6106 818
rect 6128 816 6130 818
rect 6134 816 6136 818
rect 6158 816 6160 818
rect 6164 816 6166 818
rect 6234 816 6236 818
rect 6240 816 6242 818
rect 6264 816 6266 818
rect 6270 816 6272 818
rect 6294 816 6296 818
rect 6300 816 6302 818
rect 6324 816 6326 818
rect 6330 816 6332 818
rect 6354 816 6356 818
rect 6360 816 6362 818
rect 6384 816 6386 818
rect 6390 816 6392 818
rect 6414 816 6416 818
rect 6420 816 6422 818
rect 6578 816 6580 818
rect 6584 816 6586 818
rect 6608 816 6610 818
rect 6614 816 6616 818
rect 6638 816 6640 818
rect 6644 816 6646 818
rect 6668 816 6670 818
rect 6674 816 6676 818
rect 6698 816 6700 818
rect 6704 816 6706 818
rect 6728 816 6730 818
rect 6734 816 6736 818
rect 6758 816 6760 818
rect 6764 816 6766 818
rect 1632 814 1634 816
rect 1692 814 1694 816
rect 1702 814 1704 816
rect 1742 814 1744 816
rect 1772 814 1774 816
rect 1802 814 1804 816
rect 1832 814 1834 816
rect 1862 814 1864 816
rect 1892 814 1894 816
rect 1922 814 1924 816
rect 1952 814 1954 816
rect 1982 814 1984 816
rect 3232 814 3234 816
rect 3262 814 3264 816
rect 3292 814 3294 816
rect 3322 814 3324 816
rect 3352 814 3354 816
rect 3382 814 3384 816
rect 3616 814 3618 816
rect 3646 814 3648 816
rect 3676 814 3678 816
rect 3706 814 3708 816
rect 3736 814 3738 816
rect 3766 814 3768 816
rect 3832 814 3834 816
rect 3862 814 3864 816
rect 3892 814 3894 816
rect 3922 814 3924 816
rect 3952 814 3954 816
rect 3982 814 3984 816
rect 4216 814 4218 816
rect 4246 814 4248 816
rect 4276 814 4278 816
rect 4306 814 4308 816
rect 4336 814 4338 816
rect 4366 814 4368 816
rect 4432 814 4434 816
rect 4462 814 4464 816
rect 4492 814 4494 816
rect 4522 814 4524 816
rect 4552 814 4554 816
rect 4582 814 4584 816
rect 4612 814 4614 816
rect 4684 814 4686 816
rect 4714 814 4716 816
rect 4786 814 4788 816
rect 4816 814 4818 816
rect 4846 814 4848 816
rect 4876 814 4878 816
rect 4906 814 4908 816
rect 4936 814 4938 816
rect 4966 814 4968 816
rect 5032 814 5034 816
rect 5062 814 5064 816
rect 5092 814 5094 816
rect 5122 814 5124 816
rect 5152 814 5154 816
rect 5182 814 5184 816
rect 5212 814 5214 816
rect 5284 814 5286 816
rect 5314 814 5316 816
rect 5386 814 5388 816
rect 5416 814 5418 816
rect 5446 814 5448 816
rect 5476 814 5478 816
rect 5506 814 5508 816
rect 5536 814 5538 816
rect 5566 814 5568 816
rect 5632 814 5634 816
rect 5662 814 5664 816
rect 5692 814 5694 816
rect 5722 814 5724 816
rect 5752 814 5754 816
rect 6046 814 6048 816
rect 6076 814 6078 816
rect 6106 814 6108 816
rect 6136 814 6138 816
rect 6166 814 6168 816
rect 6232 814 6234 816
rect 6262 814 6264 816
rect 6292 814 6294 816
rect 6322 814 6324 816
rect 6352 814 6354 816
rect 6382 814 6384 816
rect 6412 814 6414 816
rect 6586 814 6588 816
rect 6616 814 6618 816
rect 6646 814 6648 816
rect 6676 814 6678 816
rect 6706 814 6708 816
rect 6736 814 6738 816
rect 6766 814 6768 816
rect 1630 812 1632 814
rect 1684 812 1686 814
rect 1690 812 1692 814
rect 1704 812 1706 814
rect 1720 812 1722 814
rect 1744 812 1746 814
rect 1750 812 1752 814
rect 1774 812 1776 814
rect 1780 812 1782 814
rect 1804 812 1806 814
rect 1810 812 1812 814
rect 1834 812 1836 814
rect 1840 812 1842 814
rect 1864 812 1866 814
rect 1870 812 1872 814
rect 1894 812 1896 814
rect 1900 812 1902 814
rect 1924 812 1926 814
rect 1930 812 1932 814
rect 1954 812 1956 814
rect 1960 812 1962 814
rect 1984 812 1986 814
rect 1682 810 1684 812
rect 1722 810 1724 812
rect 1752 810 1754 812
rect 1782 810 1784 812
rect 1812 810 1814 812
rect 1842 810 1844 812
rect 1872 810 1874 812
rect 1902 810 1904 812
rect 1932 810 1934 812
rect 1962 810 1964 812
rect 3232 808 3234 810
rect 3262 808 3264 810
rect 3292 808 3294 810
rect 3322 808 3324 810
rect 3352 808 3354 810
rect 3382 808 3384 810
rect 3616 808 3618 810
rect 3646 808 3648 810
rect 3676 808 3678 810
rect 3706 808 3708 810
rect 3736 808 3738 810
rect 3766 808 3768 810
rect 3832 808 3834 810
rect 3862 808 3864 810
rect 3892 808 3894 810
rect 3922 808 3924 810
rect 3952 808 3954 810
rect 3982 808 3984 810
rect 4216 808 4218 810
rect 4246 808 4248 810
rect 4276 808 4278 810
rect 4306 808 4308 810
rect 4336 808 4338 810
rect 4366 808 4368 810
rect 4432 808 4434 810
rect 4462 808 4464 810
rect 4492 808 4494 810
rect 4522 808 4524 810
rect 4552 808 4554 810
rect 4582 808 4584 810
rect 4612 808 4614 810
rect 4684 808 4686 810
rect 4714 808 4716 810
rect 4786 808 4788 810
rect 4816 808 4818 810
rect 4846 808 4848 810
rect 4876 808 4878 810
rect 4906 808 4908 810
rect 4936 808 4938 810
rect 4966 808 4968 810
rect 5032 808 5034 810
rect 5062 808 5064 810
rect 5092 808 5094 810
rect 5122 808 5124 810
rect 5152 808 5154 810
rect 5182 808 5184 810
rect 5212 808 5214 810
rect 5284 808 5286 810
rect 5314 808 5316 810
rect 5386 808 5388 810
rect 5416 808 5418 810
rect 5446 808 5448 810
rect 5476 808 5478 810
rect 5506 808 5508 810
rect 5536 808 5538 810
rect 5566 808 5568 810
rect 5632 808 5634 810
rect 5662 808 5664 810
rect 5692 808 5694 810
rect 5722 808 5724 810
rect 5752 808 5754 810
rect 6046 808 6048 810
rect 6076 808 6078 810
rect 6106 808 6108 810
rect 6136 808 6138 810
rect 6166 808 6168 810
rect 6232 808 6234 810
rect 6262 808 6264 810
rect 6292 808 6294 810
rect 6322 808 6324 810
rect 6352 808 6354 810
rect 6382 808 6384 810
rect 6412 808 6414 810
rect 6586 808 6588 810
rect 6616 808 6618 810
rect 6646 808 6648 810
rect 6676 808 6678 810
rect 6706 808 6708 810
rect 6736 808 6738 810
rect 6766 808 6768 810
rect 3234 806 3236 808
rect 3240 806 3242 808
rect 3264 806 3266 808
rect 3270 806 3272 808
rect 3294 806 3296 808
rect 3300 806 3302 808
rect 3324 806 3326 808
rect 3330 806 3332 808
rect 3354 806 3356 808
rect 3360 806 3362 808
rect 3384 806 3386 808
rect 3614 806 3616 808
rect 3638 806 3640 808
rect 3644 806 3646 808
rect 3668 806 3670 808
rect 3674 806 3676 808
rect 3698 806 3700 808
rect 3704 806 3706 808
rect 3728 806 3730 808
rect 3734 806 3736 808
rect 3758 806 3760 808
rect 3764 806 3766 808
rect 3834 806 3836 808
rect 3840 806 3842 808
rect 3864 806 3866 808
rect 3870 806 3872 808
rect 3894 806 3896 808
rect 3900 806 3902 808
rect 3924 806 3926 808
rect 3930 806 3932 808
rect 3954 806 3956 808
rect 3960 806 3962 808
rect 3984 806 3986 808
rect 4214 806 4216 808
rect 4238 806 4240 808
rect 4244 806 4246 808
rect 4268 806 4270 808
rect 4274 806 4276 808
rect 4298 806 4300 808
rect 4304 806 4306 808
rect 4328 806 4330 808
rect 4334 806 4336 808
rect 4358 806 4360 808
rect 4364 806 4366 808
rect 4434 806 4436 808
rect 4440 806 4442 808
rect 4464 806 4466 808
rect 4470 806 4472 808
rect 4494 806 4496 808
rect 4500 806 4502 808
rect 4524 806 4526 808
rect 4530 806 4532 808
rect 4554 806 4556 808
rect 4560 806 4562 808
rect 4584 806 4586 808
rect 4590 806 4592 808
rect 4614 806 4616 808
rect 4620 806 4622 808
rect 4686 806 4688 808
rect 4692 806 4694 808
rect 4716 806 4718 808
rect 4722 806 4724 808
rect 4778 806 4780 808
rect 4784 806 4786 808
rect 4808 806 4810 808
rect 4814 806 4816 808
rect 4838 806 4840 808
rect 4844 806 4846 808
rect 4868 806 4870 808
rect 4874 806 4876 808
rect 4898 806 4900 808
rect 4904 806 4906 808
rect 4928 806 4930 808
rect 4934 806 4936 808
rect 4958 806 4960 808
rect 4964 806 4966 808
rect 5034 806 5036 808
rect 5040 806 5042 808
rect 5064 806 5066 808
rect 5070 806 5072 808
rect 5094 806 5096 808
rect 5100 806 5102 808
rect 5124 806 5126 808
rect 5130 806 5132 808
rect 5154 806 5156 808
rect 5160 806 5162 808
rect 5184 806 5186 808
rect 5190 806 5192 808
rect 5214 806 5216 808
rect 5220 806 5222 808
rect 5286 806 5288 808
rect 5292 806 5294 808
rect 5316 806 5318 808
rect 5322 806 5324 808
rect 5378 806 5380 808
rect 5384 806 5386 808
rect 5408 806 5410 808
rect 5414 806 5416 808
rect 5438 806 5440 808
rect 5444 806 5446 808
rect 5468 806 5470 808
rect 5474 806 5476 808
rect 5498 806 5500 808
rect 5504 806 5506 808
rect 5528 806 5530 808
rect 5534 806 5536 808
rect 5558 806 5560 808
rect 5564 806 5566 808
rect 5634 806 5636 808
rect 5640 806 5642 808
rect 5664 806 5666 808
rect 5670 806 5672 808
rect 5694 806 5696 808
rect 5700 806 5702 808
rect 5724 806 5726 808
rect 5730 806 5732 808
rect 5754 806 5756 808
rect 5760 806 5762 808
rect 6038 806 6040 808
rect 6044 806 6046 808
rect 6068 806 6070 808
rect 6074 806 6076 808
rect 6098 806 6100 808
rect 6104 806 6106 808
rect 6128 806 6130 808
rect 6134 806 6136 808
rect 6158 806 6160 808
rect 6164 806 6166 808
rect 6234 806 6236 808
rect 6240 806 6242 808
rect 6264 806 6266 808
rect 6270 806 6272 808
rect 6294 806 6296 808
rect 6300 806 6302 808
rect 6324 806 6326 808
rect 6330 806 6332 808
rect 6354 806 6356 808
rect 6360 806 6362 808
rect 6384 806 6386 808
rect 6390 806 6392 808
rect 6414 806 6416 808
rect 6420 806 6422 808
rect 6578 806 6580 808
rect 6584 806 6586 808
rect 6608 806 6610 808
rect 6614 806 6616 808
rect 6638 806 6640 808
rect 6644 806 6646 808
rect 6668 806 6670 808
rect 6674 806 6676 808
rect 6698 806 6700 808
rect 6704 806 6706 808
rect 6728 806 6730 808
rect 6734 806 6736 808
rect 6758 806 6760 808
rect 6764 806 6766 808
rect 1622 804 1624 806
rect 1682 804 1684 806
rect 1722 804 1724 806
rect 1752 804 1754 806
rect 1782 804 1784 806
rect 1812 804 1814 806
rect 1842 804 1844 806
rect 1872 804 1874 806
rect 1902 804 1904 806
rect 1932 804 1934 806
rect 1962 804 1964 806
rect 3242 804 3244 806
rect 3272 804 3274 806
rect 3302 804 3304 806
rect 3332 804 3334 806
rect 3362 804 3364 806
rect 3636 804 3638 806
rect 3666 804 3668 806
rect 3696 804 3698 806
rect 3726 804 3728 806
rect 3756 804 3758 806
rect 3842 804 3844 806
rect 3872 804 3874 806
rect 3902 804 3904 806
rect 3932 804 3934 806
rect 3962 804 3964 806
rect 4236 804 4238 806
rect 4266 804 4268 806
rect 4296 804 4298 806
rect 4326 804 4328 806
rect 4356 804 4358 806
rect 4442 804 4444 806
rect 4472 804 4474 806
rect 4502 804 4504 806
rect 4532 804 4534 806
rect 4562 804 4564 806
rect 4592 804 4594 806
rect 4622 804 4624 806
rect 4694 804 4696 806
rect 4724 804 4726 806
rect 4776 804 4778 806
rect 4806 804 4808 806
rect 4836 804 4838 806
rect 4866 804 4868 806
rect 4896 804 4898 806
rect 4926 804 4928 806
rect 4956 804 4958 806
rect 5042 804 5044 806
rect 5072 804 5074 806
rect 5102 804 5104 806
rect 5132 804 5134 806
rect 5162 804 5164 806
rect 5192 804 5194 806
rect 5222 804 5224 806
rect 5294 804 5296 806
rect 5324 804 5326 806
rect 5376 804 5378 806
rect 5406 804 5408 806
rect 5436 804 5438 806
rect 5466 804 5468 806
rect 5496 804 5498 806
rect 5526 804 5528 806
rect 5556 804 5558 806
rect 5642 804 5644 806
rect 5672 804 5674 806
rect 5702 804 5704 806
rect 5732 804 5734 806
rect 5762 804 5764 806
rect 6036 804 6038 806
rect 6066 804 6068 806
rect 6096 804 6098 806
rect 6126 804 6128 806
rect 6156 804 6158 806
rect 6242 804 6244 806
rect 6272 804 6274 806
rect 6302 804 6304 806
rect 6332 804 6334 806
rect 6362 804 6364 806
rect 6392 804 6394 806
rect 6422 804 6424 806
rect 6576 804 6578 806
rect 6606 804 6608 806
rect 6636 804 6638 806
rect 6666 804 6668 806
rect 6696 804 6698 806
rect 6726 804 6728 806
rect 6756 804 6758 806
rect 1620 802 1622 804
rect 1674 802 1676 804
rect 1680 802 1682 804
rect 1704 802 1706 804
rect 1720 802 1722 804
rect 1744 802 1746 804
rect 1750 802 1752 804
rect 1774 802 1776 804
rect 1780 802 1782 804
rect 1804 802 1806 804
rect 1810 802 1812 804
rect 1834 802 1836 804
rect 1840 802 1842 804
rect 1864 802 1866 804
rect 1870 802 1872 804
rect 1894 802 1896 804
rect 1900 802 1902 804
rect 1924 802 1926 804
rect 1930 802 1932 804
rect 1954 802 1956 804
rect 1960 802 1962 804
rect 1984 802 1986 804
rect 1672 800 1674 802
rect 1702 800 1704 802
rect 1742 800 1744 802
rect 1772 800 1774 802
rect 1802 800 1804 802
rect 1832 800 1834 802
rect 1862 800 1864 802
rect 1892 800 1894 802
rect 1922 800 1924 802
rect 1952 800 1954 802
rect 1982 800 1984 802
rect 3242 798 3244 800
rect 3272 798 3274 800
rect 3302 798 3304 800
rect 3332 798 3334 800
rect 3362 798 3364 800
rect 3636 798 3638 800
rect 3666 798 3668 800
rect 3696 798 3698 800
rect 3726 798 3728 800
rect 3756 798 3758 800
rect 3842 798 3844 800
rect 3872 798 3874 800
rect 3902 798 3904 800
rect 3932 798 3934 800
rect 3962 798 3964 800
rect 4236 798 4238 800
rect 4266 798 4268 800
rect 4296 798 4298 800
rect 4326 798 4328 800
rect 4356 798 4358 800
rect 4442 798 4444 800
rect 4472 798 4474 800
rect 4502 798 4504 800
rect 4532 798 4534 800
rect 4562 798 4564 800
rect 4592 798 4594 800
rect 4622 798 4624 800
rect 4694 798 4696 800
rect 4724 798 4726 800
rect 4776 798 4778 800
rect 4806 798 4808 800
rect 4836 798 4838 800
rect 4866 798 4868 800
rect 4896 798 4898 800
rect 4926 798 4928 800
rect 4956 798 4958 800
rect 5042 798 5044 800
rect 5072 798 5074 800
rect 5102 798 5104 800
rect 5132 798 5134 800
rect 5162 798 5164 800
rect 5192 798 5194 800
rect 5222 798 5224 800
rect 5294 798 5296 800
rect 5324 798 5326 800
rect 5376 798 5378 800
rect 5406 798 5408 800
rect 5436 798 5438 800
rect 5466 798 5468 800
rect 5496 798 5498 800
rect 5526 798 5528 800
rect 5556 798 5558 800
rect 5642 798 5644 800
rect 5672 798 5674 800
rect 5702 798 5704 800
rect 5732 798 5734 800
rect 5762 798 5764 800
rect 6036 798 6038 800
rect 6066 798 6068 800
rect 6096 798 6098 800
rect 6126 798 6128 800
rect 6156 798 6158 800
rect 6242 798 6244 800
rect 6272 798 6274 800
rect 6302 798 6304 800
rect 6332 798 6334 800
rect 6362 798 6364 800
rect 6392 798 6394 800
rect 6422 798 6424 800
rect 6576 798 6578 800
rect 6606 798 6608 800
rect 6636 798 6638 800
rect 6666 798 6668 800
rect 6696 798 6698 800
rect 6726 798 6728 800
rect 6756 798 6758 800
rect 3234 796 3236 798
rect 3240 796 3242 798
rect 3264 796 3266 798
rect 3270 796 3272 798
rect 3294 796 3296 798
rect 3300 796 3302 798
rect 3324 796 3326 798
rect 3330 796 3332 798
rect 3354 796 3356 798
rect 3360 796 3362 798
rect 3384 796 3386 798
rect 3614 796 3616 798
rect 3638 796 3640 798
rect 3644 796 3646 798
rect 3668 796 3670 798
rect 3674 796 3676 798
rect 3698 796 3700 798
rect 3704 796 3706 798
rect 3728 796 3730 798
rect 3734 796 3736 798
rect 3758 796 3760 798
rect 3764 796 3766 798
rect 3834 796 3836 798
rect 3840 796 3842 798
rect 3864 796 3866 798
rect 3870 796 3872 798
rect 3894 796 3896 798
rect 3900 796 3902 798
rect 3924 796 3926 798
rect 3930 796 3932 798
rect 3954 796 3956 798
rect 3960 796 3962 798
rect 3984 796 3986 798
rect 4214 796 4216 798
rect 4238 796 4240 798
rect 4244 796 4246 798
rect 4268 796 4270 798
rect 4274 796 4276 798
rect 4298 796 4300 798
rect 4304 796 4306 798
rect 4328 796 4330 798
rect 4334 796 4336 798
rect 4358 796 4360 798
rect 4364 796 4366 798
rect 4434 796 4436 798
rect 4440 796 4442 798
rect 4464 796 4466 798
rect 4470 796 4472 798
rect 4494 796 4496 798
rect 4500 796 4502 798
rect 4524 796 4526 798
rect 4530 796 4532 798
rect 4554 796 4556 798
rect 4560 796 4562 798
rect 4584 796 4586 798
rect 4590 796 4592 798
rect 4614 796 4616 798
rect 4620 796 4622 798
rect 4686 796 4688 798
rect 4692 796 4694 798
rect 4716 796 4718 798
rect 4722 796 4724 798
rect 4778 796 4780 798
rect 4784 796 4786 798
rect 4808 796 4810 798
rect 4814 796 4816 798
rect 4838 796 4840 798
rect 4844 796 4846 798
rect 4868 796 4870 798
rect 4874 796 4876 798
rect 4898 796 4900 798
rect 4904 796 4906 798
rect 4928 796 4930 798
rect 4934 796 4936 798
rect 4958 796 4960 798
rect 4964 796 4966 798
rect 5034 796 5036 798
rect 5040 796 5042 798
rect 5064 796 5066 798
rect 5070 796 5072 798
rect 5094 796 5096 798
rect 5100 796 5102 798
rect 5124 796 5126 798
rect 5130 796 5132 798
rect 5154 796 5156 798
rect 5160 796 5162 798
rect 5184 796 5186 798
rect 5190 796 5192 798
rect 5214 796 5216 798
rect 5220 796 5222 798
rect 5286 796 5288 798
rect 5292 796 5294 798
rect 5316 796 5318 798
rect 5322 796 5324 798
rect 5378 796 5380 798
rect 5384 796 5386 798
rect 5408 796 5410 798
rect 5414 796 5416 798
rect 5438 796 5440 798
rect 5444 796 5446 798
rect 5468 796 5470 798
rect 5474 796 5476 798
rect 5498 796 5500 798
rect 5504 796 5506 798
rect 5528 796 5530 798
rect 5534 796 5536 798
rect 5558 796 5560 798
rect 5564 796 5566 798
rect 5634 796 5636 798
rect 5640 796 5642 798
rect 5664 796 5666 798
rect 5670 796 5672 798
rect 5694 796 5696 798
rect 5700 796 5702 798
rect 5724 796 5726 798
rect 5730 796 5732 798
rect 5754 796 5756 798
rect 5760 796 5762 798
rect 6038 796 6040 798
rect 6044 796 6046 798
rect 6068 796 6070 798
rect 6074 796 6076 798
rect 6098 796 6100 798
rect 6104 796 6106 798
rect 6128 796 6130 798
rect 6134 796 6136 798
rect 6158 796 6160 798
rect 6164 796 6166 798
rect 6234 796 6236 798
rect 6240 796 6242 798
rect 6264 796 6266 798
rect 6270 796 6272 798
rect 6294 796 6296 798
rect 6300 796 6302 798
rect 6324 796 6326 798
rect 6330 796 6332 798
rect 6354 796 6356 798
rect 6360 796 6362 798
rect 6384 796 6386 798
rect 6390 796 6392 798
rect 6414 796 6416 798
rect 6420 796 6422 798
rect 6578 796 6580 798
rect 6584 796 6586 798
rect 6608 796 6610 798
rect 6614 796 6616 798
rect 6638 796 6640 798
rect 6644 796 6646 798
rect 6668 796 6670 798
rect 6674 796 6676 798
rect 6698 796 6700 798
rect 6704 796 6706 798
rect 6728 796 6730 798
rect 6734 796 6736 798
rect 6758 796 6760 798
rect 6764 796 6766 798
rect 1612 794 1614 796
rect 1672 794 1674 796
rect 1702 794 1704 796
rect 1742 794 1744 796
rect 1772 794 1774 796
rect 1802 794 1804 796
rect 1832 794 1834 796
rect 1862 794 1864 796
rect 1892 794 1894 796
rect 1922 794 1924 796
rect 1952 794 1954 796
rect 1982 794 1984 796
rect 3232 794 3234 796
rect 3262 794 3264 796
rect 3292 794 3294 796
rect 3322 794 3324 796
rect 3352 794 3354 796
rect 3382 794 3384 796
rect 3616 794 3618 796
rect 3646 794 3648 796
rect 3676 794 3678 796
rect 3706 794 3708 796
rect 3736 794 3738 796
rect 3766 794 3768 796
rect 3832 794 3834 796
rect 3862 794 3864 796
rect 3892 794 3894 796
rect 3922 794 3924 796
rect 3952 794 3954 796
rect 3982 794 3984 796
rect 4216 794 4218 796
rect 4246 794 4248 796
rect 4276 794 4278 796
rect 4306 794 4308 796
rect 4336 794 4338 796
rect 4366 794 4368 796
rect 4432 794 4434 796
rect 4462 794 4464 796
rect 4492 794 4494 796
rect 4522 794 4524 796
rect 4552 794 4554 796
rect 4582 794 4584 796
rect 4612 794 4614 796
rect 4684 794 4686 796
rect 4714 794 4716 796
rect 4786 794 4788 796
rect 4816 794 4818 796
rect 4846 794 4848 796
rect 4876 794 4878 796
rect 4906 794 4908 796
rect 4936 794 4938 796
rect 4966 794 4968 796
rect 5032 794 5034 796
rect 5062 794 5064 796
rect 5092 794 5094 796
rect 5122 794 5124 796
rect 5152 794 5154 796
rect 5182 794 5184 796
rect 5212 794 5214 796
rect 5284 794 5286 796
rect 5314 794 5316 796
rect 5386 794 5388 796
rect 5416 794 5418 796
rect 5446 794 5448 796
rect 5476 794 5478 796
rect 5506 794 5508 796
rect 5536 794 5538 796
rect 5566 794 5568 796
rect 5632 794 5634 796
rect 5662 794 5664 796
rect 5692 794 5694 796
rect 5722 794 5724 796
rect 5752 794 5754 796
rect 6046 794 6048 796
rect 6076 794 6078 796
rect 6106 794 6108 796
rect 6136 794 6138 796
rect 6166 794 6168 796
rect 6232 794 6234 796
rect 6262 794 6264 796
rect 6292 794 6294 796
rect 6322 794 6324 796
rect 6352 794 6354 796
rect 6382 794 6384 796
rect 6412 794 6414 796
rect 6586 794 6588 796
rect 6616 794 6618 796
rect 6646 794 6648 796
rect 6676 794 6678 796
rect 6706 794 6708 796
rect 6736 794 6738 796
rect 6766 794 6768 796
rect 1610 792 1612 794
rect 1664 792 1666 794
rect 1670 792 1672 794
rect 1704 792 1706 794
rect 1720 792 1722 794
rect 1744 792 1746 794
rect 1750 792 1752 794
rect 1774 792 1776 794
rect 1780 792 1782 794
rect 1804 792 1806 794
rect 1810 792 1812 794
rect 1834 792 1836 794
rect 1840 792 1842 794
rect 1864 792 1866 794
rect 1870 792 1872 794
rect 1894 792 1896 794
rect 1900 792 1902 794
rect 1924 792 1926 794
rect 1930 792 1932 794
rect 1954 792 1956 794
rect 1960 792 1962 794
rect 1984 792 1986 794
rect 1662 790 1664 792
rect 1722 790 1724 792
rect 1752 790 1754 792
rect 1782 790 1784 792
rect 1812 790 1814 792
rect 1842 790 1844 792
rect 1872 790 1874 792
rect 1902 790 1904 792
rect 1932 790 1934 792
rect 1962 790 1964 792
rect 3232 788 3234 790
rect 3262 788 3264 790
rect 3292 788 3294 790
rect 3322 788 3324 790
rect 3352 788 3354 790
rect 3382 788 3384 790
rect 3616 788 3618 790
rect 3646 788 3648 790
rect 3676 788 3678 790
rect 3706 788 3708 790
rect 3736 788 3738 790
rect 3766 788 3768 790
rect 3832 788 3834 790
rect 3862 788 3864 790
rect 3892 788 3894 790
rect 3922 788 3924 790
rect 3952 788 3954 790
rect 3982 788 3984 790
rect 4216 788 4218 790
rect 4246 788 4248 790
rect 4276 788 4278 790
rect 4306 788 4308 790
rect 4336 788 4338 790
rect 4366 788 4368 790
rect 4432 788 4434 790
rect 4462 788 4464 790
rect 4492 788 4494 790
rect 4522 788 4524 790
rect 4552 788 4554 790
rect 4582 788 4584 790
rect 4612 788 4614 790
rect 4684 788 4686 790
rect 4714 788 4716 790
rect 4786 788 4788 790
rect 4816 788 4818 790
rect 4846 788 4848 790
rect 4876 788 4878 790
rect 4906 788 4908 790
rect 4936 788 4938 790
rect 4966 788 4968 790
rect 5032 788 5034 790
rect 5062 788 5064 790
rect 5092 788 5094 790
rect 5122 788 5124 790
rect 5152 788 5154 790
rect 5182 788 5184 790
rect 5212 788 5214 790
rect 5284 788 5286 790
rect 5314 788 5316 790
rect 5386 788 5388 790
rect 5416 788 5418 790
rect 5446 788 5448 790
rect 5476 788 5478 790
rect 5506 788 5508 790
rect 5536 788 5538 790
rect 5566 788 5568 790
rect 5632 788 5634 790
rect 5662 788 5664 790
rect 5692 788 5694 790
rect 5722 788 5724 790
rect 5752 788 5754 790
rect 6046 788 6048 790
rect 6076 788 6078 790
rect 6106 788 6108 790
rect 6136 788 6138 790
rect 6166 788 6168 790
rect 6232 788 6234 790
rect 6262 788 6264 790
rect 6292 788 6294 790
rect 6322 788 6324 790
rect 6352 788 6354 790
rect 6382 788 6384 790
rect 6412 788 6414 790
rect 6586 788 6588 790
rect 6616 788 6618 790
rect 6646 788 6648 790
rect 6676 788 6678 790
rect 6706 788 6708 790
rect 6736 788 6738 790
rect 6766 788 6768 790
rect 3234 786 3236 788
rect 3240 786 3242 788
rect 3264 786 3266 788
rect 3270 786 3272 788
rect 3294 786 3296 788
rect 3300 786 3302 788
rect 3324 786 3326 788
rect 3330 786 3332 788
rect 3354 786 3356 788
rect 3360 786 3362 788
rect 3384 786 3386 788
rect 3614 786 3616 788
rect 3638 786 3640 788
rect 3644 786 3646 788
rect 3668 786 3670 788
rect 3674 786 3676 788
rect 3698 786 3700 788
rect 3704 786 3706 788
rect 3728 786 3730 788
rect 3734 786 3736 788
rect 3758 786 3760 788
rect 3764 786 3766 788
rect 3834 786 3836 788
rect 3840 786 3842 788
rect 3864 786 3866 788
rect 3870 786 3872 788
rect 3894 786 3896 788
rect 3900 786 3902 788
rect 3924 786 3926 788
rect 3930 786 3932 788
rect 3954 786 3956 788
rect 3960 786 3962 788
rect 3984 786 3986 788
rect 4214 786 4216 788
rect 4238 786 4240 788
rect 4244 786 4246 788
rect 4268 786 4270 788
rect 4274 786 4276 788
rect 4298 786 4300 788
rect 4304 786 4306 788
rect 4328 786 4330 788
rect 4334 786 4336 788
rect 4358 786 4360 788
rect 4364 786 4366 788
rect 4434 786 4436 788
rect 4440 786 4442 788
rect 4464 786 4466 788
rect 4470 786 4472 788
rect 4494 786 4496 788
rect 4500 786 4502 788
rect 4524 786 4526 788
rect 4530 786 4532 788
rect 4554 786 4556 788
rect 4560 786 4562 788
rect 4584 786 4586 788
rect 4590 786 4592 788
rect 4614 786 4616 788
rect 4620 786 4622 788
rect 4686 786 4688 788
rect 4692 786 4694 788
rect 4716 786 4718 788
rect 4722 786 4724 788
rect 4778 786 4780 788
rect 4784 786 4786 788
rect 4808 786 4810 788
rect 4814 786 4816 788
rect 4838 786 4840 788
rect 4844 786 4846 788
rect 4868 786 4870 788
rect 4874 786 4876 788
rect 4898 786 4900 788
rect 4904 786 4906 788
rect 4928 786 4930 788
rect 4934 786 4936 788
rect 4958 786 4960 788
rect 4964 786 4966 788
rect 5034 786 5036 788
rect 5040 786 5042 788
rect 5064 786 5066 788
rect 5070 786 5072 788
rect 5094 786 5096 788
rect 5100 786 5102 788
rect 5124 786 5126 788
rect 5130 786 5132 788
rect 5154 786 5156 788
rect 5160 786 5162 788
rect 5184 786 5186 788
rect 5190 786 5192 788
rect 5214 786 5216 788
rect 5220 786 5222 788
rect 5286 786 5288 788
rect 5292 786 5294 788
rect 5316 786 5318 788
rect 5322 786 5324 788
rect 5378 786 5380 788
rect 5384 786 5386 788
rect 5408 786 5410 788
rect 5414 786 5416 788
rect 5438 786 5440 788
rect 5444 786 5446 788
rect 5468 786 5470 788
rect 5474 786 5476 788
rect 5498 786 5500 788
rect 5504 786 5506 788
rect 5528 786 5530 788
rect 5534 786 5536 788
rect 5558 786 5560 788
rect 5564 786 5566 788
rect 5634 786 5636 788
rect 5640 786 5642 788
rect 5664 786 5666 788
rect 5670 786 5672 788
rect 5694 786 5696 788
rect 5700 786 5702 788
rect 5724 786 5726 788
rect 5730 786 5732 788
rect 5754 786 5756 788
rect 5760 786 5762 788
rect 6038 786 6040 788
rect 6044 786 6046 788
rect 6068 786 6070 788
rect 6074 786 6076 788
rect 6098 786 6100 788
rect 6104 786 6106 788
rect 6128 786 6130 788
rect 6134 786 6136 788
rect 6158 786 6160 788
rect 6164 786 6166 788
rect 6234 786 6236 788
rect 6240 786 6242 788
rect 6264 786 6266 788
rect 6270 786 6272 788
rect 6294 786 6296 788
rect 6300 786 6302 788
rect 6324 786 6326 788
rect 6330 786 6332 788
rect 6354 786 6356 788
rect 6360 786 6362 788
rect 6384 786 6386 788
rect 6390 786 6392 788
rect 6414 786 6416 788
rect 6420 786 6422 788
rect 6578 786 6580 788
rect 6584 786 6586 788
rect 6608 786 6610 788
rect 6614 786 6616 788
rect 6638 786 6640 788
rect 6644 786 6646 788
rect 6668 786 6670 788
rect 6674 786 6676 788
rect 6698 786 6700 788
rect 6704 786 6706 788
rect 6728 786 6730 788
rect 6734 786 6736 788
rect 6758 786 6760 788
rect 6764 786 6766 788
rect 1602 784 1604 786
rect 1662 784 1664 786
rect 1722 784 1724 786
rect 1752 784 1754 786
rect 1782 784 1784 786
rect 1812 784 1814 786
rect 1842 784 1844 786
rect 1872 784 1874 786
rect 1902 784 1904 786
rect 1932 784 1934 786
rect 1962 784 1964 786
rect 3242 784 3244 786
rect 3272 784 3274 786
rect 3302 784 3304 786
rect 3332 784 3334 786
rect 3362 784 3364 786
rect 3636 784 3638 786
rect 3666 784 3668 786
rect 3696 784 3698 786
rect 3726 784 3728 786
rect 3756 784 3758 786
rect 3842 784 3844 786
rect 3872 784 3874 786
rect 3902 784 3904 786
rect 3932 784 3934 786
rect 3962 784 3964 786
rect 4236 784 4238 786
rect 4266 784 4268 786
rect 4296 784 4298 786
rect 4326 784 4328 786
rect 4356 784 4358 786
rect 4442 784 4444 786
rect 4472 784 4474 786
rect 4502 784 4504 786
rect 4532 784 4534 786
rect 4562 784 4564 786
rect 4592 784 4594 786
rect 4622 784 4624 786
rect 4694 784 4696 786
rect 4724 784 4726 786
rect 4776 784 4778 786
rect 4806 784 4808 786
rect 4836 784 4838 786
rect 4866 784 4868 786
rect 4896 784 4898 786
rect 4926 784 4928 786
rect 4956 784 4958 786
rect 5042 784 5044 786
rect 5072 784 5074 786
rect 5102 784 5104 786
rect 5132 784 5134 786
rect 5162 784 5164 786
rect 5192 784 5194 786
rect 5222 784 5224 786
rect 5294 784 5296 786
rect 5324 784 5326 786
rect 5376 784 5378 786
rect 5406 784 5408 786
rect 5436 784 5438 786
rect 5466 784 5468 786
rect 5496 784 5498 786
rect 5526 784 5528 786
rect 5556 784 5558 786
rect 5642 784 5644 786
rect 5672 784 5674 786
rect 5702 784 5704 786
rect 5732 784 5734 786
rect 5762 784 5764 786
rect 6036 784 6038 786
rect 6066 784 6068 786
rect 6096 784 6098 786
rect 6126 784 6128 786
rect 6156 784 6158 786
rect 6242 784 6244 786
rect 6272 784 6274 786
rect 6302 784 6304 786
rect 6332 784 6334 786
rect 6362 784 6364 786
rect 6392 784 6394 786
rect 6422 784 6424 786
rect 6576 784 6578 786
rect 6606 784 6608 786
rect 6636 784 6638 786
rect 6666 784 6668 786
rect 6696 784 6698 786
rect 6726 784 6728 786
rect 6756 784 6758 786
rect 1600 782 1602 784
rect 1654 782 1656 784
rect 1660 782 1662 784
rect 1704 782 1706 784
rect 1720 782 1722 784
rect 1744 782 1746 784
rect 1750 782 1752 784
rect 1774 782 1776 784
rect 1780 782 1782 784
rect 1804 782 1806 784
rect 1810 782 1812 784
rect 1834 782 1836 784
rect 1840 782 1842 784
rect 1864 782 1866 784
rect 1870 782 1872 784
rect 1894 782 1896 784
rect 1900 782 1902 784
rect 1924 782 1926 784
rect 1930 782 1932 784
rect 1954 782 1956 784
rect 1960 782 1962 784
rect 1984 782 1986 784
rect 1652 780 1654 782
rect 1702 780 1704 782
rect 1742 780 1744 782
rect 1772 780 1774 782
rect 1802 780 1804 782
rect 1832 780 1834 782
rect 1862 780 1864 782
rect 1892 780 1894 782
rect 1922 780 1924 782
rect 1952 780 1954 782
rect 1982 780 1984 782
rect 2404 781 2415 782
rect 3004 781 3015 782
rect 3242 778 3244 780
rect 3272 778 3274 780
rect 3726 778 3728 780
rect 3756 778 3758 780
rect 3842 778 3844 780
rect 3872 778 3874 780
rect 4326 778 4328 780
rect 4356 778 4358 780
rect 4442 778 4444 780
rect 4472 778 4474 780
rect 4926 778 4928 780
rect 4956 778 4958 780
rect 5042 778 5044 780
rect 5072 778 5074 780
rect 5526 778 5528 780
rect 5556 778 5558 780
rect 5642 778 5644 780
rect 5672 778 5674 780
rect 6126 778 6128 780
rect 6156 778 6158 780
rect 6242 778 6244 780
rect 6272 778 6274 780
rect 6726 778 6728 780
rect 6756 778 6758 780
rect 3234 776 3236 778
rect 3240 776 3242 778
rect 3264 776 3266 778
rect 3270 776 3272 778
rect 3294 776 3296 778
rect 3310 776 3312 778
rect 3324 776 3326 778
rect 3340 776 3342 778
rect 3354 776 3356 778
rect 3370 776 3372 778
rect 3384 776 3386 778
rect 3614 776 3616 778
rect 3628 776 3630 778
rect 3644 776 3646 778
rect 3658 776 3660 778
rect 3674 776 3676 778
rect 3688 776 3690 778
rect 3704 776 3706 778
rect 3728 776 3730 778
rect 3734 776 3736 778
rect 3758 776 3760 778
rect 3764 776 3766 778
rect 3834 776 3836 778
rect 3840 776 3842 778
rect 3864 776 3866 778
rect 3870 776 3872 778
rect 3894 776 3896 778
rect 3910 776 3912 778
rect 3924 776 3926 778
rect 3940 776 3942 778
rect 3954 776 3956 778
rect 3970 776 3972 778
rect 3984 776 3986 778
rect 4214 776 4216 778
rect 4228 776 4230 778
rect 4244 776 4246 778
rect 4258 776 4260 778
rect 4274 776 4276 778
rect 4288 776 4290 778
rect 4304 776 4306 778
rect 4328 776 4330 778
rect 4334 776 4336 778
rect 4358 776 4360 778
rect 4364 776 4366 778
rect 4434 776 4436 778
rect 4440 776 4442 778
rect 4464 776 4466 778
rect 4470 776 4472 778
rect 4494 776 4496 778
rect 4510 776 4512 778
rect 4524 776 4526 778
rect 4540 776 4542 778
rect 4554 776 4556 778
rect 4570 776 4572 778
rect 4584 776 4586 778
rect 4600 776 4602 778
rect 4614 776 4616 778
rect 4630 776 4632 778
rect 4644 776 4646 778
rect 4666 776 4668 778
rect 4672 776 4674 778
rect 4686 776 4688 778
rect 4702 776 4704 778
rect 4716 776 4718 778
rect 4732 776 4734 778
rect 4754 776 4756 778
rect 4768 776 4770 778
rect 4784 776 4786 778
rect 4798 776 4800 778
rect 4814 776 4816 778
rect 4828 776 4830 778
rect 4844 776 4846 778
rect 4858 776 4860 778
rect 4874 776 4876 778
rect 4888 776 4890 778
rect 4904 776 4906 778
rect 4928 776 4930 778
rect 4934 776 4936 778
rect 4958 776 4960 778
rect 4964 776 4966 778
rect 5034 776 5036 778
rect 5040 776 5042 778
rect 5064 776 5066 778
rect 5070 776 5072 778
rect 5094 776 5096 778
rect 5110 776 5112 778
rect 5124 776 5126 778
rect 5140 776 5142 778
rect 5154 776 5156 778
rect 5170 776 5172 778
rect 5184 776 5186 778
rect 5200 776 5202 778
rect 5214 776 5216 778
rect 5230 776 5232 778
rect 5244 776 5246 778
rect 5266 776 5268 778
rect 5272 776 5274 778
rect 5286 776 5288 778
rect 5302 776 5304 778
rect 5316 776 5318 778
rect 5332 776 5334 778
rect 5354 776 5356 778
rect 5368 776 5370 778
rect 5384 776 5386 778
rect 5398 776 5400 778
rect 5414 776 5416 778
rect 5428 776 5430 778
rect 5444 776 5446 778
rect 5458 776 5460 778
rect 5474 776 5476 778
rect 5488 776 5490 778
rect 5504 776 5506 778
rect 5528 776 5530 778
rect 5534 776 5536 778
rect 5558 776 5560 778
rect 5564 776 5566 778
rect 5634 776 5636 778
rect 5640 776 5642 778
rect 5664 776 5666 778
rect 5670 776 5672 778
rect 5694 776 5696 778
rect 5710 776 5712 778
rect 5724 776 5726 778
rect 5740 776 5742 778
rect 5754 776 5756 778
rect 5770 776 5772 778
rect 5784 776 5786 778
rect 5892 776 5894 778
rect 5906 776 5908 778
rect 6014 776 6016 778
rect 6028 776 6030 778
rect 6044 776 6046 778
rect 6058 776 6060 778
rect 6074 776 6076 778
rect 6088 776 6090 778
rect 6104 776 6106 778
rect 6128 776 6130 778
rect 6134 776 6136 778
rect 6158 776 6160 778
rect 6164 776 6166 778
rect 6234 776 6236 778
rect 6240 776 6242 778
rect 6264 776 6266 778
rect 6270 776 6272 778
rect 6294 776 6296 778
rect 6310 776 6312 778
rect 6324 776 6326 778
rect 6340 776 6342 778
rect 6354 776 6356 778
rect 6370 776 6372 778
rect 6384 776 6386 778
rect 6400 776 6402 778
rect 6414 776 6416 778
rect 6430 776 6432 778
rect 6444 776 6446 778
rect 6460 776 6462 778
rect 6474 776 6476 778
rect 6480 776 6482 778
rect 6518 776 6520 778
rect 6524 776 6526 778
rect 6538 776 6540 778
rect 6554 776 6556 778
rect 6568 776 6570 778
rect 6584 776 6586 778
rect 6598 776 6600 778
rect 6614 776 6616 778
rect 6628 776 6630 778
rect 6644 776 6646 778
rect 6658 776 6660 778
rect 6674 776 6676 778
rect 6688 776 6690 778
rect 6704 776 6706 778
rect 6728 776 6730 778
rect 6734 776 6736 778
rect 6758 776 6760 778
rect 6764 776 6766 778
rect 1652 774 1654 776
rect 1742 774 1744 776
rect 1772 774 1774 776
rect 1802 774 1804 776
rect 1832 774 1834 776
rect 1862 774 1864 776
rect 1892 774 1894 776
rect 1922 774 1924 776
rect 1952 774 1954 776
rect 1982 774 1984 776
rect 3232 774 3234 776
rect 3262 774 3264 776
rect 3292 774 3294 776
rect 3312 774 3314 776
rect 3322 774 3324 776
rect 3342 774 3344 776
rect 3352 774 3354 776
rect 3372 774 3374 776
rect 3382 774 3384 776
rect 3616 774 3618 776
rect 3626 774 3628 776
rect 3646 774 3648 776
rect 3656 774 3658 776
rect 3676 774 3678 776
rect 3686 774 3688 776
rect 3706 774 3708 776
rect 3736 774 3738 776
rect 3766 774 3768 776
rect 3832 774 3834 776
rect 3862 774 3864 776
rect 3892 774 3894 776
rect 3912 774 3914 776
rect 3922 774 3924 776
rect 3942 774 3944 776
rect 3952 774 3954 776
rect 3972 774 3974 776
rect 3982 774 3984 776
rect 4216 774 4218 776
rect 4226 774 4228 776
rect 4246 774 4248 776
rect 4256 774 4258 776
rect 4276 774 4278 776
rect 4286 774 4288 776
rect 4306 774 4308 776
rect 4336 774 4338 776
rect 4366 774 4368 776
rect 4432 774 4434 776
rect 4462 774 4464 776
rect 4492 774 4494 776
rect 4512 774 4514 776
rect 4522 774 4524 776
rect 4542 774 4544 776
rect 4552 774 4554 776
rect 4572 774 4574 776
rect 4582 774 4584 776
rect 4602 774 4604 776
rect 4612 774 4614 776
rect 4632 774 4634 776
rect 4642 774 4644 776
rect 4664 774 4666 776
rect 4674 774 4676 776
rect 4684 774 4686 776
rect 4704 774 4706 776
rect 4714 774 4716 776
rect 4734 774 4736 776
rect 4756 774 4758 776
rect 4766 774 4768 776
rect 4786 774 4788 776
rect 4796 774 4798 776
rect 4816 774 4818 776
rect 4826 774 4828 776
rect 4846 774 4848 776
rect 4856 774 4858 776
rect 4876 774 4878 776
rect 4886 774 4888 776
rect 4906 774 4908 776
rect 4936 774 4938 776
rect 4966 774 4968 776
rect 5032 774 5034 776
rect 5062 774 5064 776
rect 5092 774 5094 776
rect 5112 774 5114 776
rect 5122 774 5124 776
rect 5142 774 5144 776
rect 5152 774 5154 776
rect 5172 774 5174 776
rect 5182 774 5184 776
rect 5202 774 5204 776
rect 5212 774 5214 776
rect 5232 774 5234 776
rect 5242 774 5244 776
rect 5264 774 5266 776
rect 5274 774 5276 776
rect 5284 774 5286 776
rect 5304 774 5306 776
rect 5314 774 5316 776
rect 5334 774 5336 776
rect 5356 774 5358 776
rect 5366 774 5368 776
rect 5386 774 5388 776
rect 5396 774 5398 776
rect 5416 774 5418 776
rect 5426 774 5428 776
rect 5446 774 5448 776
rect 5456 774 5458 776
rect 5476 774 5478 776
rect 5486 774 5488 776
rect 5506 774 5508 776
rect 5536 774 5538 776
rect 5566 774 5568 776
rect 5632 774 5634 776
rect 5662 774 5664 776
rect 5692 774 5694 776
rect 5712 774 5714 776
rect 5722 774 5724 776
rect 5742 774 5744 776
rect 5752 774 5754 776
rect 5772 774 5774 776
rect 5782 774 5784 776
rect 5894 774 5896 776
rect 5904 774 5906 776
rect 6016 774 6018 776
rect 6026 774 6028 776
rect 6046 774 6048 776
rect 6056 774 6058 776
rect 6076 774 6078 776
rect 6086 774 6088 776
rect 6106 774 6108 776
rect 6136 774 6138 776
rect 6166 774 6168 776
rect 6232 774 6234 776
rect 6262 774 6264 776
rect 6292 774 6294 776
rect 6312 774 6314 776
rect 6322 774 6324 776
rect 6342 774 6344 776
rect 6352 774 6354 776
rect 6372 774 6374 776
rect 6382 774 6384 776
rect 6402 774 6404 776
rect 6412 774 6414 776
rect 6432 774 6434 776
rect 6442 774 6444 776
rect 6462 774 6464 776
rect 6472 774 6474 776
rect 6482 774 6484 776
rect 6516 774 6518 776
rect 6526 774 6528 776
rect 6536 774 6538 776
rect 6556 774 6558 776
rect 6566 774 6568 776
rect 6586 774 6588 776
rect 6596 774 6598 776
rect 6616 774 6618 776
rect 6626 774 6628 776
rect 6646 774 6648 776
rect 6656 774 6658 776
rect 6676 774 6678 776
rect 6686 774 6688 776
rect 6706 774 6708 776
rect 6736 774 6738 776
rect 6766 774 6768 776
rect 1644 772 1646 774
rect 1650 772 1652 774
rect 1694 772 1696 774
rect 1720 772 1722 774
rect 1744 772 1746 774
rect 1750 772 1752 774
rect 1774 772 1776 774
rect 1780 772 1782 774
rect 1804 772 1806 774
rect 1810 772 1812 774
rect 1834 772 1836 774
rect 1840 772 1842 774
rect 1864 772 1866 774
rect 1870 772 1872 774
rect 1894 772 1896 774
rect 1900 772 1902 774
rect 1924 772 1926 774
rect 1930 772 1932 774
rect 1954 772 1956 774
rect 1960 772 1962 774
rect 1984 772 1986 774
rect 1642 770 1644 772
rect 1692 770 1694 772
rect 1722 770 1724 772
rect 1752 770 1754 772
rect 1782 770 1784 772
rect 1812 770 1814 772
rect 1842 770 1844 772
rect 1872 770 1874 772
rect 1902 770 1904 772
rect 1932 770 1934 772
rect 1962 770 1964 772
rect 3232 768 3234 770
rect 3262 768 3264 770
rect 3292 768 3294 770
rect 3312 768 3314 770
rect 3322 768 3324 770
rect 3342 768 3344 770
rect 3352 768 3354 770
rect 3372 768 3374 770
rect 3382 768 3384 770
rect 3616 768 3618 770
rect 3626 768 3628 770
rect 3646 768 3648 770
rect 3656 768 3658 770
rect 3676 768 3678 770
rect 3686 768 3688 770
rect 3706 768 3708 770
rect 3736 768 3738 770
rect 3766 768 3768 770
rect 3832 768 3834 770
rect 3862 768 3864 770
rect 3892 768 3894 770
rect 3912 768 3914 770
rect 3922 768 3924 770
rect 3942 768 3944 770
rect 3952 768 3954 770
rect 3972 768 3974 770
rect 3982 768 3984 770
rect 4216 768 4218 770
rect 4226 768 4228 770
rect 4246 768 4248 770
rect 4256 768 4258 770
rect 4276 768 4278 770
rect 4286 768 4288 770
rect 4306 768 4308 770
rect 4336 768 4338 770
rect 4366 768 4368 770
rect 4432 768 4434 770
rect 4462 768 4464 770
rect 4492 768 4494 770
rect 4512 768 4514 770
rect 4522 768 4524 770
rect 4542 768 4544 770
rect 4552 768 4554 770
rect 4572 768 4574 770
rect 4582 768 4584 770
rect 4602 768 4604 770
rect 4612 768 4614 770
rect 4632 768 4634 770
rect 4642 768 4644 770
rect 4664 768 4666 770
rect 4674 768 4676 770
rect 4684 768 4686 770
rect 4704 768 4706 770
rect 4714 768 4716 770
rect 4734 768 4736 770
rect 4756 768 4758 770
rect 4766 768 4768 770
rect 4786 768 4788 770
rect 4796 768 4798 770
rect 4816 768 4818 770
rect 4826 768 4828 770
rect 4846 768 4848 770
rect 4856 768 4858 770
rect 4876 768 4878 770
rect 4886 768 4888 770
rect 4906 768 4908 770
rect 4936 768 4938 770
rect 4966 768 4968 770
rect 5032 768 5034 770
rect 5062 768 5064 770
rect 5092 768 5094 770
rect 5112 768 5114 770
rect 5122 768 5124 770
rect 5142 768 5144 770
rect 5152 768 5154 770
rect 5172 768 5174 770
rect 5182 768 5184 770
rect 5202 768 5204 770
rect 5212 768 5214 770
rect 5232 768 5234 770
rect 5242 768 5244 770
rect 5264 768 5266 770
rect 5274 768 5276 770
rect 5284 768 5286 770
rect 5304 768 5306 770
rect 5314 768 5316 770
rect 5334 768 5336 770
rect 5356 768 5358 770
rect 5366 768 5368 770
rect 5386 768 5388 770
rect 5396 768 5398 770
rect 5416 768 5418 770
rect 5426 768 5428 770
rect 5446 768 5448 770
rect 5456 768 5458 770
rect 5476 768 5478 770
rect 5486 768 5488 770
rect 5506 768 5508 770
rect 5536 768 5538 770
rect 5566 768 5568 770
rect 5632 768 5634 770
rect 5662 768 5664 770
rect 5692 768 5694 770
rect 5712 768 5714 770
rect 5722 768 5724 770
rect 5742 768 5744 770
rect 5752 768 5754 770
rect 5772 768 5774 770
rect 5782 768 5784 770
rect 5894 768 5896 770
rect 5904 768 5906 770
rect 6016 768 6018 770
rect 6026 768 6028 770
rect 6046 768 6048 770
rect 6056 768 6058 770
rect 6076 768 6078 770
rect 6086 768 6088 770
rect 6106 768 6108 770
rect 6136 768 6138 770
rect 6166 768 6168 770
rect 6232 768 6234 770
rect 6262 768 6264 770
rect 6292 768 6294 770
rect 6312 768 6314 770
rect 6322 768 6324 770
rect 6342 768 6344 770
rect 6352 768 6354 770
rect 6372 768 6374 770
rect 6382 768 6384 770
rect 6402 768 6404 770
rect 6412 768 6414 770
rect 6432 768 6434 770
rect 6442 768 6444 770
rect 6462 768 6464 770
rect 6472 768 6474 770
rect 6482 768 6484 770
rect 6516 768 6518 770
rect 6526 768 6528 770
rect 6536 768 6538 770
rect 6556 768 6558 770
rect 6566 768 6568 770
rect 6586 768 6588 770
rect 6596 768 6598 770
rect 6616 768 6618 770
rect 6626 768 6628 770
rect 6646 768 6648 770
rect 6656 768 6658 770
rect 6676 768 6678 770
rect 6686 768 6688 770
rect 6706 768 6708 770
rect 6736 768 6738 770
rect 6766 768 6768 770
rect 3234 766 3236 768
rect 3240 766 3242 768
rect 3264 766 3266 768
rect 3270 766 3272 768
rect 3294 766 3296 768
rect 3310 766 3312 768
rect 3324 766 3326 768
rect 3340 766 3342 768
rect 3354 766 3356 768
rect 3370 766 3372 768
rect 3384 766 3386 768
rect 3614 766 3616 768
rect 3628 766 3630 768
rect 3644 766 3646 768
rect 3658 766 3660 768
rect 3674 766 3676 768
rect 3688 766 3690 768
rect 3704 766 3706 768
rect 3728 766 3730 768
rect 3734 766 3736 768
rect 3758 766 3760 768
rect 3764 766 3766 768
rect 3834 766 3836 768
rect 3840 766 3842 768
rect 3864 766 3866 768
rect 3870 766 3872 768
rect 3894 766 3896 768
rect 3910 766 3912 768
rect 3924 766 3926 768
rect 3940 766 3942 768
rect 3954 766 3956 768
rect 3970 766 3972 768
rect 3984 766 3986 768
rect 4214 766 4216 768
rect 4228 766 4230 768
rect 4244 766 4246 768
rect 4258 766 4260 768
rect 4274 766 4276 768
rect 4288 766 4290 768
rect 4304 766 4306 768
rect 4328 766 4330 768
rect 4334 766 4336 768
rect 4358 766 4360 768
rect 4364 766 4366 768
rect 4434 766 4436 768
rect 4440 766 4442 768
rect 4464 766 4466 768
rect 4470 766 4472 768
rect 4494 766 4496 768
rect 4510 766 4512 768
rect 4524 766 4526 768
rect 4540 766 4542 768
rect 4554 766 4556 768
rect 4570 766 4572 768
rect 4584 766 4586 768
rect 4600 766 4602 768
rect 4614 766 4616 768
rect 4630 766 4632 768
rect 4644 766 4646 768
rect 4666 766 4668 768
rect 4672 766 4674 768
rect 4686 766 4688 768
rect 4702 766 4704 768
rect 4716 766 4718 768
rect 4732 766 4734 768
rect 4754 766 4756 768
rect 4768 766 4770 768
rect 4784 766 4786 768
rect 4798 766 4800 768
rect 4814 766 4816 768
rect 4828 766 4830 768
rect 4844 766 4846 768
rect 4858 766 4860 768
rect 4874 766 4876 768
rect 4888 766 4890 768
rect 4904 766 4906 768
rect 4928 766 4930 768
rect 4934 766 4936 768
rect 4958 766 4960 768
rect 4964 766 4966 768
rect 5034 766 5036 768
rect 5040 766 5042 768
rect 5064 766 5066 768
rect 5070 766 5072 768
rect 5094 766 5096 768
rect 5110 766 5112 768
rect 5124 766 5126 768
rect 5140 766 5142 768
rect 5154 766 5156 768
rect 5170 766 5172 768
rect 5184 766 5186 768
rect 5200 766 5202 768
rect 5214 766 5216 768
rect 5230 766 5232 768
rect 5244 766 5246 768
rect 5266 766 5268 768
rect 5272 766 5274 768
rect 5286 766 5288 768
rect 5302 766 5304 768
rect 5316 766 5318 768
rect 5332 766 5334 768
rect 5354 766 5356 768
rect 5368 766 5370 768
rect 5384 766 5386 768
rect 5398 766 5400 768
rect 5414 766 5416 768
rect 5428 766 5430 768
rect 5444 766 5446 768
rect 5458 766 5460 768
rect 5474 766 5476 768
rect 5488 766 5490 768
rect 5504 766 5506 768
rect 5528 766 5530 768
rect 5534 766 5536 768
rect 5558 766 5560 768
rect 5564 766 5566 768
rect 5634 766 5636 768
rect 5640 766 5642 768
rect 5664 766 5666 768
rect 5670 766 5672 768
rect 5694 766 5696 768
rect 5710 766 5712 768
rect 5724 766 5726 768
rect 5740 766 5742 768
rect 5754 766 5756 768
rect 5770 766 5772 768
rect 5784 766 5786 768
rect 5896 766 5898 768
rect 5902 766 5904 768
rect 6014 766 6016 768
rect 6028 766 6030 768
rect 6044 766 6046 768
rect 6058 766 6060 768
rect 6074 766 6076 768
rect 6088 766 6090 768
rect 6104 766 6106 768
rect 6128 766 6130 768
rect 6134 766 6136 768
rect 6158 766 6160 768
rect 6164 766 6166 768
rect 6234 766 6236 768
rect 6240 766 6242 768
rect 6264 766 6266 768
rect 6270 766 6272 768
rect 6294 766 6296 768
rect 6310 766 6312 768
rect 6324 766 6326 768
rect 6340 766 6342 768
rect 6354 766 6356 768
rect 6370 766 6372 768
rect 6384 766 6386 768
rect 6400 766 6402 768
rect 6414 766 6416 768
rect 6430 766 6432 768
rect 6444 766 6446 768
rect 6460 766 6462 768
rect 6474 766 6476 768
rect 6480 766 6482 768
rect 6518 766 6520 768
rect 6524 766 6526 768
rect 6538 766 6540 768
rect 6554 766 6556 768
rect 6568 766 6570 768
rect 6584 766 6586 768
rect 6598 766 6600 768
rect 6614 766 6616 768
rect 6628 766 6630 768
rect 6644 766 6646 768
rect 6658 766 6660 768
rect 6674 766 6676 768
rect 6688 766 6690 768
rect 6704 766 6706 768
rect 6728 766 6730 768
rect 6734 766 6736 768
rect 6758 766 6760 768
rect 6764 766 6766 768
rect 1642 764 1644 766
rect 1692 764 1694 766
rect 1702 764 1704 766
rect 1722 764 1724 766
rect 1752 764 1754 766
rect 1782 764 1784 766
rect 1812 764 1814 766
rect 1842 764 1844 766
rect 1872 764 1874 766
rect 1902 764 1904 766
rect 1932 764 1934 766
rect 1962 764 1964 766
rect 3242 764 3244 766
rect 3272 764 3274 766
rect 3726 764 3728 766
rect 3756 764 3758 766
rect 3842 764 3844 766
rect 3872 764 3874 766
rect 4326 764 4328 766
rect 4356 764 4358 766
rect 4442 764 4444 766
rect 4472 764 4474 766
rect 4926 764 4928 766
rect 4956 764 4958 766
rect 5042 764 5044 766
rect 5072 764 5074 766
rect 5526 764 5528 766
rect 5556 764 5558 766
rect 5642 764 5644 766
rect 5672 764 5674 766
rect 6126 764 6128 766
rect 6156 764 6158 766
rect 6242 764 6244 766
rect 6272 764 6274 766
rect 6726 764 6728 766
rect 6756 764 6758 766
rect 1634 762 1636 764
rect 1640 762 1642 764
rect 1684 762 1686 764
rect 1690 762 1692 764
rect 1704 762 1706 764
rect 1720 762 1722 764
rect 1744 762 1746 764
rect 1750 762 1752 764
rect 1774 762 1776 764
rect 1780 762 1782 764
rect 1804 762 1806 764
rect 1810 762 1812 764
rect 1834 762 1836 764
rect 1840 762 1842 764
rect 1864 762 1866 764
rect 1870 762 1872 764
rect 1894 762 1896 764
rect 1900 762 1902 764
rect 1924 762 1926 764
rect 1930 762 1932 764
rect 1954 762 1956 764
rect 1960 762 1962 764
rect 1984 762 1986 764
rect 1632 760 1634 762
rect 1682 760 1684 762
rect 1742 760 1744 762
rect 1772 760 1774 762
rect 1802 760 1804 762
rect 1832 760 1834 762
rect 1862 760 1864 762
rect 1892 760 1894 762
rect 1922 760 1924 762
rect 1952 760 1954 762
rect 1982 760 1984 762
rect 3242 758 3244 760
rect 3272 758 3274 760
rect 3302 758 3304 760
rect 3332 758 3334 760
rect 3362 758 3364 760
rect 3636 758 3638 760
rect 3666 758 3668 760
rect 3696 758 3698 760
rect 3726 758 3728 760
rect 3756 758 3758 760
rect 3842 758 3844 760
rect 3872 758 3874 760
rect 3902 758 3904 760
rect 3932 758 3934 760
rect 3962 758 3964 760
rect 4236 758 4238 760
rect 4266 758 4268 760
rect 4296 758 4298 760
rect 4326 758 4328 760
rect 4356 758 4358 760
rect 4442 758 4444 760
rect 4472 758 4474 760
rect 4502 758 4504 760
rect 4532 758 4534 760
rect 4562 758 4564 760
rect 4592 758 4594 760
rect 4622 758 4624 760
rect 4694 758 4696 760
rect 4724 758 4726 760
rect 4776 758 4778 760
rect 4806 758 4808 760
rect 4836 758 4838 760
rect 4866 758 4868 760
rect 4896 758 4898 760
rect 4926 758 4928 760
rect 4956 758 4958 760
rect 5042 758 5044 760
rect 5072 758 5074 760
rect 5102 758 5104 760
rect 5132 758 5134 760
rect 5162 758 5164 760
rect 5192 758 5194 760
rect 5222 758 5224 760
rect 5294 758 5296 760
rect 5324 758 5326 760
rect 5376 758 5378 760
rect 5406 758 5408 760
rect 5436 758 5438 760
rect 5466 758 5468 760
rect 5496 758 5498 760
rect 5526 758 5528 760
rect 5556 758 5558 760
rect 5642 758 5644 760
rect 5672 758 5674 760
rect 5702 758 5704 760
rect 5732 758 5734 760
rect 5762 758 5764 760
rect 6036 758 6038 760
rect 6066 758 6068 760
rect 6096 758 6098 760
rect 6126 758 6128 760
rect 6156 758 6158 760
rect 6242 758 6244 760
rect 6272 758 6274 760
rect 6302 758 6304 760
rect 6332 758 6334 760
rect 6362 758 6364 760
rect 6392 758 6394 760
rect 6422 758 6424 760
rect 6576 758 6578 760
rect 6606 758 6608 760
rect 6636 758 6638 760
rect 6666 758 6668 760
rect 6696 758 6698 760
rect 6726 758 6728 760
rect 6756 758 6758 760
rect 3234 756 3236 758
rect 3240 756 3242 758
rect 3264 756 3266 758
rect 3270 756 3272 758
rect 3294 756 3296 758
rect 3300 756 3302 758
rect 3324 756 3326 758
rect 3330 756 3332 758
rect 3354 756 3356 758
rect 3360 756 3362 758
rect 3384 756 3386 758
rect 3614 756 3616 758
rect 3638 756 3640 758
rect 3644 756 3646 758
rect 3668 756 3670 758
rect 3674 756 3676 758
rect 3698 756 3700 758
rect 3704 756 3706 758
rect 3728 756 3730 758
rect 3734 756 3736 758
rect 3758 756 3760 758
rect 3764 756 3766 758
rect 3834 756 3836 758
rect 3840 756 3842 758
rect 3864 756 3866 758
rect 3870 756 3872 758
rect 3894 756 3896 758
rect 3900 756 3902 758
rect 3924 756 3926 758
rect 3930 756 3932 758
rect 3954 756 3956 758
rect 3960 756 3962 758
rect 3984 756 3986 758
rect 4214 756 4216 758
rect 4238 756 4240 758
rect 4244 756 4246 758
rect 4268 756 4270 758
rect 4274 756 4276 758
rect 4298 756 4300 758
rect 4304 756 4306 758
rect 4328 756 4330 758
rect 4334 756 4336 758
rect 4358 756 4360 758
rect 4364 756 4366 758
rect 4434 756 4436 758
rect 4440 756 4442 758
rect 4464 756 4466 758
rect 4470 756 4472 758
rect 4494 756 4496 758
rect 4500 756 4502 758
rect 4524 756 4526 758
rect 4530 756 4532 758
rect 4554 756 4556 758
rect 4560 756 4562 758
rect 4584 756 4586 758
rect 4590 756 4592 758
rect 4614 756 4616 758
rect 4620 756 4622 758
rect 4686 756 4688 758
rect 4692 756 4694 758
rect 4716 756 4718 758
rect 4722 756 4724 758
rect 4778 756 4780 758
rect 4784 756 4786 758
rect 4808 756 4810 758
rect 4814 756 4816 758
rect 4838 756 4840 758
rect 4844 756 4846 758
rect 4868 756 4870 758
rect 4874 756 4876 758
rect 4898 756 4900 758
rect 4904 756 4906 758
rect 4928 756 4930 758
rect 4934 756 4936 758
rect 4958 756 4960 758
rect 4964 756 4966 758
rect 5034 756 5036 758
rect 5040 756 5042 758
rect 5064 756 5066 758
rect 5070 756 5072 758
rect 5094 756 5096 758
rect 5100 756 5102 758
rect 5124 756 5126 758
rect 5130 756 5132 758
rect 5154 756 5156 758
rect 5160 756 5162 758
rect 5184 756 5186 758
rect 5190 756 5192 758
rect 5214 756 5216 758
rect 5220 756 5222 758
rect 5286 756 5288 758
rect 5292 756 5294 758
rect 5316 756 5318 758
rect 5322 756 5324 758
rect 5378 756 5380 758
rect 5384 756 5386 758
rect 5408 756 5410 758
rect 5414 756 5416 758
rect 5438 756 5440 758
rect 5444 756 5446 758
rect 5468 756 5470 758
rect 5474 756 5476 758
rect 5498 756 5500 758
rect 5504 756 5506 758
rect 5528 756 5530 758
rect 5534 756 5536 758
rect 5558 756 5560 758
rect 5564 756 5566 758
rect 5634 756 5636 758
rect 5640 756 5642 758
rect 5664 756 5666 758
rect 5670 756 5672 758
rect 5694 756 5696 758
rect 5700 756 5702 758
rect 5724 756 5726 758
rect 5730 756 5732 758
rect 5754 756 5756 758
rect 5760 756 5762 758
rect 6038 756 6040 758
rect 6044 756 6046 758
rect 6068 756 6070 758
rect 6074 756 6076 758
rect 6098 756 6100 758
rect 6104 756 6106 758
rect 6128 756 6130 758
rect 6134 756 6136 758
rect 6158 756 6160 758
rect 6164 756 6166 758
rect 6234 756 6236 758
rect 6240 756 6242 758
rect 6264 756 6266 758
rect 6270 756 6272 758
rect 6294 756 6296 758
rect 6300 756 6302 758
rect 6324 756 6326 758
rect 6330 756 6332 758
rect 6354 756 6356 758
rect 6360 756 6362 758
rect 6384 756 6386 758
rect 6390 756 6392 758
rect 6414 756 6416 758
rect 6420 756 6422 758
rect 6578 756 6580 758
rect 6584 756 6586 758
rect 6608 756 6610 758
rect 6614 756 6616 758
rect 6638 756 6640 758
rect 6644 756 6646 758
rect 6668 756 6670 758
rect 6674 756 6676 758
rect 6698 756 6700 758
rect 6704 756 6706 758
rect 6728 756 6730 758
rect 6734 756 6736 758
rect 6758 756 6760 758
rect 6764 756 6766 758
rect 1632 754 1634 756
rect 1682 754 1684 756
rect 1742 754 1744 756
rect 1772 754 1774 756
rect 1802 754 1804 756
rect 1832 754 1834 756
rect 1862 754 1864 756
rect 1892 754 1894 756
rect 1922 754 1924 756
rect 1952 754 1954 756
rect 1982 754 1984 756
rect 3232 754 3234 756
rect 3262 754 3264 756
rect 3292 754 3294 756
rect 3322 754 3324 756
rect 3352 754 3354 756
rect 3382 754 3384 756
rect 3616 754 3618 756
rect 3646 754 3648 756
rect 3676 754 3678 756
rect 3706 754 3708 756
rect 3736 754 3738 756
rect 3766 754 3768 756
rect 3832 754 3834 756
rect 3862 754 3864 756
rect 3892 754 3894 756
rect 3922 754 3924 756
rect 3952 754 3954 756
rect 3982 754 3984 756
rect 4216 754 4218 756
rect 4246 754 4248 756
rect 4276 754 4278 756
rect 4306 754 4308 756
rect 4336 754 4338 756
rect 4366 754 4368 756
rect 4432 754 4434 756
rect 4462 754 4464 756
rect 4492 754 4494 756
rect 4522 754 4524 756
rect 4552 754 4554 756
rect 4582 754 4584 756
rect 4612 754 4614 756
rect 4684 754 4686 756
rect 4714 754 4716 756
rect 4786 754 4788 756
rect 4816 754 4818 756
rect 4846 754 4848 756
rect 4876 754 4878 756
rect 4906 754 4908 756
rect 4936 754 4938 756
rect 4966 754 4968 756
rect 5032 754 5034 756
rect 5062 754 5064 756
rect 5092 754 5094 756
rect 5122 754 5124 756
rect 5152 754 5154 756
rect 5182 754 5184 756
rect 5212 754 5214 756
rect 5284 754 5286 756
rect 5314 754 5316 756
rect 5386 754 5388 756
rect 5416 754 5418 756
rect 5446 754 5448 756
rect 5476 754 5478 756
rect 5506 754 5508 756
rect 5536 754 5538 756
rect 5566 754 5568 756
rect 5632 754 5634 756
rect 5662 754 5664 756
rect 5692 754 5694 756
rect 5722 754 5724 756
rect 5752 754 5754 756
rect 6046 754 6048 756
rect 6076 754 6078 756
rect 6106 754 6108 756
rect 6136 754 6138 756
rect 6166 754 6168 756
rect 6232 754 6234 756
rect 6262 754 6264 756
rect 6292 754 6294 756
rect 6322 754 6324 756
rect 6352 754 6354 756
rect 6382 754 6384 756
rect 6412 754 6414 756
rect 6586 754 6588 756
rect 6616 754 6618 756
rect 6646 754 6648 756
rect 6676 754 6678 756
rect 6706 754 6708 756
rect 6736 754 6738 756
rect 6766 754 6768 756
rect 1624 752 1626 754
rect 1630 752 1632 754
rect 1674 752 1676 754
rect 1680 752 1682 754
rect 1704 752 1706 754
rect 1720 752 1722 754
rect 1744 752 1746 754
rect 1750 752 1752 754
rect 1774 752 1776 754
rect 1780 752 1782 754
rect 1804 752 1806 754
rect 1810 752 1812 754
rect 1834 752 1836 754
rect 1840 752 1842 754
rect 1864 752 1866 754
rect 1870 752 1872 754
rect 1894 752 1896 754
rect 1900 752 1902 754
rect 1924 752 1926 754
rect 1930 752 1932 754
rect 1954 752 1956 754
rect 1960 752 1962 754
rect 1984 752 1986 754
rect 1622 750 1624 752
rect 1672 750 1674 752
rect 1702 750 1704 752
rect 1722 750 1724 752
rect 1752 750 1754 752
rect 1782 750 1784 752
rect 1812 750 1814 752
rect 1842 750 1844 752
rect 1872 750 1874 752
rect 1902 750 1904 752
rect 1932 750 1934 752
rect 1962 750 1964 752
rect 3232 748 3234 750
rect 3262 748 3264 750
rect 3292 748 3294 750
rect 3322 748 3324 750
rect 3352 748 3354 750
rect 3382 748 3384 750
rect 3616 748 3618 750
rect 3646 748 3648 750
rect 3676 748 3678 750
rect 3706 748 3708 750
rect 3736 748 3738 750
rect 3766 748 3768 750
rect 3832 748 3834 750
rect 3862 748 3864 750
rect 3892 748 3894 750
rect 3922 748 3924 750
rect 3952 748 3954 750
rect 3982 748 3984 750
rect 4216 748 4218 750
rect 4246 748 4248 750
rect 4276 748 4278 750
rect 4306 748 4308 750
rect 4336 748 4338 750
rect 4366 748 4368 750
rect 4432 748 4434 750
rect 4462 748 4464 750
rect 4492 748 4494 750
rect 4522 748 4524 750
rect 4552 748 4554 750
rect 4582 748 4584 750
rect 4612 748 4614 750
rect 4684 748 4686 750
rect 4714 748 4716 750
rect 4786 748 4788 750
rect 4816 748 4818 750
rect 4846 748 4848 750
rect 4876 748 4878 750
rect 4906 748 4908 750
rect 4936 748 4938 750
rect 4966 748 4968 750
rect 5032 748 5034 750
rect 5062 748 5064 750
rect 5092 748 5094 750
rect 5122 748 5124 750
rect 5152 748 5154 750
rect 5182 748 5184 750
rect 5212 748 5214 750
rect 5284 748 5286 750
rect 5314 748 5316 750
rect 5386 748 5388 750
rect 5416 748 5418 750
rect 5446 748 5448 750
rect 5476 748 5478 750
rect 5506 748 5508 750
rect 5536 748 5538 750
rect 5566 748 5568 750
rect 5632 748 5634 750
rect 5662 748 5664 750
rect 5692 748 5694 750
rect 5722 748 5724 750
rect 5752 748 5754 750
rect 6046 748 6048 750
rect 6076 748 6078 750
rect 6106 748 6108 750
rect 6136 748 6138 750
rect 6166 748 6168 750
rect 6232 748 6234 750
rect 6262 748 6264 750
rect 6292 748 6294 750
rect 6322 748 6324 750
rect 6352 748 6354 750
rect 6382 748 6384 750
rect 6412 748 6414 750
rect 6586 748 6588 750
rect 6616 748 6618 750
rect 6646 748 6648 750
rect 6676 748 6678 750
rect 6706 748 6708 750
rect 6736 748 6738 750
rect 6766 748 6768 750
rect 3234 746 3236 748
rect 3240 746 3242 748
rect 3264 746 3266 748
rect 3270 746 3272 748
rect 3294 746 3296 748
rect 3300 746 3302 748
rect 3324 746 3326 748
rect 3330 746 3332 748
rect 3354 746 3356 748
rect 3360 746 3362 748
rect 3384 746 3386 748
rect 3614 746 3616 748
rect 3638 746 3640 748
rect 3644 746 3646 748
rect 3668 746 3670 748
rect 3674 746 3676 748
rect 3698 746 3700 748
rect 3704 746 3706 748
rect 3728 746 3730 748
rect 3734 746 3736 748
rect 3758 746 3760 748
rect 3764 746 3766 748
rect 3834 746 3836 748
rect 3840 746 3842 748
rect 3864 746 3866 748
rect 3870 746 3872 748
rect 3894 746 3896 748
rect 3900 746 3902 748
rect 3924 746 3926 748
rect 3930 746 3932 748
rect 3954 746 3956 748
rect 3960 746 3962 748
rect 3984 746 3986 748
rect 4214 746 4216 748
rect 4238 746 4240 748
rect 4244 746 4246 748
rect 4268 746 4270 748
rect 4274 746 4276 748
rect 4298 746 4300 748
rect 4304 746 4306 748
rect 4328 746 4330 748
rect 4334 746 4336 748
rect 4358 746 4360 748
rect 4364 746 4366 748
rect 4434 746 4436 748
rect 4440 746 4442 748
rect 4464 746 4466 748
rect 4470 746 4472 748
rect 4494 746 4496 748
rect 4500 746 4502 748
rect 4524 746 4526 748
rect 4530 746 4532 748
rect 4554 746 4556 748
rect 4560 746 4562 748
rect 4584 746 4586 748
rect 4590 746 4592 748
rect 4614 746 4616 748
rect 4620 746 4622 748
rect 4686 746 4688 748
rect 4692 746 4694 748
rect 4716 746 4718 748
rect 4722 746 4724 748
rect 4778 746 4780 748
rect 4784 746 4786 748
rect 4808 746 4810 748
rect 4814 746 4816 748
rect 4838 746 4840 748
rect 4844 746 4846 748
rect 4868 746 4870 748
rect 4874 746 4876 748
rect 4898 746 4900 748
rect 4904 746 4906 748
rect 4928 746 4930 748
rect 4934 746 4936 748
rect 4958 746 4960 748
rect 4964 746 4966 748
rect 5034 746 5036 748
rect 5040 746 5042 748
rect 5064 746 5066 748
rect 5070 746 5072 748
rect 5094 746 5096 748
rect 5100 746 5102 748
rect 5124 746 5126 748
rect 5130 746 5132 748
rect 5154 746 5156 748
rect 5160 746 5162 748
rect 5184 746 5186 748
rect 5190 746 5192 748
rect 5214 746 5216 748
rect 5220 746 5222 748
rect 5286 746 5288 748
rect 5292 746 5294 748
rect 5316 746 5318 748
rect 5322 746 5324 748
rect 5378 746 5380 748
rect 5384 746 5386 748
rect 5408 746 5410 748
rect 5414 746 5416 748
rect 5438 746 5440 748
rect 5444 746 5446 748
rect 5468 746 5470 748
rect 5474 746 5476 748
rect 5498 746 5500 748
rect 5504 746 5506 748
rect 5528 746 5530 748
rect 5534 746 5536 748
rect 5558 746 5560 748
rect 5564 746 5566 748
rect 5634 746 5636 748
rect 5640 746 5642 748
rect 5664 746 5666 748
rect 5670 746 5672 748
rect 5694 746 5696 748
rect 5700 746 5702 748
rect 5724 746 5726 748
rect 5730 746 5732 748
rect 5754 746 5756 748
rect 5760 746 5762 748
rect 6038 746 6040 748
rect 6044 746 6046 748
rect 6068 746 6070 748
rect 6074 746 6076 748
rect 6098 746 6100 748
rect 6104 746 6106 748
rect 6128 746 6130 748
rect 6134 746 6136 748
rect 6158 746 6160 748
rect 6164 746 6166 748
rect 6234 746 6236 748
rect 6240 746 6242 748
rect 6264 746 6266 748
rect 6270 746 6272 748
rect 6294 746 6296 748
rect 6300 746 6302 748
rect 6324 746 6326 748
rect 6330 746 6332 748
rect 6354 746 6356 748
rect 6360 746 6362 748
rect 6384 746 6386 748
rect 6390 746 6392 748
rect 6414 746 6416 748
rect 6420 746 6422 748
rect 6578 746 6580 748
rect 6584 746 6586 748
rect 6608 746 6610 748
rect 6614 746 6616 748
rect 6638 746 6640 748
rect 6644 746 6646 748
rect 6668 746 6670 748
rect 6674 746 6676 748
rect 6698 746 6700 748
rect 6704 746 6706 748
rect 6728 746 6730 748
rect 6734 746 6736 748
rect 6758 746 6760 748
rect 6764 746 6766 748
rect 1622 744 1624 746
rect 1672 744 1674 746
rect 1722 744 1724 746
rect 1752 744 1754 746
rect 1782 744 1784 746
rect 1812 744 1814 746
rect 1842 744 1844 746
rect 1872 744 1874 746
rect 1902 744 1904 746
rect 1932 744 1934 746
rect 1962 744 1964 746
rect 3242 744 3244 746
rect 3272 744 3274 746
rect 3302 744 3304 746
rect 3332 744 3334 746
rect 3362 744 3364 746
rect 3636 744 3638 746
rect 3666 744 3668 746
rect 3696 744 3698 746
rect 3726 744 3728 746
rect 3756 744 3758 746
rect 3842 744 3844 746
rect 3872 744 3874 746
rect 3902 744 3904 746
rect 3932 744 3934 746
rect 3962 744 3964 746
rect 4236 744 4238 746
rect 4266 744 4268 746
rect 4296 744 4298 746
rect 4326 744 4328 746
rect 4356 744 4358 746
rect 4442 744 4444 746
rect 4472 744 4474 746
rect 4502 744 4504 746
rect 4532 744 4534 746
rect 4562 744 4564 746
rect 4592 744 4594 746
rect 4622 744 4624 746
rect 4694 744 4696 746
rect 4724 744 4726 746
rect 4776 744 4778 746
rect 4806 744 4808 746
rect 4836 744 4838 746
rect 4866 744 4868 746
rect 4896 744 4898 746
rect 4926 744 4928 746
rect 4956 744 4958 746
rect 5042 744 5044 746
rect 5072 744 5074 746
rect 5102 744 5104 746
rect 5132 744 5134 746
rect 5162 744 5164 746
rect 5192 744 5194 746
rect 5222 744 5224 746
rect 5294 744 5296 746
rect 5324 744 5326 746
rect 5376 744 5378 746
rect 5406 744 5408 746
rect 5436 744 5438 746
rect 5466 744 5468 746
rect 5496 744 5498 746
rect 5526 744 5528 746
rect 5556 744 5558 746
rect 5642 744 5644 746
rect 5672 744 5674 746
rect 5702 744 5704 746
rect 5732 744 5734 746
rect 5762 744 5764 746
rect 6036 744 6038 746
rect 6066 744 6068 746
rect 6096 744 6098 746
rect 6126 744 6128 746
rect 6156 744 6158 746
rect 6242 744 6244 746
rect 6272 744 6274 746
rect 6302 744 6304 746
rect 6332 744 6334 746
rect 6362 744 6364 746
rect 6392 744 6394 746
rect 6422 744 6424 746
rect 6576 744 6578 746
rect 6606 744 6608 746
rect 6636 744 6638 746
rect 6666 744 6668 746
rect 6696 744 6698 746
rect 6726 744 6728 746
rect 6756 744 6758 746
rect 1614 742 1616 744
rect 1620 742 1622 744
rect 1664 742 1666 744
rect 1670 742 1672 744
rect 1694 742 1696 744
rect 1720 742 1722 744
rect 1744 742 1746 744
rect 1750 742 1752 744
rect 1774 742 1776 744
rect 1780 742 1782 744
rect 1804 742 1806 744
rect 1810 742 1812 744
rect 1834 742 1836 744
rect 1840 742 1842 744
rect 1864 742 1866 744
rect 1870 742 1872 744
rect 1894 742 1896 744
rect 1900 742 1902 744
rect 1924 742 1926 744
rect 1930 742 1932 744
rect 1954 742 1956 744
rect 1960 742 1962 744
rect 1984 742 1986 744
rect 1612 740 1614 742
rect 1662 740 1664 742
rect 1692 740 1694 742
rect 1742 740 1744 742
rect 1772 740 1774 742
rect 1802 740 1804 742
rect 1832 740 1834 742
rect 1862 740 1864 742
rect 1892 740 1894 742
rect 1922 740 1924 742
rect 1952 740 1954 742
rect 1982 740 1984 742
rect 4622 738 4624 740
rect 4694 738 4696 740
rect 4724 738 4726 740
rect 4776 738 4778 740
rect 5222 738 5224 740
rect 5294 738 5296 740
rect 5324 738 5326 740
rect 5376 738 5378 740
rect 6422 738 6424 740
rect 6576 738 6578 740
rect 4620 736 4622 738
rect 4686 736 4688 738
rect 4692 736 4694 738
rect 4716 736 4718 738
rect 4722 736 4724 738
rect 4778 736 4780 738
rect 5220 736 5222 738
rect 5286 736 5288 738
rect 5292 736 5294 738
rect 5316 736 5318 738
rect 5322 736 5324 738
rect 5378 736 5380 738
rect 6420 736 6422 738
rect 6578 736 6580 738
rect 1612 734 1614 736
rect 1662 734 1664 736
rect 1742 734 1744 736
rect 1772 734 1774 736
rect 1802 734 1804 736
rect 1832 734 1834 736
rect 1862 734 1864 736
rect 1892 734 1894 736
rect 1922 734 1924 736
rect 1952 734 1954 736
rect 1982 734 1984 736
rect 4684 734 4686 736
rect 4714 734 4716 736
rect 5284 734 5286 736
rect 5314 734 5316 736
rect 1604 732 1606 734
rect 1610 732 1612 734
rect 1654 732 1656 734
rect 1660 732 1662 734
rect 1684 732 1686 734
rect 1720 732 1722 734
rect 1744 732 1746 734
rect 1750 732 1752 734
rect 1774 732 1776 734
rect 1780 732 1782 734
rect 1804 732 1806 734
rect 1810 732 1812 734
rect 1834 732 1836 734
rect 1840 732 1842 734
rect 1864 732 1866 734
rect 1870 732 1872 734
rect 1894 732 1896 734
rect 1900 732 1902 734
rect 1924 732 1926 734
rect 1930 732 1932 734
rect 1954 732 1956 734
rect 1960 732 1962 734
rect 1984 732 1986 734
rect 1602 730 1604 732
rect 1652 730 1654 732
rect 1682 730 1684 732
rect 1722 730 1724 732
rect 1752 730 1754 732
rect 1782 730 1784 732
rect 1812 730 1814 732
rect 1842 730 1844 732
rect 1872 730 1874 732
rect 1902 730 1904 732
rect 1932 730 1934 732
rect 1962 730 1964 732
rect 4684 728 4686 730
rect 4714 728 4716 730
rect 5284 728 5286 730
rect 5314 728 5316 730
rect 4620 726 4622 728
rect 4686 726 4688 728
rect 4692 726 4694 728
rect 4716 726 4718 728
rect 4722 726 4724 728
rect 4778 726 4780 728
rect 5220 726 5222 728
rect 5286 726 5288 728
rect 5292 726 5294 728
rect 5316 726 5318 728
rect 5322 726 5324 728
rect 5378 726 5380 728
rect 6420 726 6422 728
rect 6578 726 6580 728
rect 1602 724 1604 726
rect 1652 724 1654 726
rect 1722 724 1724 726
rect 1752 724 1754 726
rect 1782 724 1784 726
rect 1812 724 1814 726
rect 1842 724 1844 726
rect 1872 724 1874 726
rect 1902 724 1904 726
rect 1932 724 1934 726
rect 1962 724 1964 726
rect 4622 724 4624 726
rect 4694 724 4696 726
rect 4724 724 4726 726
rect 4776 724 4778 726
rect 5222 724 5224 726
rect 5294 724 5296 726
rect 5324 724 5326 726
rect 5376 724 5378 726
rect 6422 724 6424 726
rect 6576 724 6578 726
rect 1600 722 1602 724
rect 1644 722 1646 724
rect 1650 722 1652 724
rect 1674 722 1676 724
rect 1720 722 1722 724
rect 1744 722 1746 724
rect 1750 722 1752 724
rect 1774 722 1776 724
rect 1780 722 1782 724
rect 1804 722 1806 724
rect 1810 722 1812 724
rect 1834 722 1836 724
rect 1840 722 1842 724
rect 1864 722 1866 724
rect 1870 722 1872 724
rect 1894 722 1896 724
rect 1900 722 1902 724
rect 1924 722 1926 724
rect 1930 722 1932 724
rect 1954 722 1956 724
rect 1960 722 1962 724
rect 1984 722 1986 724
rect 1642 720 1644 722
rect 1672 720 1674 722
rect 1742 720 1744 722
rect 1772 720 1774 722
rect 1802 720 1804 722
rect 1832 720 1834 722
rect 1862 720 1864 722
rect 1892 720 1894 722
rect 1922 720 1924 722
rect 1952 720 1954 722
rect 1982 720 1984 722
rect 3242 718 3244 720
rect 3272 718 3274 720
rect 3302 718 3304 720
rect 3332 718 3334 720
rect 3362 718 3364 720
rect 3636 718 3638 720
rect 3666 718 3668 720
rect 3696 718 3698 720
rect 3726 718 3728 720
rect 3756 718 3758 720
rect 3842 718 3844 720
rect 3872 718 3874 720
rect 3902 718 3904 720
rect 3932 718 3934 720
rect 3962 718 3964 720
rect 4236 718 4238 720
rect 4266 718 4268 720
rect 4296 718 4298 720
rect 4326 718 4328 720
rect 4356 718 4358 720
rect 4442 718 4444 720
rect 4472 718 4474 720
rect 4502 718 4504 720
rect 4532 718 4534 720
rect 4562 718 4564 720
rect 4592 718 4594 720
rect 4622 718 4624 720
rect 4694 718 4696 720
rect 4724 718 4726 720
rect 4776 718 4778 720
rect 4806 718 4808 720
rect 4836 718 4838 720
rect 4866 718 4868 720
rect 4896 718 4898 720
rect 4926 718 4928 720
rect 4956 718 4958 720
rect 5042 718 5044 720
rect 5072 718 5074 720
rect 5102 718 5104 720
rect 5132 718 5134 720
rect 5162 718 5164 720
rect 5192 718 5194 720
rect 5222 718 5224 720
rect 5294 718 5296 720
rect 5324 718 5326 720
rect 5376 718 5378 720
rect 5406 718 5408 720
rect 5436 718 5438 720
rect 5466 718 5468 720
rect 5496 718 5498 720
rect 5526 718 5528 720
rect 5556 718 5558 720
rect 5642 718 5644 720
rect 5672 718 5674 720
rect 5702 718 5704 720
rect 5732 718 5734 720
rect 5762 718 5764 720
rect 6036 718 6038 720
rect 6066 718 6068 720
rect 6096 718 6098 720
rect 6126 718 6128 720
rect 6156 718 6158 720
rect 6242 718 6244 720
rect 6272 718 6274 720
rect 6302 718 6304 720
rect 6332 718 6334 720
rect 6362 718 6364 720
rect 6392 718 6394 720
rect 6422 718 6424 720
rect 6576 718 6578 720
rect 6606 718 6608 720
rect 6636 718 6638 720
rect 6666 718 6668 720
rect 6696 718 6698 720
rect 6726 718 6728 720
rect 6756 718 6758 720
rect 3234 716 3236 718
rect 3240 716 3242 718
rect 3264 716 3266 718
rect 3270 716 3272 718
rect 3294 716 3296 718
rect 3300 716 3302 718
rect 3324 716 3326 718
rect 3330 716 3332 718
rect 3354 716 3356 718
rect 3360 716 3362 718
rect 3384 716 3386 718
rect 3614 716 3616 718
rect 3638 716 3640 718
rect 3644 716 3646 718
rect 3668 716 3670 718
rect 3674 716 3676 718
rect 3698 716 3700 718
rect 3704 716 3706 718
rect 3728 716 3730 718
rect 3734 716 3736 718
rect 3758 716 3760 718
rect 3764 716 3766 718
rect 3834 716 3836 718
rect 3840 716 3842 718
rect 3864 716 3866 718
rect 3870 716 3872 718
rect 3894 716 3896 718
rect 3900 716 3902 718
rect 3924 716 3926 718
rect 3930 716 3932 718
rect 3954 716 3956 718
rect 3960 716 3962 718
rect 3984 716 3986 718
rect 4214 716 4216 718
rect 4238 716 4240 718
rect 4244 716 4246 718
rect 4268 716 4270 718
rect 4274 716 4276 718
rect 4298 716 4300 718
rect 4304 716 4306 718
rect 4328 716 4330 718
rect 4334 716 4336 718
rect 4358 716 4360 718
rect 4364 716 4366 718
rect 4434 716 4436 718
rect 4440 716 4442 718
rect 4464 716 4466 718
rect 4470 716 4472 718
rect 4494 716 4496 718
rect 4500 716 4502 718
rect 4524 716 4526 718
rect 4530 716 4532 718
rect 4554 716 4556 718
rect 4560 716 4562 718
rect 4584 716 4586 718
rect 4590 716 4592 718
rect 4614 716 4616 718
rect 4620 716 4622 718
rect 4686 716 4688 718
rect 4692 716 4694 718
rect 4716 716 4718 718
rect 4722 716 4724 718
rect 4778 716 4780 718
rect 4784 716 4786 718
rect 4808 716 4810 718
rect 4814 716 4816 718
rect 4838 716 4840 718
rect 4844 716 4846 718
rect 4868 716 4870 718
rect 4874 716 4876 718
rect 4898 716 4900 718
rect 4904 716 4906 718
rect 4928 716 4930 718
rect 4934 716 4936 718
rect 4958 716 4960 718
rect 4964 716 4966 718
rect 5034 716 5036 718
rect 5040 716 5042 718
rect 5064 716 5066 718
rect 5070 716 5072 718
rect 5094 716 5096 718
rect 5100 716 5102 718
rect 5124 716 5126 718
rect 5130 716 5132 718
rect 5154 716 5156 718
rect 5160 716 5162 718
rect 5184 716 5186 718
rect 5190 716 5192 718
rect 5214 716 5216 718
rect 5220 716 5222 718
rect 5286 716 5288 718
rect 5292 716 5294 718
rect 5316 716 5318 718
rect 5322 716 5324 718
rect 5378 716 5380 718
rect 5384 716 5386 718
rect 5408 716 5410 718
rect 5414 716 5416 718
rect 5438 716 5440 718
rect 5444 716 5446 718
rect 5468 716 5470 718
rect 5474 716 5476 718
rect 5498 716 5500 718
rect 5504 716 5506 718
rect 5528 716 5530 718
rect 5534 716 5536 718
rect 5558 716 5560 718
rect 5564 716 5566 718
rect 5634 716 5636 718
rect 5640 716 5642 718
rect 5664 716 5666 718
rect 5670 716 5672 718
rect 5694 716 5696 718
rect 5700 716 5702 718
rect 5724 716 5726 718
rect 5730 716 5732 718
rect 5754 716 5756 718
rect 5760 716 5762 718
rect 6038 716 6040 718
rect 6044 716 6046 718
rect 6068 716 6070 718
rect 6074 716 6076 718
rect 6098 716 6100 718
rect 6104 716 6106 718
rect 6128 716 6130 718
rect 6134 716 6136 718
rect 6158 716 6160 718
rect 6164 716 6166 718
rect 6234 716 6236 718
rect 6240 716 6242 718
rect 6264 716 6266 718
rect 6270 716 6272 718
rect 6294 716 6296 718
rect 6300 716 6302 718
rect 6324 716 6326 718
rect 6330 716 6332 718
rect 6354 716 6356 718
rect 6360 716 6362 718
rect 6384 716 6386 718
rect 6390 716 6392 718
rect 6414 716 6416 718
rect 6420 716 6422 718
rect 6578 716 6580 718
rect 6584 716 6586 718
rect 6608 716 6610 718
rect 6614 716 6616 718
rect 6638 716 6640 718
rect 6644 716 6646 718
rect 6668 716 6670 718
rect 6674 716 6676 718
rect 6698 716 6700 718
rect 6704 716 6706 718
rect 6728 716 6730 718
rect 6734 716 6736 718
rect 6758 716 6760 718
rect 6764 716 6766 718
rect 1642 714 1644 716
rect 1742 714 1744 716
rect 1772 714 1774 716
rect 1802 714 1804 716
rect 1832 714 1834 716
rect 1862 714 1864 716
rect 1892 714 1894 716
rect 1922 714 1924 716
rect 1952 714 1954 716
rect 1982 714 1984 716
rect 3232 714 3234 716
rect 3262 714 3264 716
rect 3292 714 3294 716
rect 3322 714 3324 716
rect 3352 714 3354 716
rect 3382 714 3384 716
rect 3616 714 3618 716
rect 3646 714 3648 716
rect 3676 714 3678 716
rect 3706 714 3708 716
rect 3736 714 3738 716
rect 3766 714 3768 716
rect 3832 714 3834 716
rect 3862 714 3864 716
rect 3892 714 3894 716
rect 3922 714 3924 716
rect 3952 714 3954 716
rect 3982 714 3984 716
rect 4216 714 4218 716
rect 4246 714 4248 716
rect 4276 714 4278 716
rect 4306 714 4308 716
rect 4336 714 4338 716
rect 4366 714 4368 716
rect 4432 714 4434 716
rect 4462 714 4464 716
rect 4492 714 4494 716
rect 4522 714 4524 716
rect 4552 714 4554 716
rect 4582 714 4584 716
rect 4612 714 4614 716
rect 4684 714 4686 716
rect 4714 714 4716 716
rect 4786 714 4788 716
rect 4816 714 4818 716
rect 4846 714 4848 716
rect 4876 714 4878 716
rect 4906 714 4908 716
rect 4936 714 4938 716
rect 4966 714 4968 716
rect 5032 714 5034 716
rect 5062 714 5064 716
rect 5092 714 5094 716
rect 5122 714 5124 716
rect 5152 714 5154 716
rect 5182 714 5184 716
rect 5212 714 5214 716
rect 5284 714 5286 716
rect 5314 714 5316 716
rect 5386 714 5388 716
rect 5416 714 5418 716
rect 5446 714 5448 716
rect 5476 714 5478 716
rect 5506 714 5508 716
rect 5536 714 5538 716
rect 5566 714 5568 716
rect 5632 714 5634 716
rect 5662 714 5664 716
rect 5692 714 5694 716
rect 5722 714 5724 716
rect 5752 714 5754 716
rect 6046 714 6048 716
rect 6076 714 6078 716
rect 6106 714 6108 716
rect 6136 714 6138 716
rect 6166 714 6168 716
rect 6232 714 6234 716
rect 6262 714 6264 716
rect 6292 714 6294 716
rect 6322 714 6324 716
rect 6352 714 6354 716
rect 6382 714 6384 716
rect 6412 714 6414 716
rect 6586 714 6588 716
rect 6616 714 6618 716
rect 6646 714 6648 716
rect 6676 714 6678 716
rect 6706 714 6708 716
rect 6736 714 6738 716
rect 6766 714 6768 716
rect 1634 712 1636 714
rect 1640 712 1642 714
rect 1664 712 1666 714
rect 1720 712 1722 714
rect 1744 712 1746 714
rect 1750 712 1752 714
rect 1774 712 1776 714
rect 1780 712 1782 714
rect 1804 712 1806 714
rect 1810 712 1812 714
rect 1834 712 1836 714
rect 1840 712 1842 714
rect 1864 712 1866 714
rect 1870 712 1872 714
rect 1894 712 1896 714
rect 1900 712 1902 714
rect 1924 712 1926 714
rect 1930 712 1932 714
rect 1954 712 1956 714
rect 1960 712 1962 714
rect 1984 712 1986 714
rect 1632 710 1634 712
rect 1662 710 1664 712
rect 1722 710 1724 712
rect 1752 710 1754 712
rect 1782 710 1784 712
rect 1812 710 1814 712
rect 1842 710 1844 712
rect 1872 710 1874 712
rect 1902 710 1904 712
rect 1932 710 1934 712
rect 1962 710 1964 712
rect 3232 708 3234 710
rect 3262 708 3264 710
rect 3292 708 3294 710
rect 3322 708 3324 710
rect 3352 708 3354 710
rect 3382 708 3384 710
rect 3616 708 3618 710
rect 3646 708 3648 710
rect 3676 708 3678 710
rect 3706 708 3708 710
rect 3736 708 3738 710
rect 3766 708 3768 710
rect 3832 708 3834 710
rect 3862 708 3864 710
rect 3892 708 3894 710
rect 3922 708 3924 710
rect 3952 708 3954 710
rect 3982 708 3984 710
rect 4216 708 4218 710
rect 4246 708 4248 710
rect 4276 708 4278 710
rect 4306 708 4308 710
rect 4336 708 4338 710
rect 4366 708 4368 710
rect 4432 708 4434 710
rect 4462 708 4464 710
rect 4492 708 4494 710
rect 4522 708 4524 710
rect 4552 708 4554 710
rect 4582 708 4584 710
rect 4612 708 4614 710
rect 4684 708 4686 710
rect 4714 708 4716 710
rect 4786 708 4788 710
rect 4816 708 4818 710
rect 4846 708 4848 710
rect 4876 708 4878 710
rect 4906 708 4908 710
rect 4936 708 4938 710
rect 4966 708 4968 710
rect 5032 708 5034 710
rect 5062 708 5064 710
rect 5092 708 5094 710
rect 5122 708 5124 710
rect 5152 708 5154 710
rect 5182 708 5184 710
rect 5212 708 5214 710
rect 5284 708 5286 710
rect 5314 708 5316 710
rect 5386 708 5388 710
rect 5416 708 5418 710
rect 5446 708 5448 710
rect 5476 708 5478 710
rect 5506 708 5508 710
rect 5536 708 5538 710
rect 5566 708 5568 710
rect 5632 708 5634 710
rect 5662 708 5664 710
rect 5692 708 5694 710
rect 5722 708 5724 710
rect 5752 708 5754 710
rect 6046 708 6048 710
rect 6076 708 6078 710
rect 6106 708 6108 710
rect 6136 708 6138 710
rect 6166 708 6168 710
rect 6232 708 6234 710
rect 6262 708 6264 710
rect 6292 708 6294 710
rect 6322 708 6324 710
rect 6352 708 6354 710
rect 6382 708 6384 710
rect 6412 708 6414 710
rect 6586 708 6588 710
rect 6616 708 6618 710
rect 6646 708 6648 710
rect 6676 708 6678 710
rect 6706 708 6708 710
rect 6736 708 6738 710
rect 6766 708 6768 710
rect 3234 706 3236 708
rect 3240 706 3242 708
rect 3264 706 3266 708
rect 3270 706 3272 708
rect 3294 706 3296 708
rect 3300 706 3302 708
rect 3324 706 3326 708
rect 3330 706 3332 708
rect 3354 706 3356 708
rect 3360 706 3362 708
rect 3384 706 3386 708
rect 3614 706 3616 708
rect 3638 706 3640 708
rect 3644 706 3646 708
rect 3668 706 3670 708
rect 3674 706 3676 708
rect 3698 706 3700 708
rect 3704 706 3706 708
rect 3728 706 3730 708
rect 3734 706 3736 708
rect 3758 706 3760 708
rect 3764 706 3766 708
rect 3834 706 3836 708
rect 3840 706 3842 708
rect 3864 706 3866 708
rect 3870 706 3872 708
rect 3894 706 3896 708
rect 3900 706 3902 708
rect 3924 706 3926 708
rect 3930 706 3932 708
rect 3954 706 3956 708
rect 3960 706 3962 708
rect 3984 706 3986 708
rect 4214 706 4216 708
rect 4238 706 4240 708
rect 4244 706 4246 708
rect 4268 706 4270 708
rect 4274 706 4276 708
rect 4298 706 4300 708
rect 4304 706 4306 708
rect 4328 706 4330 708
rect 4334 706 4336 708
rect 4358 706 4360 708
rect 4364 706 4366 708
rect 4434 706 4436 708
rect 4440 706 4442 708
rect 4464 706 4466 708
rect 4470 706 4472 708
rect 4494 706 4496 708
rect 4500 706 4502 708
rect 4524 706 4526 708
rect 4530 706 4532 708
rect 4554 706 4556 708
rect 4560 706 4562 708
rect 4584 706 4586 708
rect 4590 706 4592 708
rect 4614 706 4616 708
rect 4620 706 4622 708
rect 4686 706 4688 708
rect 4692 706 4694 708
rect 4716 706 4718 708
rect 4722 706 4724 708
rect 4778 706 4780 708
rect 4784 706 4786 708
rect 4808 706 4810 708
rect 4814 706 4816 708
rect 4838 706 4840 708
rect 4844 706 4846 708
rect 4868 706 4870 708
rect 4874 706 4876 708
rect 4898 706 4900 708
rect 4904 706 4906 708
rect 4928 706 4930 708
rect 4934 706 4936 708
rect 4958 706 4960 708
rect 4964 706 4966 708
rect 5034 706 5036 708
rect 5040 706 5042 708
rect 5064 706 5066 708
rect 5070 706 5072 708
rect 5094 706 5096 708
rect 5100 706 5102 708
rect 5124 706 5126 708
rect 5130 706 5132 708
rect 5154 706 5156 708
rect 5160 706 5162 708
rect 5184 706 5186 708
rect 5190 706 5192 708
rect 5214 706 5216 708
rect 5220 706 5222 708
rect 5286 706 5288 708
rect 5292 706 5294 708
rect 5316 706 5318 708
rect 5322 706 5324 708
rect 5378 706 5380 708
rect 5384 706 5386 708
rect 5408 706 5410 708
rect 5414 706 5416 708
rect 5438 706 5440 708
rect 5444 706 5446 708
rect 5468 706 5470 708
rect 5474 706 5476 708
rect 5498 706 5500 708
rect 5504 706 5506 708
rect 5528 706 5530 708
rect 5534 706 5536 708
rect 5558 706 5560 708
rect 5564 706 5566 708
rect 5634 706 5636 708
rect 5640 706 5642 708
rect 5664 706 5666 708
rect 5670 706 5672 708
rect 5694 706 5696 708
rect 5700 706 5702 708
rect 5724 706 5726 708
rect 5730 706 5732 708
rect 5754 706 5756 708
rect 5760 706 5762 708
rect 5896 706 5898 708
rect 5902 706 5904 708
rect 6038 706 6040 708
rect 6044 706 6046 708
rect 6068 706 6070 708
rect 6074 706 6076 708
rect 6098 706 6100 708
rect 6104 706 6106 708
rect 6128 706 6130 708
rect 6134 706 6136 708
rect 6158 706 6160 708
rect 6164 706 6166 708
rect 6234 706 6236 708
rect 6240 706 6242 708
rect 6264 706 6266 708
rect 6270 706 6272 708
rect 6294 706 6296 708
rect 6300 706 6302 708
rect 6324 706 6326 708
rect 6330 706 6332 708
rect 6354 706 6356 708
rect 6360 706 6362 708
rect 6384 706 6386 708
rect 6390 706 6392 708
rect 6414 706 6416 708
rect 6420 706 6422 708
rect 6578 706 6580 708
rect 6584 706 6586 708
rect 6608 706 6610 708
rect 6614 706 6616 708
rect 6638 706 6640 708
rect 6644 706 6646 708
rect 6668 706 6670 708
rect 6674 706 6676 708
rect 6698 706 6700 708
rect 6704 706 6706 708
rect 6728 706 6730 708
rect 6734 706 6736 708
rect 6758 706 6760 708
rect 6764 706 6766 708
rect 1632 704 1634 706
rect 1692 704 1694 706
rect 1702 704 1704 706
rect 1722 704 1724 706
rect 1752 704 1754 706
rect 1782 704 1784 706
rect 1812 704 1814 706
rect 1842 704 1844 706
rect 1872 704 1874 706
rect 1902 704 1904 706
rect 1932 704 1934 706
rect 1962 704 1964 706
rect 1624 702 1626 704
rect 1630 702 1632 704
rect 1654 702 1656 704
rect 1690 702 1692 704
rect 1704 702 1706 704
rect 1720 702 1722 704
rect 1744 702 1746 704
rect 1750 702 1752 704
rect 1774 702 1776 704
rect 1780 702 1782 704
rect 1804 702 1806 704
rect 1810 702 1812 704
rect 1834 702 1836 704
rect 1840 702 1842 704
rect 1864 702 1866 704
rect 1870 702 1872 704
rect 1894 702 1896 704
rect 1900 702 1902 704
rect 1924 702 1926 704
rect 1930 702 1932 704
rect 1954 702 1956 704
rect 1960 702 1962 704
rect 1984 702 1986 704
rect 2586 703 2598 705
rect 3186 703 3198 705
rect 3242 704 3244 706
rect 3272 704 3274 706
rect 3302 704 3304 706
rect 3332 704 3334 706
rect 3362 704 3364 706
rect 3636 704 3638 706
rect 3666 704 3668 706
rect 3696 704 3698 706
rect 3726 704 3728 706
rect 3756 704 3758 706
rect 3842 704 3844 706
rect 3872 704 3874 706
rect 3902 704 3904 706
rect 3932 704 3934 706
rect 3962 704 3964 706
rect 4236 704 4238 706
rect 4266 704 4268 706
rect 4296 704 4298 706
rect 4326 704 4328 706
rect 4356 704 4358 706
rect 4442 704 4444 706
rect 4472 704 4474 706
rect 4502 704 4504 706
rect 4532 704 4534 706
rect 4562 704 4564 706
rect 4592 704 4594 706
rect 4622 704 4624 706
rect 4694 704 4696 706
rect 4724 704 4726 706
rect 4776 704 4778 706
rect 4806 704 4808 706
rect 4836 704 4838 706
rect 4866 704 4868 706
rect 4896 704 4898 706
rect 4926 704 4928 706
rect 4956 704 4958 706
rect 5042 704 5044 706
rect 5072 704 5074 706
rect 5102 704 5104 706
rect 5132 704 5134 706
rect 5162 704 5164 706
rect 5192 704 5194 706
rect 5222 704 5224 706
rect 5294 704 5296 706
rect 5324 704 5326 706
rect 5376 704 5378 706
rect 5406 704 5408 706
rect 5436 704 5438 706
rect 5466 704 5468 706
rect 5496 704 5498 706
rect 5526 704 5528 706
rect 5556 704 5558 706
rect 5642 704 5644 706
rect 5672 704 5674 706
rect 5702 704 5704 706
rect 5732 704 5734 706
rect 5762 704 5764 706
rect 5894 704 5896 706
rect 5904 704 5906 706
rect 6036 704 6038 706
rect 6066 704 6068 706
rect 6096 704 6098 706
rect 6126 704 6128 706
rect 6156 704 6158 706
rect 6242 704 6244 706
rect 6272 704 6274 706
rect 6302 704 6304 706
rect 6332 704 6334 706
rect 6362 704 6364 706
rect 6392 704 6394 706
rect 6422 704 6424 706
rect 6576 704 6578 706
rect 6606 704 6608 706
rect 6636 704 6638 706
rect 6666 704 6668 706
rect 6696 704 6698 706
rect 6726 704 6728 706
rect 6756 704 6758 706
rect 1622 700 1624 702
rect 1652 700 1654 702
rect 1742 700 1744 702
rect 1772 700 1774 702
rect 1802 700 1804 702
rect 1832 700 1834 702
rect 1862 700 1864 702
rect 1892 700 1894 702
rect 1922 700 1924 702
rect 1952 700 1954 702
rect 1982 700 1984 702
rect 2588 701 2590 703
rect 3188 701 3190 703
rect 2094 700 2096 701
rect 2126 700 2128 701
rect 2132 700 2134 701
rect 2158 700 2160 701
rect 2164 700 2166 701
rect 2222 700 2224 701
rect 2228 700 2230 701
rect 2694 700 2696 701
rect 2726 700 2728 701
rect 2732 700 2734 701
rect 2758 700 2760 701
rect 2764 700 2766 701
rect 2822 700 2824 701
rect 2828 700 2830 701
rect 6894 700 6896 701
rect 6926 700 6928 701
rect 6932 700 6934 701
rect 6958 700 6960 701
rect 6964 700 6966 701
rect 7022 700 7024 701
rect 7028 700 7030 701
rect 2588 697 2590 699
rect 3188 697 3190 699
rect 3242 698 3244 700
rect 3272 698 3274 700
rect 3302 698 3304 700
rect 3332 698 3334 700
rect 3362 698 3364 700
rect 3636 698 3638 700
rect 3666 698 3668 700
rect 3696 698 3698 700
rect 3726 698 3728 700
rect 3756 698 3758 700
rect 3842 698 3844 700
rect 3872 698 3874 700
rect 3902 698 3904 700
rect 3932 698 3934 700
rect 3962 698 3964 700
rect 4236 698 4238 700
rect 4266 698 4268 700
rect 4296 698 4298 700
rect 4326 698 4328 700
rect 4356 698 4358 700
rect 4442 698 4444 700
rect 4472 698 4474 700
rect 4502 698 4504 700
rect 4532 698 4534 700
rect 4562 698 4564 700
rect 4592 698 4594 700
rect 4622 698 4624 700
rect 4694 698 4696 700
rect 4724 698 4726 700
rect 4776 698 4778 700
rect 4806 698 4808 700
rect 4836 698 4838 700
rect 4866 698 4868 700
rect 4896 698 4898 700
rect 4926 698 4928 700
rect 4956 698 4958 700
rect 5042 698 5044 700
rect 5072 698 5074 700
rect 5102 698 5104 700
rect 5132 698 5134 700
rect 5162 698 5164 700
rect 5192 698 5194 700
rect 5222 698 5224 700
rect 5294 698 5296 700
rect 5324 698 5326 700
rect 5376 698 5378 700
rect 5406 698 5408 700
rect 5436 698 5438 700
rect 5466 698 5468 700
rect 5496 698 5498 700
rect 5526 698 5528 700
rect 5556 698 5558 700
rect 5642 698 5644 700
rect 5672 698 5674 700
rect 5702 698 5704 700
rect 5732 698 5734 700
rect 5762 698 5764 700
rect 6036 698 6038 700
rect 6066 698 6068 700
rect 6096 698 6098 700
rect 6126 698 6128 700
rect 6156 698 6158 700
rect 6242 698 6244 700
rect 6272 698 6274 700
rect 6302 698 6304 700
rect 6332 698 6334 700
rect 6362 698 6364 700
rect 6392 698 6394 700
rect 6422 698 6424 700
rect 6576 698 6578 700
rect 6606 698 6608 700
rect 6636 698 6638 700
rect 6666 698 6668 700
rect 6696 698 6698 700
rect 6726 698 6728 700
rect 6756 698 6758 700
rect 1622 694 1624 696
rect 1682 694 1684 696
rect 1712 694 1714 696
rect 1742 694 1744 696
rect 1772 694 1774 696
rect 2590 695 2592 697
rect 3190 695 3192 697
rect 3234 696 3236 698
rect 3240 696 3242 698
rect 3264 696 3266 698
rect 3270 696 3272 698
rect 3294 696 3296 698
rect 3300 696 3302 698
rect 3324 696 3326 698
rect 3330 696 3332 698
rect 3354 696 3356 698
rect 3360 696 3362 698
rect 3384 696 3386 698
rect 3614 696 3616 698
rect 3638 696 3640 698
rect 3644 696 3646 698
rect 3668 696 3670 698
rect 3674 696 3676 698
rect 3698 696 3700 698
rect 3704 696 3706 698
rect 3728 696 3730 698
rect 3734 696 3736 698
rect 3758 696 3760 698
rect 3764 696 3766 698
rect 3834 696 3836 698
rect 3840 696 3842 698
rect 3864 696 3866 698
rect 3870 696 3872 698
rect 3894 696 3896 698
rect 3900 696 3902 698
rect 3924 696 3926 698
rect 3930 696 3932 698
rect 3954 696 3956 698
rect 3960 696 3962 698
rect 3984 696 3986 698
rect 4214 696 4216 698
rect 4238 696 4240 698
rect 4244 696 4246 698
rect 4268 696 4270 698
rect 4274 696 4276 698
rect 4298 696 4300 698
rect 4304 696 4306 698
rect 4328 696 4330 698
rect 4334 696 4336 698
rect 4358 696 4360 698
rect 4364 696 4366 698
rect 4434 696 4436 698
rect 4440 696 4442 698
rect 4464 696 4466 698
rect 4470 696 4472 698
rect 4494 696 4496 698
rect 4500 696 4502 698
rect 4524 696 4526 698
rect 4530 696 4532 698
rect 4554 696 4556 698
rect 4560 696 4562 698
rect 4584 696 4586 698
rect 4590 696 4592 698
rect 4614 696 4616 698
rect 4620 696 4622 698
rect 4686 696 4688 698
rect 4692 696 4694 698
rect 4716 696 4718 698
rect 4722 696 4724 698
rect 4778 696 4780 698
rect 4784 696 4786 698
rect 4808 696 4810 698
rect 4814 696 4816 698
rect 4838 696 4840 698
rect 4844 696 4846 698
rect 4868 696 4870 698
rect 4874 696 4876 698
rect 4898 696 4900 698
rect 4904 696 4906 698
rect 4928 696 4930 698
rect 4934 696 4936 698
rect 4958 696 4960 698
rect 4964 696 4966 698
rect 5034 696 5036 698
rect 5040 696 5042 698
rect 5064 696 5066 698
rect 5070 696 5072 698
rect 5094 696 5096 698
rect 5100 696 5102 698
rect 5124 696 5126 698
rect 5130 696 5132 698
rect 5154 696 5156 698
rect 5160 696 5162 698
rect 5184 696 5186 698
rect 5190 696 5192 698
rect 5214 696 5216 698
rect 5220 696 5222 698
rect 5286 696 5288 698
rect 5292 696 5294 698
rect 5316 696 5318 698
rect 5322 696 5324 698
rect 5378 696 5380 698
rect 5384 696 5386 698
rect 5408 696 5410 698
rect 5414 696 5416 698
rect 5438 696 5440 698
rect 5444 696 5446 698
rect 5468 696 5470 698
rect 5474 696 5476 698
rect 5498 696 5500 698
rect 5504 696 5506 698
rect 5528 696 5530 698
rect 5534 696 5536 698
rect 5558 696 5560 698
rect 5564 696 5566 698
rect 5634 696 5636 698
rect 5640 696 5642 698
rect 5664 696 5666 698
rect 5670 696 5672 698
rect 5694 696 5696 698
rect 5700 696 5702 698
rect 5724 696 5726 698
rect 5730 696 5732 698
rect 5754 696 5756 698
rect 5760 696 5762 698
rect 6038 696 6040 698
rect 6044 696 6046 698
rect 6068 696 6070 698
rect 6074 696 6076 698
rect 6098 696 6100 698
rect 6104 696 6106 698
rect 6128 696 6130 698
rect 6134 696 6136 698
rect 6158 696 6160 698
rect 6164 696 6166 698
rect 6234 696 6236 698
rect 6240 696 6242 698
rect 6264 696 6266 698
rect 6270 696 6272 698
rect 6294 696 6296 698
rect 6300 696 6302 698
rect 6324 696 6326 698
rect 6330 696 6332 698
rect 6354 696 6356 698
rect 6360 696 6362 698
rect 6384 696 6386 698
rect 6390 696 6392 698
rect 6414 696 6416 698
rect 6420 696 6422 698
rect 6578 696 6580 698
rect 6584 696 6586 698
rect 6608 696 6610 698
rect 6614 696 6616 698
rect 6638 696 6640 698
rect 6644 696 6646 698
rect 6668 696 6670 698
rect 6674 696 6676 698
rect 6698 696 6700 698
rect 6704 696 6706 698
rect 6728 696 6730 698
rect 6734 696 6736 698
rect 6758 696 6760 698
rect 6764 696 6766 698
rect 3232 694 3234 696
rect 3262 694 3264 696
rect 3292 694 3294 696
rect 3322 694 3324 696
rect 3352 694 3354 696
rect 3382 694 3384 696
rect 3616 694 3618 696
rect 3646 694 3648 696
rect 3676 694 3678 696
rect 3706 694 3708 696
rect 3736 694 3738 696
rect 3766 694 3768 696
rect 3832 694 3834 696
rect 3862 694 3864 696
rect 3892 694 3894 696
rect 3922 694 3924 696
rect 3952 694 3954 696
rect 3982 694 3984 696
rect 4216 694 4218 696
rect 4246 694 4248 696
rect 4276 694 4278 696
rect 4306 694 4308 696
rect 4336 694 4338 696
rect 4366 694 4368 696
rect 4432 694 4434 696
rect 4462 694 4464 696
rect 4492 694 4494 696
rect 4522 694 4524 696
rect 4552 694 4554 696
rect 4582 694 4584 696
rect 4612 694 4614 696
rect 4684 694 4686 696
rect 4714 694 4716 696
rect 4786 694 4788 696
rect 4816 694 4818 696
rect 4846 694 4848 696
rect 4876 694 4878 696
rect 4906 694 4908 696
rect 4936 694 4938 696
rect 4966 694 4968 696
rect 5032 694 5034 696
rect 5062 694 5064 696
rect 5092 694 5094 696
rect 5122 694 5124 696
rect 5152 694 5154 696
rect 5182 694 5184 696
rect 5212 694 5214 696
rect 5284 694 5286 696
rect 5314 694 5316 696
rect 5386 694 5388 696
rect 5416 694 5418 696
rect 5446 694 5448 696
rect 5476 694 5478 696
rect 5506 694 5508 696
rect 5536 694 5538 696
rect 5566 694 5568 696
rect 5632 694 5634 696
rect 5662 694 5664 696
rect 5692 694 5694 696
rect 5722 694 5724 696
rect 5752 694 5754 696
rect 6046 694 6048 696
rect 6076 694 6078 696
rect 6106 694 6108 696
rect 6136 694 6138 696
rect 6166 694 6168 696
rect 6232 694 6234 696
rect 6262 694 6264 696
rect 6292 694 6294 696
rect 6322 694 6324 696
rect 6352 694 6354 696
rect 6382 694 6384 696
rect 6412 694 6414 696
rect 6586 694 6588 696
rect 6616 694 6618 696
rect 6646 694 6648 696
rect 6676 694 6678 696
rect 6706 694 6708 696
rect 6736 694 6738 696
rect 6766 694 6768 696
rect 1624 692 1626 694
rect 1680 692 1682 694
rect 1714 692 1716 694
rect 1740 692 1742 694
rect 1774 692 1776 694
rect 1672 684 1674 686
rect 1644 682 1646 684
rect 1670 682 1672 684
rect 2549 683 2550 684
rect 3149 683 3150 684
rect 1642 680 1644 682
rect 1662 674 1664 676
rect 1634 672 1636 674
rect 1660 672 1662 674
rect 1632 670 1634 672
rect 2555 670 2556 671
rect 3155 670 3156 671
rect 1652 664 1654 666
rect 1624 662 1626 664
rect 1650 662 1652 664
rect 1622 660 1624 662
rect 2588 656 2590 658
rect 3188 656 3190 658
rect 1642 654 1644 656
rect 2590 654 2592 656
rect 3190 654 3192 656
rect 1614 652 1616 654
rect 1640 652 1642 654
rect 1612 650 1614 652
rect 1632 644 1634 646
rect 3232 644 3234 646
rect 3262 644 3264 646
rect 3292 644 3294 646
rect 3322 644 3324 646
rect 3352 644 3354 646
rect 3382 644 3384 646
rect 3616 644 3618 646
rect 3646 644 3648 646
rect 3676 644 3678 646
rect 3706 644 3708 646
rect 3736 644 3738 646
rect 3766 644 3768 646
rect 3832 644 3834 646
rect 3862 644 3864 646
rect 3892 644 3894 646
rect 3922 644 3924 646
rect 3952 644 3954 646
rect 3982 644 3984 646
rect 4216 644 4218 646
rect 4246 644 4248 646
rect 4276 644 4278 646
rect 4306 644 4308 646
rect 4336 644 4338 646
rect 4366 644 4368 646
rect 4432 644 4434 646
rect 4462 644 4464 646
rect 4492 644 4494 646
rect 4522 644 4524 646
rect 4552 644 4554 646
rect 4582 644 4584 646
rect 4612 644 4614 646
rect 4684 644 4686 646
rect 4714 644 4716 646
rect 4786 644 4788 646
rect 4816 644 4818 646
rect 4846 644 4848 646
rect 4876 644 4878 646
rect 4906 644 4908 646
rect 4936 644 4938 646
rect 4966 644 4968 646
rect 5032 644 5034 646
rect 5062 644 5064 646
rect 5092 644 5094 646
rect 5122 644 5124 646
rect 5152 644 5154 646
rect 5182 644 5184 646
rect 5212 644 5214 646
rect 5284 644 5286 646
rect 5314 644 5316 646
rect 5386 644 5388 646
rect 5416 644 5418 646
rect 5446 644 5448 646
rect 5476 644 5478 646
rect 5506 644 5508 646
rect 5536 644 5538 646
rect 5566 644 5568 646
rect 5632 644 5634 646
rect 5662 644 5664 646
rect 5692 644 5694 646
rect 5722 644 5724 646
rect 5752 644 5754 646
rect 5782 644 5784 646
rect 5812 644 5814 646
rect 5884 644 5886 646
rect 5914 644 5916 646
rect 5986 644 5988 646
rect 6016 644 6018 646
rect 6046 644 6048 646
rect 6076 644 6078 646
rect 6106 644 6108 646
rect 6136 644 6138 646
rect 6166 644 6168 646
rect 6232 644 6234 646
rect 6262 644 6264 646
rect 6292 644 6294 646
rect 6322 644 6324 646
rect 6352 644 6354 646
rect 6382 644 6384 646
rect 6616 644 6618 646
rect 6646 644 6648 646
rect 6676 644 6678 646
rect 6706 644 6708 646
rect 6736 644 6738 646
rect 6766 644 6768 646
rect 1604 642 1606 644
rect 1630 642 1632 644
rect 3234 642 3236 644
rect 3240 642 3242 644
rect 3264 642 3266 644
rect 3270 642 3272 644
rect 3294 642 3296 644
rect 3300 642 3302 644
rect 3324 642 3326 644
rect 3330 642 3332 644
rect 3354 642 3356 644
rect 3360 642 3362 644
rect 3384 642 3386 644
rect 3614 642 3616 644
rect 3638 642 3640 644
rect 3644 642 3646 644
rect 3668 642 3670 644
rect 3674 642 3676 644
rect 3698 642 3700 644
rect 3704 642 3706 644
rect 3728 642 3730 644
rect 3734 642 3736 644
rect 3758 642 3760 644
rect 3764 642 3766 644
rect 3834 642 3836 644
rect 3840 642 3842 644
rect 3864 642 3866 644
rect 3870 642 3872 644
rect 3894 642 3896 644
rect 3900 642 3902 644
rect 3924 642 3926 644
rect 3930 642 3932 644
rect 3954 642 3956 644
rect 3960 642 3962 644
rect 3984 642 3986 644
rect 4214 642 4216 644
rect 4238 642 4240 644
rect 4244 642 4246 644
rect 4268 642 4270 644
rect 4274 642 4276 644
rect 4298 642 4300 644
rect 4304 642 4306 644
rect 4328 642 4330 644
rect 4334 642 4336 644
rect 4358 642 4360 644
rect 4364 642 4366 644
rect 4434 642 4436 644
rect 4440 642 4442 644
rect 4464 642 4466 644
rect 4470 642 4472 644
rect 4494 642 4496 644
rect 4500 642 4502 644
rect 4524 642 4526 644
rect 4530 642 4532 644
rect 4554 642 4556 644
rect 4560 642 4562 644
rect 4584 642 4586 644
rect 4590 642 4592 644
rect 4614 642 4616 644
rect 4620 642 4622 644
rect 4686 642 4688 644
rect 4692 642 4694 644
rect 4716 642 4718 644
rect 4722 642 4724 644
rect 4778 642 4780 644
rect 4784 642 4786 644
rect 4808 642 4810 644
rect 4814 642 4816 644
rect 4838 642 4840 644
rect 4844 642 4846 644
rect 4868 642 4870 644
rect 4874 642 4876 644
rect 4898 642 4900 644
rect 4904 642 4906 644
rect 4928 642 4930 644
rect 4934 642 4936 644
rect 4958 642 4960 644
rect 4964 642 4966 644
rect 5034 642 5036 644
rect 5040 642 5042 644
rect 5064 642 5066 644
rect 5070 642 5072 644
rect 5094 642 5096 644
rect 5100 642 5102 644
rect 5124 642 5126 644
rect 5130 642 5132 644
rect 5154 642 5156 644
rect 5160 642 5162 644
rect 5184 642 5186 644
rect 5190 642 5192 644
rect 5214 642 5216 644
rect 5220 642 5222 644
rect 5286 642 5288 644
rect 5292 642 5294 644
rect 5316 642 5318 644
rect 5322 642 5324 644
rect 5378 642 5380 644
rect 5384 642 5386 644
rect 5408 642 5410 644
rect 5414 642 5416 644
rect 5438 642 5440 644
rect 5444 642 5446 644
rect 5468 642 5470 644
rect 5474 642 5476 644
rect 5498 642 5500 644
rect 5504 642 5506 644
rect 5528 642 5530 644
rect 5534 642 5536 644
rect 5558 642 5560 644
rect 5564 642 5566 644
rect 5634 642 5636 644
rect 5640 642 5642 644
rect 5664 642 5666 644
rect 5670 642 5672 644
rect 5694 642 5696 644
rect 5700 642 5702 644
rect 5724 642 5726 644
rect 5730 642 5732 644
rect 5754 642 5756 644
rect 5760 642 5762 644
rect 5784 642 5786 644
rect 5790 642 5792 644
rect 5814 642 5816 644
rect 5820 642 5822 644
rect 5886 642 5888 644
rect 5892 642 5894 644
rect 5916 642 5918 644
rect 5922 642 5924 644
rect 5978 642 5980 644
rect 5984 642 5986 644
rect 6008 642 6010 644
rect 6014 642 6016 644
rect 6038 642 6040 644
rect 6044 642 6046 644
rect 6068 642 6070 644
rect 6074 642 6076 644
rect 6098 642 6100 644
rect 6104 642 6106 644
rect 6128 642 6130 644
rect 6134 642 6136 644
rect 6158 642 6160 644
rect 6164 642 6166 644
rect 6234 642 6236 644
rect 6240 642 6242 644
rect 6264 642 6266 644
rect 6270 642 6272 644
rect 6294 642 6296 644
rect 6300 642 6302 644
rect 6324 642 6326 644
rect 6330 642 6332 644
rect 6354 642 6356 644
rect 6360 642 6362 644
rect 6384 642 6386 644
rect 6614 642 6616 644
rect 6638 642 6640 644
rect 6644 642 6646 644
rect 6668 642 6670 644
rect 6674 642 6676 644
rect 6698 642 6700 644
rect 6704 642 6706 644
rect 6728 642 6730 644
rect 6734 642 6736 644
rect 6758 642 6760 644
rect 6764 642 6766 644
rect 1602 640 1604 642
rect 3242 640 3244 642
rect 3272 640 3274 642
rect 3302 640 3304 642
rect 3332 640 3334 642
rect 3362 640 3364 642
rect 3636 640 3638 642
rect 3666 640 3668 642
rect 3696 640 3698 642
rect 3726 640 3728 642
rect 3756 640 3758 642
rect 3842 640 3844 642
rect 3872 640 3874 642
rect 3902 640 3904 642
rect 3932 640 3934 642
rect 3962 640 3964 642
rect 4236 640 4238 642
rect 4266 640 4268 642
rect 4296 640 4298 642
rect 4326 640 4328 642
rect 4356 640 4358 642
rect 4442 640 4444 642
rect 4472 640 4474 642
rect 4502 640 4504 642
rect 4532 640 4534 642
rect 4562 640 4564 642
rect 4592 640 4594 642
rect 4622 640 4624 642
rect 4694 640 4696 642
rect 4724 640 4726 642
rect 4776 640 4778 642
rect 4806 640 4808 642
rect 4836 640 4838 642
rect 4866 640 4868 642
rect 4896 640 4898 642
rect 4926 640 4928 642
rect 4956 640 4958 642
rect 5042 640 5044 642
rect 5072 640 5074 642
rect 5102 640 5104 642
rect 5132 640 5134 642
rect 5162 640 5164 642
rect 5192 640 5194 642
rect 5222 640 5224 642
rect 5294 640 5296 642
rect 5324 640 5326 642
rect 5376 640 5378 642
rect 5406 640 5408 642
rect 5436 640 5438 642
rect 5466 640 5468 642
rect 5496 640 5498 642
rect 5526 640 5528 642
rect 5556 640 5558 642
rect 5642 640 5644 642
rect 5672 640 5674 642
rect 5702 640 5704 642
rect 5732 640 5734 642
rect 5762 640 5764 642
rect 5792 640 5794 642
rect 5822 640 5824 642
rect 5894 640 5896 642
rect 5924 640 5926 642
rect 5976 640 5978 642
rect 6006 640 6008 642
rect 6036 640 6038 642
rect 6066 640 6068 642
rect 6096 640 6098 642
rect 6126 640 6128 642
rect 6156 640 6158 642
rect 6242 640 6244 642
rect 6272 640 6274 642
rect 6302 640 6304 642
rect 6332 640 6334 642
rect 6362 640 6364 642
rect 6636 640 6638 642
rect 6666 640 6668 642
rect 6696 640 6698 642
rect 6726 640 6728 642
rect 6756 640 6758 642
rect 1622 634 1624 636
rect 1848 634 1850 636
rect 1878 634 1880 636
rect 1908 634 1910 636
rect 1938 634 1940 636
rect 1968 634 1970 636
rect 3242 634 3244 636
rect 3272 634 3274 636
rect 3302 634 3304 636
rect 3332 634 3334 636
rect 3362 634 3364 636
rect 3636 634 3638 636
rect 3666 634 3668 636
rect 3696 634 3698 636
rect 3726 634 3728 636
rect 3756 634 3758 636
rect 3842 634 3844 636
rect 3872 634 3874 636
rect 3902 634 3904 636
rect 3932 634 3934 636
rect 3962 634 3964 636
rect 4236 634 4238 636
rect 4266 634 4268 636
rect 4296 634 4298 636
rect 4326 634 4328 636
rect 4356 634 4358 636
rect 4442 634 4444 636
rect 4472 634 4474 636
rect 4502 634 4504 636
rect 4532 634 4534 636
rect 4562 634 4564 636
rect 4592 634 4594 636
rect 4622 634 4624 636
rect 4694 634 4696 636
rect 4724 634 4726 636
rect 4776 634 4778 636
rect 4806 634 4808 636
rect 4836 634 4838 636
rect 4866 634 4868 636
rect 4896 634 4898 636
rect 4926 634 4928 636
rect 4956 634 4958 636
rect 5042 634 5044 636
rect 5072 634 5074 636
rect 5102 634 5104 636
rect 5132 634 5134 636
rect 5162 634 5164 636
rect 5192 634 5194 636
rect 5222 634 5224 636
rect 5294 634 5296 636
rect 5324 634 5326 636
rect 5376 634 5378 636
rect 5406 634 5408 636
rect 5436 634 5438 636
rect 5466 634 5468 636
rect 5496 634 5498 636
rect 5526 634 5528 636
rect 5556 634 5558 636
rect 5642 634 5644 636
rect 5672 634 5674 636
rect 5702 634 5704 636
rect 5732 634 5734 636
rect 5762 634 5764 636
rect 5792 634 5794 636
rect 5822 634 5824 636
rect 5894 634 5896 636
rect 5924 634 5926 636
rect 5976 634 5978 636
rect 6006 634 6008 636
rect 6036 634 6038 636
rect 6066 634 6068 636
rect 6096 634 6098 636
rect 6126 634 6128 636
rect 6156 634 6158 636
rect 6242 634 6244 636
rect 6272 634 6274 636
rect 6302 634 6304 636
rect 6332 634 6334 636
rect 6362 634 6364 636
rect 6636 634 6638 636
rect 6666 634 6668 636
rect 6696 634 6698 636
rect 6726 634 6728 636
rect 6756 634 6758 636
rect 1620 632 1622 634
rect 1820 632 1822 634
rect 1826 632 1828 634
rect 1850 632 1852 634
rect 1856 632 1858 634
rect 1880 632 1882 634
rect 1886 632 1888 634
rect 1910 632 1912 634
rect 1916 632 1918 634
rect 1940 632 1942 634
rect 1946 632 1948 634
rect 1970 632 1972 634
rect 1976 632 1978 634
rect 3234 632 3236 634
rect 3240 632 3242 634
rect 3264 632 3266 634
rect 3270 632 3272 634
rect 3294 632 3296 634
rect 3300 632 3302 634
rect 3324 632 3326 634
rect 3330 632 3332 634
rect 3354 632 3356 634
rect 3360 632 3362 634
rect 3384 632 3386 634
rect 3614 632 3616 634
rect 3638 632 3640 634
rect 3644 632 3646 634
rect 3668 632 3670 634
rect 3674 632 3676 634
rect 3698 632 3700 634
rect 3704 632 3706 634
rect 3728 632 3730 634
rect 3734 632 3736 634
rect 3758 632 3760 634
rect 3764 632 3766 634
rect 3834 632 3836 634
rect 3840 632 3842 634
rect 3864 632 3866 634
rect 3870 632 3872 634
rect 3894 632 3896 634
rect 3900 632 3902 634
rect 3924 632 3926 634
rect 3930 632 3932 634
rect 3954 632 3956 634
rect 3960 632 3962 634
rect 3984 632 3986 634
rect 4214 632 4216 634
rect 4238 632 4240 634
rect 4244 632 4246 634
rect 4268 632 4270 634
rect 4274 632 4276 634
rect 4298 632 4300 634
rect 4304 632 4306 634
rect 4328 632 4330 634
rect 4334 632 4336 634
rect 4358 632 4360 634
rect 4364 632 4366 634
rect 4434 632 4436 634
rect 4440 632 4442 634
rect 4464 632 4466 634
rect 4470 632 4472 634
rect 4494 632 4496 634
rect 4500 632 4502 634
rect 4524 632 4526 634
rect 4530 632 4532 634
rect 4554 632 4556 634
rect 4560 632 4562 634
rect 4584 632 4586 634
rect 4590 632 4592 634
rect 4614 632 4616 634
rect 4620 632 4622 634
rect 4686 632 4688 634
rect 4692 632 4694 634
rect 4716 632 4718 634
rect 4722 632 4724 634
rect 4778 632 4780 634
rect 4784 632 4786 634
rect 4808 632 4810 634
rect 4814 632 4816 634
rect 4838 632 4840 634
rect 4844 632 4846 634
rect 4868 632 4870 634
rect 4874 632 4876 634
rect 4898 632 4900 634
rect 4904 632 4906 634
rect 4928 632 4930 634
rect 4934 632 4936 634
rect 4958 632 4960 634
rect 4964 632 4966 634
rect 5034 632 5036 634
rect 5040 632 5042 634
rect 5064 632 5066 634
rect 5070 632 5072 634
rect 5094 632 5096 634
rect 5100 632 5102 634
rect 5124 632 5126 634
rect 5130 632 5132 634
rect 5154 632 5156 634
rect 5160 632 5162 634
rect 5184 632 5186 634
rect 5190 632 5192 634
rect 5214 632 5216 634
rect 5220 632 5222 634
rect 5286 632 5288 634
rect 5292 632 5294 634
rect 5316 632 5318 634
rect 5322 632 5324 634
rect 5378 632 5380 634
rect 5384 632 5386 634
rect 5408 632 5410 634
rect 5414 632 5416 634
rect 5438 632 5440 634
rect 5444 632 5446 634
rect 5468 632 5470 634
rect 5474 632 5476 634
rect 5498 632 5500 634
rect 5504 632 5506 634
rect 5528 632 5530 634
rect 5534 632 5536 634
rect 5558 632 5560 634
rect 5564 632 5566 634
rect 5634 632 5636 634
rect 5640 632 5642 634
rect 5664 632 5666 634
rect 5670 632 5672 634
rect 5694 632 5696 634
rect 5700 632 5702 634
rect 5724 632 5726 634
rect 5730 632 5732 634
rect 5754 632 5756 634
rect 5760 632 5762 634
rect 5784 632 5786 634
rect 5790 632 5792 634
rect 5814 632 5816 634
rect 5820 632 5822 634
rect 5886 632 5888 634
rect 5892 632 5894 634
rect 5916 632 5918 634
rect 5922 632 5924 634
rect 5978 632 5980 634
rect 5984 632 5986 634
rect 6008 632 6010 634
rect 6014 632 6016 634
rect 6038 632 6040 634
rect 6044 632 6046 634
rect 6068 632 6070 634
rect 6074 632 6076 634
rect 6098 632 6100 634
rect 6104 632 6106 634
rect 6128 632 6130 634
rect 6134 632 6136 634
rect 6158 632 6160 634
rect 6164 632 6166 634
rect 6234 632 6236 634
rect 6240 632 6242 634
rect 6264 632 6266 634
rect 6270 632 6272 634
rect 6294 632 6296 634
rect 6300 632 6302 634
rect 6324 632 6326 634
rect 6330 632 6332 634
rect 6354 632 6356 634
rect 6360 632 6362 634
rect 6384 632 6386 634
rect 6614 632 6616 634
rect 6638 632 6640 634
rect 6644 632 6646 634
rect 6668 632 6670 634
rect 6674 632 6676 634
rect 6698 632 6700 634
rect 6704 632 6706 634
rect 6728 632 6730 634
rect 6734 632 6736 634
rect 6758 632 6760 634
rect 6764 632 6766 634
rect 1818 630 1820 632
rect 1828 630 1830 632
rect 1858 630 1860 632
rect 1888 630 1890 632
rect 1918 630 1920 632
rect 1948 630 1950 632
rect 1978 630 1980 632
rect 3232 630 3234 632
rect 3262 630 3264 632
rect 3292 630 3294 632
rect 3322 630 3324 632
rect 3352 630 3354 632
rect 3382 630 3384 632
rect 3616 630 3618 632
rect 3646 630 3648 632
rect 3676 630 3678 632
rect 3706 630 3708 632
rect 3736 630 3738 632
rect 3766 630 3768 632
rect 3832 630 3834 632
rect 3862 630 3864 632
rect 3892 630 3894 632
rect 3922 630 3924 632
rect 3952 630 3954 632
rect 3982 630 3984 632
rect 4216 630 4218 632
rect 4246 630 4248 632
rect 4276 630 4278 632
rect 4306 630 4308 632
rect 4336 630 4338 632
rect 4366 630 4368 632
rect 4432 630 4434 632
rect 4462 630 4464 632
rect 4492 630 4494 632
rect 4522 630 4524 632
rect 4552 630 4554 632
rect 4582 630 4584 632
rect 4612 630 4614 632
rect 4684 630 4686 632
rect 4714 630 4716 632
rect 4786 630 4788 632
rect 4816 630 4818 632
rect 4846 630 4848 632
rect 4876 630 4878 632
rect 4906 630 4908 632
rect 4936 630 4938 632
rect 4966 630 4968 632
rect 5032 630 5034 632
rect 5062 630 5064 632
rect 5092 630 5094 632
rect 5122 630 5124 632
rect 5152 630 5154 632
rect 5182 630 5184 632
rect 5212 630 5214 632
rect 5284 630 5286 632
rect 5314 630 5316 632
rect 5386 630 5388 632
rect 5416 630 5418 632
rect 5446 630 5448 632
rect 5476 630 5478 632
rect 5506 630 5508 632
rect 5536 630 5538 632
rect 5566 630 5568 632
rect 5632 630 5634 632
rect 5662 630 5664 632
rect 5692 630 5694 632
rect 5722 630 5724 632
rect 5752 630 5754 632
rect 5782 630 5784 632
rect 5812 630 5814 632
rect 5884 630 5886 632
rect 5914 630 5916 632
rect 5986 630 5988 632
rect 6016 630 6018 632
rect 6046 630 6048 632
rect 6076 630 6078 632
rect 6106 630 6108 632
rect 6136 630 6138 632
rect 6166 630 6168 632
rect 6232 630 6234 632
rect 6262 630 6264 632
rect 6292 630 6294 632
rect 6322 630 6324 632
rect 6352 630 6354 632
rect 6382 630 6384 632
rect 6616 630 6618 632
rect 6646 630 6648 632
rect 6676 630 6678 632
rect 6706 630 6708 632
rect 6736 630 6738 632
rect 6766 630 6768 632
rect 1612 624 1614 626
rect 1828 624 1830 626
rect 1858 624 1860 626
rect 1888 624 1890 626
rect 1918 624 1920 626
rect 1948 624 1950 626
rect 1978 624 1980 626
rect 3232 624 3234 626
rect 3262 624 3264 626
rect 3292 624 3294 626
rect 3322 624 3324 626
rect 3352 624 3354 626
rect 3382 624 3384 626
rect 3616 624 3618 626
rect 3646 624 3648 626
rect 3676 624 3678 626
rect 3706 624 3708 626
rect 3736 624 3738 626
rect 3766 624 3768 626
rect 3832 624 3834 626
rect 3862 624 3864 626
rect 3892 624 3894 626
rect 3922 624 3924 626
rect 3952 624 3954 626
rect 3982 624 3984 626
rect 4216 624 4218 626
rect 4246 624 4248 626
rect 4276 624 4278 626
rect 4306 624 4308 626
rect 4336 624 4338 626
rect 4366 624 4368 626
rect 4432 624 4434 626
rect 4462 624 4464 626
rect 4492 624 4494 626
rect 4522 624 4524 626
rect 4552 624 4554 626
rect 4582 624 4584 626
rect 4612 624 4614 626
rect 4684 624 4686 626
rect 4714 624 4716 626
rect 4786 624 4788 626
rect 4816 624 4818 626
rect 4846 624 4848 626
rect 4876 624 4878 626
rect 4906 624 4908 626
rect 4936 624 4938 626
rect 4966 624 4968 626
rect 5032 624 5034 626
rect 5062 624 5064 626
rect 5092 624 5094 626
rect 5122 624 5124 626
rect 5152 624 5154 626
rect 5182 624 5184 626
rect 5212 624 5214 626
rect 5284 624 5286 626
rect 5314 624 5316 626
rect 5386 624 5388 626
rect 5416 624 5418 626
rect 5446 624 5448 626
rect 5476 624 5478 626
rect 5506 624 5508 626
rect 5536 624 5538 626
rect 5566 624 5568 626
rect 5632 624 5634 626
rect 5662 624 5664 626
rect 5692 624 5694 626
rect 5722 624 5724 626
rect 5752 624 5754 626
rect 5782 624 5784 626
rect 5812 624 5814 626
rect 5884 624 5886 626
rect 5914 624 5916 626
rect 5986 624 5988 626
rect 6016 624 6018 626
rect 6046 624 6048 626
rect 6076 624 6078 626
rect 6106 624 6108 626
rect 6136 624 6138 626
rect 6166 624 6168 626
rect 6232 624 6234 626
rect 6262 624 6264 626
rect 6292 624 6294 626
rect 6322 624 6324 626
rect 6352 624 6354 626
rect 6382 624 6384 626
rect 6616 624 6618 626
rect 6646 624 6648 626
rect 6676 624 6678 626
rect 6706 624 6708 626
rect 6736 624 6738 626
rect 6766 624 6768 626
rect 1610 622 1612 624
rect 1810 622 1812 624
rect 1826 622 1828 624
rect 1850 622 1852 624
rect 1856 622 1858 624
rect 1880 622 1882 624
rect 1886 622 1888 624
rect 1910 622 1912 624
rect 1916 622 1918 624
rect 1940 622 1942 624
rect 1946 622 1948 624
rect 1970 622 1972 624
rect 1976 622 1978 624
rect 3234 622 3236 624
rect 3240 622 3242 624
rect 3264 622 3266 624
rect 3270 622 3272 624
rect 3294 622 3296 624
rect 3300 622 3302 624
rect 3324 622 3326 624
rect 3330 622 3332 624
rect 3354 622 3356 624
rect 3360 622 3362 624
rect 3384 622 3386 624
rect 3614 622 3616 624
rect 3638 622 3640 624
rect 3644 622 3646 624
rect 3668 622 3670 624
rect 3674 622 3676 624
rect 3698 622 3700 624
rect 3704 622 3706 624
rect 3728 622 3730 624
rect 3734 622 3736 624
rect 3758 622 3760 624
rect 3764 622 3766 624
rect 3834 622 3836 624
rect 3840 622 3842 624
rect 3864 622 3866 624
rect 3870 622 3872 624
rect 3894 622 3896 624
rect 3900 622 3902 624
rect 3924 622 3926 624
rect 3930 622 3932 624
rect 3954 622 3956 624
rect 3960 622 3962 624
rect 3984 622 3986 624
rect 4214 622 4216 624
rect 4238 622 4240 624
rect 4244 622 4246 624
rect 4268 622 4270 624
rect 4274 622 4276 624
rect 4298 622 4300 624
rect 4304 622 4306 624
rect 4328 622 4330 624
rect 4334 622 4336 624
rect 4358 622 4360 624
rect 4364 622 4366 624
rect 4434 622 4436 624
rect 4440 622 4442 624
rect 4464 622 4466 624
rect 4470 622 4472 624
rect 4494 622 4496 624
rect 4500 622 4502 624
rect 4524 622 4526 624
rect 4530 622 4532 624
rect 4554 622 4556 624
rect 4560 622 4562 624
rect 4584 622 4586 624
rect 4590 622 4592 624
rect 4614 622 4616 624
rect 4620 622 4622 624
rect 4686 622 4688 624
rect 4692 622 4694 624
rect 4716 622 4718 624
rect 4722 622 4724 624
rect 4778 622 4780 624
rect 4784 622 4786 624
rect 4808 622 4810 624
rect 4814 622 4816 624
rect 4838 622 4840 624
rect 4844 622 4846 624
rect 4868 622 4870 624
rect 4874 622 4876 624
rect 4898 622 4900 624
rect 4904 622 4906 624
rect 4928 622 4930 624
rect 4934 622 4936 624
rect 4958 622 4960 624
rect 4964 622 4966 624
rect 5034 622 5036 624
rect 5040 622 5042 624
rect 5064 622 5066 624
rect 5070 622 5072 624
rect 5094 622 5096 624
rect 5100 622 5102 624
rect 5124 622 5126 624
rect 5130 622 5132 624
rect 5154 622 5156 624
rect 5160 622 5162 624
rect 5184 622 5186 624
rect 5190 622 5192 624
rect 5214 622 5216 624
rect 5220 622 5222 624
rect 5286 622 5288 624
rect 5292 622 5294 624
rect 5316 622 5318 624
rect 5322 622 5324 624
rect 5378 622 5380 624
rect 5384 622 5386 624
rect 5408 622 5410 624
rect 5414 622 5416 624
rect 5438 622 5440 624
rect 5444 622 5446 624
rect 5468 622 5470 624
rect 5474 622 5476 624
rect 5498 622 5500 624
rect 5504 622 5506 624
rect 5528 622 5530 624
rect 5534 622 5536 624
rect 5558 622 5560 624
rect 5564 622 5566 624
rect 5634 622 5636 624
rect 5640 622 5642 624
rect 5664 622 5666 624
rect 5670 622 5672 624
rect 5694 622 5696 624
rect 5700 622 5702 624
rect 5724 622 5726 624
rect 5730 622 5732 624
rect 5754 622 5756 624
rect 5760 622 5762 624
rect 5784 622 5786 624
rect 5790 622 5792 624
rect 5814 622 5816 624
rect 5820 622 5822 624
rect 5886 622 5888 624
rect 5892 622 5894 624
rect 5916 622 5918 624
rect 5922 622 5924 624
rect 5978 622 5980 624
rect 5984 622 5986 624
rect 6008 622 6010 624
rect 6014 622 6016 624
rect 6038 622 6040 624
rect 6044 622 6046 624
rect 6068 622 6070 624
rect 6074 622 6076 624
rect 6098 622 6100 624
rect 6104 622 6106 624
rect 6128 622 6130 624
rect 6134 622 6136 624
rect 6158 622 6160 624
rect 6164 622 6166 624
rect 6234 622 6236 624
rect 6240 622 6242 624
rect 6264 622 6266 624
rect 6270 622 6272 624
rect 6294 622 6296 624
rect 6300 622 6302 624
rect 6324 622 6326 624
rect 6330 622 6332 624
rect 6354 622 6356 624
rect 6360 622 6362 624
rect 6384 622 6386 624
rect 6614 622 6616 624
rect 6638 622 6640 624
rect 6644 622 6646 624
rect 6668 622 6670 624
rect 6674 622 6676 624
rect 6698 622 6700 624
rect 6704 622 6706 624
rect 6728 622 6730 624
rect 6734 622 6736 624
rect 6758 622 6760 624
rect 6764 622 6766 624
rect 1808 620 1810 622
rect 1848 620 1850 622
rect 1878 620 1880 622
rect 1908 620 1910 622
rect 1938 620 1940 622
rect 1968 620 1970 622
rect 3242 620 3244 622
rect 3272 620 3274 622
rect 3302 620 3304 622
rect 3332 620 3334 622
rect 3362 620 3364 622
rect 3636 620 3638 622
rect 3666 620 3668 622
rect 3696 620 3698 622
rect 3726 620 3728 622
rect 3756 620 3758 622
rect 3842 620 3844 622
rect 3872 620 3874 622
rect 3902 620 3904 622
rect 3932 620 3934 622
rect 3962 620 3964 622
rect 4236 620 4238 622
rect 4266 620 4268 622
rect 4296 620 4298 622
rect 4326 620 4328 622
rect 4356 620 4358 622
rect 4442 620 4444 622
rect 4472 620 4474 622
rect 4502 620 4504 622
rect 4532 620 4534 622
rect 4562 620 4564 622
rect 4592 620 4594 622
rect 4622 620 4624 622
rect 4694 620 4696 622
rect 4724 620 4726 622
rect 4776 620 4778 622
rect 4806 620 4808 622
rect 4836 620 4838 622
rect 4866 620 4868 622
rect 4896 620 4898 622
rect 4926 620 4928 622
rect 4956 620 4958 622
rect 5042 620 5044 622
rect 5072 620 5074 622
rect 5102 620 5104 622
rect 5132 620 5134 622
rect 5162 620 5164 622
rect 5192 620 5194 622
rect 5222 620 5224 622
rect 5294 620 5296 622
rect 5324 620 5326 622
rect 5376 620 5378 622
rect 5406 620 5408 622
rect 5436 620 5438 622
rect 5466 620 5468 622
rect 5496 620 5498 622
rect 5526 620 5528 622
rect 5556 620 5558 622
rect 5642 620 5644 622
rect 5672 620 5674 622
rect 5702 620 5704 622
rect 5732 620 5734 622
rect 5762 620 5764 622
rect 5792 620 5794 622
rect 5822 620 5824 622
rect 5894 620 5896 622
rect 5924 620 5926 622
rect 5976 620 5978 622
rect 6006 620 6008 622
rect 6036 620 6038 622
rect 6066 620 6068 622
rect 6096 620 6098 622
rect 6126 620 6128 622
rect 6156 620 6158 622
rect 6242 620 6244 622
rect 6272 620 6274 622
rect 6302 620 6304 622
rect 6332 620 6334 622
rect 6362 620 6364 622
rect 6636 620 6638 622
rect 6666 620 6668 622
rect 6696 620 6698 622
rect 6726 620 6728 622
rect 6756 620 6758 622
rect 1602 614 1604 616
rect 1808 614 1810 616
rect 1818 614 1820 616
rect 1848 614 1850 616
rect 1878 614 1880 616
rect 1908 614 1910 616
rect 1938 614 1940 616
rect 1968 614 1970 616
rect 4622 614 4624 616
rect 4694 614 4696 616
rect 4724 614 4726 616
rect 4776 614 4778 616
rect 5222 614 5224 616
rect 5294 614 5296 616
rect 5324 614 5326 616
rect 5376 614 5378 616
rect 5822 614 5824 616
rect 5894 614 5896 616
rect 5924 614 5926 616
rect 5976 614 5978 616
rect 1600 612 1602 614
rect 1800 612 1802 614
rect 1806 612 1808 614
rect 1820 612 1822 614
rect 1826 612 1828 614
rect 1850 612 1852 614
rect 1856 612 1858 614
rect 1880 612 1882 614
rect 1886 612 1888 614
rect 1910 612 1912 614
rect 1916 612 1918 614
rect 1940 612 1942 614
rect 1946 612 1948 614
rect 1970 612 1972 614
rect 1976 612 1978 614
rect 4620 612 4622 614
rect 4686 612 4688 614
rect 4692 612 4694 614
rect 4716 612 4718 614
rect 4722 612 4724 614
rect 4778 612 4780 614
rect 5220 612 5222 614
rect 5286 612 5288 614
rect 5292 612 5294 614
rect 5316 612 5318 614
rect 5322 612 5324 614
rect 5378 612 5380 614
rect 5820 612 5822 614
rect 5886 612 5888 614
rect 5892 612 5894 614
rect 5916 612 5918 614
rect 5922 612 5924 614
rect 5978 612 5980 614
rect 1798 610 1800 612
rect 1828 610 1830 612
rect 1858 610 1860 612
rect 1888 610 1890 612
rect 1918 610 1920 612
rect 1948 610 1950 612
rect 1978 610 1980 612
rect 4684 610 4686 612
rect 4714 610 4716 612
rect 5284 610 5286 612
rect 5314 610 5316 612
rect 5884 610 5886 612
rect 5914 610 5916 612
rect 1798 604 1800 606
rect 1828 604 1830 606
rect 1858 604 1860 606
rect 1888 604 1890 606
rect 1918 604 1920 606
rect 1948 604 1950 606
rect 1978 604 1980 606
rect 4684 604 4686 606
rect 4714 604 4716 606
rect 5284 604 5286 606
rect 5314 604 5316 606
rect 5884 604 5886 606
rect 5914 604 5916 606
rect 1790 602 1792 604
rect 1796 602 1798 604
rect 1820 602 1822 604
rect 1826 602 1828 604
rect 1850 602 1852 604
rect 1856 602 1858 604
rect 1880 602 1882 604
rect 1886 602 1888 604
rect 1910 602 1912 604
rect 1916 602 1918 604
rect 1940 602 1942 604
rect 1946 602 1948 604
rect 1970 602 1972 604
rect 1976 602 1978 604
rect 4620 602 4622 604
rect 4686 602 4688 604
rect 4692 602 4694 604
rect 4716 602 4718 604
rect 4722 602 4724 604
rect 4778 602 4780 604
rect 5220 602 5222 604
rect 5286 602 5288 604
rect 5292 602 5294 604
rect 5316 602 5318 604
rect 5322 602 5324 604
rect 5378 602 5380 604
rect 5820 602 5822 604
rect 5886 602 5888 604
rect 5892 602 5894 604
rect 5916 602 5918 604
rect 5922 602 5924 604
rect 5978 602 5980 604
rect 1788 600 1790 602
rect 1818 600 1820 602
rect 1848 600 1850 602
rect 1878 600 1880 602
rect 1908 600 1910 602
rect 1938 600 1940 602
rect 1968 600 1970 602
rect 4622 600 4624 602
rect 4694 600 4696 602
rect 4724 600 4726 602
rect 4776 600 4778 602
rect 5222 600 5224 602
rect 5294 600 5296 602
rect 5324 600 5326 602
rect 5376 600 5378 602
rect 5822 600 5824 602
rect 5894 600 5896 602
rect 5924 600 5926 602
rect 5976 600 5978 602
rect 1788 594 1790 596
rect 1848 594 1850 596
rect 1878 594 1880 596
rect 1908 594 1910 596
rect 1938 594 1940 596
rect 1968 594 1970 596
rect 3242 594 3244 596
rect 3272 594 3274 596
rect 3302 594 3304 596
rect 3332 594 3334 596
rect 3362 594 3364 596
rect 3636 594 3638 596
rect 3666 594 3668 596
rect 3696 594 3698 596
rect 3726 594 3728 596
rect 3756 594 3758 596
rect 3842 594 3844 596
rect 3872 594 3874 596
rect 3902 594 3904 596
rect 3932 594 3934 596
rect 3962 594 3964 596
rect 4236 594 4238 596
rect 4266 594 4268 596
rect 4296 594 4298 596
rect 4326 594 4328 596
rect 4356 594 4358 596
rect 4442 594 4444 596
rect 4472 594 4474 596
rect 4502 594 4504 596
rect 4532 594 4534 596
rect 4562 594 4564 596
rect 4592 594 4594 596
rect 4622 594 4624 596
rect 4776 594 4778 596
rect 4806 594 4808 596
rect 4836 594 4838 596
rect 4866 594 4868 596
rect 4896 594 4898 596
rect 4926 594 4928 596
rect 4956 594 4958 596
rect 5042 594 5044 596
rect 5072 594 5074 596
rect 5102 594 5104 596
rect 5132 594 5134 596
rect 5162 594 5164 596
rect 5192 594 5194 596
rect 5222 594 5224 596
rect 5376 594 5378 596
rect 5406 594 5408 596
rect 5436 594 5438 596
rect 5466 594 5468 596
rect 5496 594 5498 596
rect 5526 594 5528 596
rect 5556 594 5558 596
rect 5642 594 5644 596
rect 5672 594 5674 596
rect 5702 594 5704 596
rect 5732 594 5734 596
rect 5762 594 5764 596
rect 5792 594 5794 596
rect 5822 594 5824 596
rect 5976 594 5978 596
rect 6006 594 6008 596
rect 6036 594 6038 596
rect 6066 594 6068 596
rect 6096 594 6098 596
rect 6126 594 6128 596
rect 6156 594 6158 596
rect 6242 594 6244 596
rect 6272 594 6274 596
rect 6302 594 6304 596
rect 6332 594 6334 596
rect 6362 594 6364 596
rect 6636 594 6638 596
rect 6666 594 6668 596
rect 6696 594 6698 596
rect 6726 594 6728 596
rect 6756 594 6758 596
rect 1780 592 1782 594
rect 1786 592 1788 594
rect 1810 592 1812 594
rect 1826 592 1828 594
rect 1850 592 1852 594
rect 1856 592 1858 594
rect 1880 592 1882 594
rect 1886 592 1888 594
rect 1910 592 1912 594
rect 1916 592 1918 594
rect 1940 592 1942 594
rect 1946 592 1948 594
rect 1970 592 1972 594
rect 1976 592 1978 594
rect 3234 592 3236 594
rect 3240 592 3242 594
rect 3264 592 3266 594
rect 3270 592 3272 594
rect 3294 592 3296 594
rect 3300 592 3302 594
rect 3324 592 3326 594
rect 3330 592 3332 594
rect 3354 592 3356 594
rect 3360 592 3362 594
rect 3384 592 3386 594
rect 3614 592 3616 594
rect 3638 592 3640 594
rect 3644 592 3646 594
rect 3668 592 3670 594
rect 3674 592 3676 594
rect 3698 592 3700 594
rect 3704 592 3706 594
rect 3728 592 3730 594
rect 3734 592 3736 594
rect 3758 592 3760 594
rect 3764 592 3766 594
rect 3834 592 3836 594
rect 3840 592 3842 594
rect 3864 592 3866 594
rect 3870 592 3872 594
rect 3894 592 3896 594
rect 3900 592 3902 594
rect 3924 592 3926 594
rect 3930 592 3932 594
rect 3954 592 3956 594
rect 3960 592 3962 594
rect 3984 592 3986 594
rect 4214 592 4216 594
rect 4238 592 4240 594
rect 4244 592 4246 594
rect 4268 592 4270 594
rect 4274 592 4276 594
rect 4298 592 4300 594
rect 4304 592 4306 594
rect 4328 592 4330 594
rect 4334 592 4336 594
rect 4358 592 4360 594
rect 4364 592 4366 594
rect 4434 592 4436 594
rect 4440 592 4442 594
rect 4464 592 4466 594
rect 4470 592 4472 594
rect 4494 592 4496 594
rect 4500 592 4502 594
rect 4524 592 4526 594
rect 4530 592 4532 594
rect 4554 592 4556 594
rect 4560 592 4562 594
rect 4584 592 4586 594
rect 4590 592 4592 594
rect 4614 592 4616 594
rect 4620 592 4622 594
rect 4666 592 4668 594
rect 4672 592 4674 594
rect 4686 592 4688 594
rect 4702 592 4704 594
rect 4716 592 4718 594
rect 4732 592 4734 594
rect 4778 592 4780 594
rect 4784 592 4786 594
rect 4808 592 4810 594
rect 4814 592 4816 594
rect 4838 592 4840 594
rect 4844 592 4846 594
rect 4868 592 4870 594
rect 4874 592 4876 594
rect 4898 592 4900 594
rect 4904 592 4906 594
rect 4928 592 4930 594
rect 4934 592 4936 594
rect 4958 592 4960 594
rect 4964 592 4966 594
rect 5034 592 5036 594
rect 5040 592 5042 594
rect 5064 592 5066 594
rect 5070 592 5072 594
rect 5094 592 5096 594
rect 5100 592 5102 594
rect 5124 592 5126 594
rect 5130 592 5132 594
rect 5154 592 5156 594
rect 5160 592 5162 594
rect 5184 592 5186 594
rect 5190 592 5192 594
rect 5214 592 5216 594
rect 5220 592 5222 594
rect 5266 592 5268 594
rect 5272 592 5274 594
rect 5286 592 5288 594
rect 5302 592 5304 594
rect 5316 592 5318 594
rect 5332 592 5334 594
rect 5378 592 5380 594
rect 5384 592 5386 594
rect 5408 592 5410 594
rect 5414 592 5416 594
rect 5438 592 5440 594
rect 5444 592 5446 594
rect 5468 592 5470 594
rect 5474 592 5476 594
rect 5498 592 5500 594
rect 5504 592 5506 594
rect 5528 592 5530 594
rect 5534 592 5536 594
rect 5558 592 5560 594
rect 5564 592 5566 594
rect 5634 592 5636 594
rect 5640 592 5642 594
rect 5664 592 5666 594
rect 5670 592 5672 594
rect 5694 592 5696 594
rect 5700 592 5702 594
rect 5724 592 5726 594
rect 5730 592 5732 594
rect 5754 592 5756 594
rect 5760 592 5762 594
rect 5784 592 5786 594
rect 5790 592 5792 594
rect 5814 592 5816 594
rect 5820 592 5822 594
rect 5866 592 5868 594
rect 5872 592 5874 594
rect 5886 592 5888 594
rect 5902 592 5904 594
rect 5916 592 5918 594
rect 5932 592 5934 594
rect 5978 592 5980 594
rect 5984 592 5986 594
rect 6008 592 6010 594
rect 6014 592 6016 594
rect 6038 592 6040 594
rect 6044 592 6046 594
rect 6068 592 6070 594
rect 6074 592 6076 594
rect 6098 592 6100 594
rect 6104 592 6106 594
rect 6128 592 6130 594
rect 6134 592 6136 594
rect 6158 592 6160 594
rect 6164 592 6166 594
rect 6234 592 6236 594
rect 6240 592 6242 594
rect 6264 592 6266 594
rect 6270 592 6272 594
rect 6294 592 6296 594
rect 6300 592 6302 594
rect 6324 592 6326 594
rect 6330 592 6332 594
rect 6354 592 6356 594
rect 6360 592 6362 594
rect 6384 592 6386 594
rect 6614 592 6616 594
rect 6638 592 6640 594
rect 6644 592 6646 594
rect 6668 592 6670 594
rect 6674 592 6676 594
rect 6698 592 6700 594
rect 6704 592 6706 594
rect 6728 592 6730 594
rect 6734 592 6736 594
rect 6758 592 6760 594
rect 6764 592 6766 594
rect 1778 590 1780 592
rect 1808 590 1810 592
rect 1828 590 1830 592
rect 1858 590 1860 592
rect 1888 590 1890 592
rect 1918 590 1920 592
rect 1948 590 1950 592
rect 1978 590 1980 592
rect 3232 590 3234 592
rect 3262 590 3264 592
rect 3292 590 3294 592
rect 3322 590 3324 592
rect 3352 590 3354 592
rect 3382 590 3384 592
rect 3616 590 3618 592
rect 3646 590 3648 592
rect 3676 590 3678 592
rect 3706 590 3708 592
rect 3736 590 3738 592
rect 3766 590 3768 592
rect 3832 590 3834 592
rect 3862 590 3864 592
rect 3892 590 3894 592
rect 3922 590 3924 592
rect 3952 590 3954 592
rect 3982 590 3984 592
rect 4216 590 4218 592
rect 4246 590 4248 592
rect 4276 590 4278 592
rect 4306 590 4308 592
rect 4336 590 4338 592
rect 4366 590 4368 592
rect 4432 590 4434 592
rect 4462 590 4464 592
rect 4492 590 4494 592
rect 4522 590 4524 592
rect 4552 590 4554 592
rect 4582 590 4584 592
rect 4612 590 4614 592
rect 4664 590 4666 592
rect 4674 590 4676 592
rect 4684 590 4686 592
rect 4704 590 4706 592
rect 4714 590 4716 592
rect 4734 590 4736 592
rect 4786 590 4788 592
rect 4816 590 4818 592
rect 4846 590 4848 592
rect 4876 590 4878 592
rect 4906 590 4908 592
rect 4936 590 4938 592
rect 4966 590 4968 592
rect 5032 590 5034 592
rect 5062 590 5064 592
rect 5092 590 5094 592
rect 5122 590 5124 592
rect 5152 590 5154 592
rect 5182 590 5184 592
rect 5212 590 5214 592
rect 5264 590 5266 592
rect 5274 590 5276 592
rect 5284 590 5286 592
rect 5304 590 5306 592
rect 5314 590 5316 592
rect 5334 590 5336 592
rect 5386 590 5388 592
rect 5416 590 5418 592
rect 5446 590 5448 592
rect 5476 590 5478 592
rect 5506 590 5508 592
rect 5536 590 5538 592
rect 5566 590 5568 592
rect 5632 590 5634 592
rect 5662 590 5664 592
rect 5692 590 5694 592
rect 5722 590 5724 592
rect 5752 590 5754 592
rect 5782 590 5784 592
rect 5812 590 5814 592
rect 5864 590 5866 592
rect 5874 590 5876 592
rect 5884 590 5886 592
rect 5904 590 5906 592
rect 5914 590 5916 592
rect 5934 590 5936 592
rect 5986 590 5988 592
rect 6016 590 6018 592
rect 6046 590 6048 592
rect 6076 590 6078 592
rect 6106 590 6108 592
rect 6136 590 6138 592
rect 6166 590 6168 592
rect 6232 590 6234 592
rect 6262 590 6264 592
rect 6292 590 6294 592
rect 6322 590 6324 592
rect 6352 590 6354 592
rect 6382 590 6384 592
rect 6616 590 6618 592
rect 6646 590 6648 592
rect 6676 590 6678 592
rect 6706 590 6708 592
rect 6736 590 6738 592
rect 6766 590 6768 592
rect 1778 584 1780 586
rect 1808 584 1810 586
rect 1818 584 1820 586
rect 1828 584 1830 586
rect 1888 584 1890 586
rect 1918 584 1920 586
rect 1948 584 1950 586
rect 1978 584 1980 586
rect 3232 584 3234 586
rect 3262 584 3264 586
rect 3292 584 3294 586
rect 3706 584 3708 586
rect 3736 584 3738 586
rect 3766 584 3768 586
rect 3832 584 3834 586
rect 3862 584 3864 586
rect 3892 584 3894 586
rect 4306 584 4308 586
rect 4336 584 4338 586
rect 4366 584 4368 586
rect 4432 584 4434 586
rect 4462 584 4464 586
rect 4492 584 4494 586
rect 4906 584 4908 586
rect 4936 584 4938 586
rect 4966 584 4968 586
rect 5032 584 5034 586
rect 5062 584 5064 586
rect 5092 584 5094 586
rect 5506 584 5508 586
rect 5536 584 5538 586
rect 5566 584 5568 586
rect 5632 584 5634 586
rect 5662 584 5664 586
rect 5692 584 5694 586
rect 6106 584 6108 586
rect 6136 584 6138 586
rect 6166 584 6168 586
rect 6232 584 6234 586
rect 6262 584 6264 586
rect 6292 584 6294 586
rect 6706 584 6708 586
rect 6736 584 6738 586
rect 6766 584 6768 586
rect 1770 582 1772 584
rect 1776 582 1778 584
rect 1800 582 1802 584
rect 1806 582 1808 584
rect 1820 582 1822 584
rect 1826 582 1828 584
rect 1850 582 1852 584
rect 1866 582 1868 584
rect 1880 582 1882 584
rect 1886 582 1888 584
rect 1910 582 1912 584
rect 1916 582 1918 584
rect 1940 582 1942 584
rect 1946 582 1948 584
rect 1970 582 1972 584
rect 1976 582 1978 584
rect 3234 582 3236 584
rect 3240 582 3242 584
rect 3264 582 3266 584
rect 3270 582 3272 584
rect 3294 582 3296 584
rect 3300 582 3302 584
rect 3314 582 3316 584
rect 3330 582 3332 584
rect 3344 582 3346 584
rect 3360 582 3362 584
rect 3374 582 3376 584
rect 3624 582 3626 584
rect 3638 582 3640 584
rect 3654 582 3656 584
rect 3668 582 3670 584
rect 3684 582 3686 584
rect 3698 582 3700 584
rect 3704 582 3706 584
rect 3728 582 3730 584
rect 3734 582 3736 584
rect 3758 582 3760 584
rect 3764 582 3766 584
rect 3834 582 3836 584
rect 3840 582 3842 584
rect 3864 582 3866 584
rect 3870 582 3872 584
rect 3894 582 3896 584
rect 3900 582 3902 584
rect 3914 582 3916 584
rect 3930 582 3932 584
rect 3944 582 3946 584
rect 3960 582 3962 584
rect 3974 582 3976 584
rect 4224 582 4226 584
rect 4238 582 4240 584
rect 4254 582 4256 584
rect 4268 582 4270 584
rect 4284 582 4286 584
rect 4298 582 4300 584
rect 4304 582 4306 584
rect 4328 582 4330 584
rect 4334 582 4336 584
rect 4358 582 4360 584
rect 4364 582 4366 584
rect 4434 582 4436 584
rect 4440 582 4442 584
rect 4464 582 4466 584
rect 4470 582 4472 584
rect 4494 582 4496 584
rect 4500 582 4502 584
rect 4514 582 4516 584
rect 4530 582 4532 584
rect 4544 582 4546 584
rect 4560 582 4562 584
rect 4574 582 4576 584
rect 4590 582 4592 584
rect 4604 582 4606 584
rect 4620 582 4622 584
rect 4634 582 4636 584
rect 4640 582 4642 584
rect 4758 582 4760 584
rect 4764 582 4766 584
rect 4778 582 4780 584
rect 4794 582 4796 584
rect 4808 582 4810 584
rect 4824 582 4826 584
rect 4838 582 4840 584
rect 4854 582 4856 584
rect 4868 582 4870 584
rect 4884 582 4886 584
rect 4898 582 4900 584
rect 4904 582 4906 584
rect 4928 582 4930 584
rect 4934 582 4936 584
rect 4958 582 4960 584
rect 4964 582 4966 584
rect 5034 582 5036 584
rect 5040 582 5042 584
rect 5064 582 5066 584
rect 5070 582 5072 584
rect 5094 582 5096 584
rect 5100 582 5102 584
rect 5114 582 5116 584
rect 5130 582 5132 584
rect 5144 582 5146 584
rect 5160 582 5162 584
rect 5174 582 5176 584
rect 5190 582 5192 584
rect 5204 582 5206 584
rect 5220 582 5222 584
rect 5234 582 5236 584
rect 5240 582 5242 584
rect 5358 582 5360 584
rect 5364 582 5366 584
rect 5378 582 5380 584
rect 5394 582 5396 584
rect 5408 582 5410 584
rect 5424 582 5426 584
rect 5438 582 5440 584
rect 5454 582 5456 584
rect 5468 582 5470 584
rect 5484 582 5486 584
rect 5498 582 5500 584
rect 5504 582 5506 584
rect 5528 582 5530 584
rect 5534 582 5536 584
rect 5558 582 5560 584
rect 5564 582 5566 584
rect 5634 582 5636 584
rect 5640 582 5642 584
rect 5664 582 5666 584
rect 5670 582 5672 584
rect 5694 582 5696 584
rect 5700 582 5702 584
rect 5714 582 5716 584
rect 5730 582 5732 584
rect 5744 582 5746 584
rect 5760 582 5762 584
rect 5774 582 5776 584
rect 5790 582 5792 584
rect 5804 582 5806 584
rect 5820 582 5822 584
rect 5834 582 5836 584
rect 5840 582 5842 584
rect 5958 582 5960 584
rect 5964 582 5966 584
rect 5978 582 5980 584
rect 5994 582 5996 584
rect 6008 582 6010 584
rect 6024 582 6026 584
rect 6038 582 6040 584
rect 6054 582 6056 584
rect 6068 582 6070 584
rect 6084 582 6086 584
rect 6098 582 6100 584
rect 6104 582 6106 584
rect 6128 582 6130 584
rect 6134 582 6136 584
rect 6158 582 6160 584
rect 6164 582 6166 584
rect 6234 582 6236 584
rect 6240 582 6242 584
rect 6264 582 6266 584
rect 6270 582 6272 584
rect 6294 582 6296 584
rect 6300 582 6302 584
rect 6314 582 6316 584
rect 6330 582 6332 584
rect 6344 582 6346 584
rect 6360 582 6362 584
rect 6374 582 6376 584
rect 6624 582 6626 584
rect 6638 582 6640 584
rect 6654 582 6656 584
rect 6668 582 6670 584
rect 6684 582 6686 584
rect 6698 582 6700 584
rect 6704 582 6706 584
rect 6728 582 6730 584
rect 6734 582 6736 584
rect 6758 582 6760 584
rect 6764 582 6766 584
rect 1768 580 1770 582
rect 1798 580 1800 582
rect 1848 580 1850 582
rect 1868 580 1870 582
rect 1878 580 1880 582
rect 1908 580 1910 582
rect 1938 580 1940 582
rect 1968 580 1970 582
rect 3242 580 3244 582
rect 3272 580 3274 582
rect 3302 580 3304 582
rect 3312 580 3314 582
rect 3332 580 3334 582
rect 3342 580 3344 582
rect 3362 580 3364 582
rect 3372 580 3374 582
rect 3626 580 3628 582
rect 3636 580 3638 582
rect 3656 580 3658 582
rect 3666 580 3668 582
rect 3686 580 3688 582
rect 3696 580 3698 582
rect 3726 580 3728 582
rect 3756 580 3758 582
rect 3842 580 3844 582
rect 3872 580 3874 582
rect 3902 580 3904 582
rect 3912 580 3914 582
rect 3932 580 3934 582
rect 3942 580 3944 582
rect 3962 580 3964 582
rect 3972 580 3974 582
rect 4226 580 4228 582
rect 4236 580 4238 582
rect 4256 580 4258 582
rect 4266 580 4268 582
rect 4286 580 4288 582
rect 4296 580 4298 582
rect 4326 580 4328 582
rect 4356 580 4358 582
rect 4442 580 4444 582
rect 4472 580 4474 582
rect 4502 580 4504 582
rect 4512 580 4514 582
rect 4532 580 4534 582
rect 4542 580 4544 582
rect 4562 580 4564 582
rect 4572 580 4574 582
rect 4592 580 4594 582
rect 4602 580 4604 582
rect 4622 580 4624 582
rect 4632 580 4634 582
rect 4642 580 4644 582
rect 4756 580 4758 582
rect 4766 580 4768 582
rect 4776 580 4778 582
rect 4796 580 4798 582
rect 4806 580 4808 582
rect 4826 580 4828 582
rect 4836 580 4838 582
rect 4856 580 4858 582
rect 4866 580 4868 582
rect 4886 580 4888 582
rect 4896 580 4898 582
rect 4926 580 4928 582
rect 4956 580 4958 582
rect 5042 580 5044 582
rect 5072 580 5074 582
rect 5102 580 5104 582
rect 5112 580 5114 582
rect 5132 580 5134 582
rect 5142 580 5144 582
rect 5162 580 5164 582
rect 5172 580 5174 582
rect 5192 580 5194 582
rect 5202 580 5204 582
rect 5222 580 5224 582
rect 5232 580 5234 582
rect 5242 580 5244 582
rect 5356 580 5358 582
rect 5366 580 5368 582
rect 5376 580 5378 582
rect 5396 580 5398 582
rect 5406 580 5408 582
rect 5426 580 5428 582
rect 5436 580 5438 582
rect 5456 580 5458 582
rect 5466 580 5468 582
rect 5486 580 5488 582
rect 5496 580 5498 582
rect 5526 580 5528 582
rect 5556 580 5558 582
rect 5642 580 5644 582
rect 5672 580 5674 582
rect 5702 580 5704 582
rect 5712 580 5714 582
rect 5732 580 5734 582
rect 5742 580 5744 582
rect 5762 580 5764 582
rect 5772 580 5774 582
rect 5792 580 5794 582
rect 5802 580 5804 582
rect 5822 580 5824 582
rect 5832 580 5834 582
rect 5842 580 5844 582
rect 5956 580 5958 582
rect 5966 580 5968 582
rect 5976 580 5978 582
rect 5996 580 5998 582
rect 6006 580 6008 582
rect 6026 580 6028 582
rect 6036 580 6038 582
rect 6056 580 6058 582
rect 6066 580 6068 582
rect 6086 580 6088 582
rect 6096 580 6098 582
rect 6126 580 6128 582
rect 6156 580 6158 582
rect 6242 580 6244 582
rect 6272 580 6274 582
rect 6302 580 6304 582
rect 6312 580 6314 582
rect 6332 580 6334 582
rect 6342 580 6344 582
rect 6362 580 6364 582
rect 6372 580 6374 582
rect 6626 580 6628 582
rect 6636 580 6638 582
rect 6656 580 6658 582
rect 6666 580 6668 582
rect 6686 580 6688 582
rect 6696 580 6698 582
rect 6726 580 6728 582
rect 6756 580 6758 582
rect 1768 574 1770 576
rect 1798 574 1800 576
rect 1868 574 1870 576
rect 1878 574 1880 576
rect 1908 574 1910 576
rect 1938 574 1940 576
rect 1968 574 1970 576
rect 3242 574 3244 576
rect 3272 574 3274 576
rect 3302 574 3304 576
rect 3312 574 3314 576
rect 3332 574 3334 576
rect 3342 574 3344 576
rect 3362 574 3364 576
rect 3372 574 3374 576
rect 3626 574 3628 576
rect 3636 574 3638 576
rect 3656 574 3658 576
rect 3666 574 3668 576
rect 3686 574 3688 576
rect 3696 574 3698 576
rect 3726 574 3728 576
rect 3756 574 3758 576
rect 3842 574 3844 576
rect 3872 574 3874 576
rect 3902 574 3904 576
rect 3912 574 3914 576
rect 3932 574 3934 576
rect 3942 574 3944 576
rect 3962 574 3964 576
rect 3972 574 3974 576
rect 4226 574 4228 576
rect 4236 574 4238 576
rect 4256 574 4258 576
rect 4266 574 4268 576
rect 4286 574 4288 576
rect 4296 574 4298 576
rect 4326 574 4328 576
rect 4356 574 4358 576
rect 4442 574 4444 576
rect 4472 574 4474 576
rect 4502 574 4504 576
rect 4512 574 4514 576
rect 4532 574 4534 576
rect 4542 574 4544 576
rect 4562 574 4564 576
rect 4572 574 4574 576
rect 4592 574 4594 576
rect 4602 574 4604 576
rect 4622 574 4624 576
rect 4632 574 4634 576
rect 4642 574 4644 576
rect 4664 574 4666 576
rect 4674 574 4676 576
rect 4694 574 4696 576
rect 4704 574 4706 576
rect 4724 574 4726 576
rect 4734 574 4736 576
rect 4756 574 4758 576
rect 4766 574 4768 576
rect 4776 574 4778 576
rect 4796 574 4798 576
rect 4806 574 4808 576
rect 4826 574 4828 576
rect 4836 574 4838 576
rect 4856 574 4858 576
rect 4866 574 4868 576
rect 4886 574 4888 576
rect 4896 574 4898 576
rect 4926 574 4928 576
rect 4956 574 4958 576
rect 5042 574 5044 576
rect 5072 574 5074 576
rect 5102 574 5104 576
rect 5112 574 5114 576
rect 5132 574 5134 576
rect 5142 574 5144 576
rect 5162 574 5164 576
rect 5172 574 5174 576
rect 5192 574 5194 576
rect 5202 574 5204 576
rect 5222 574 5224 576
rect 5232 574 5234 576
rect 5242 574 5244 576
rect 5264 574 5266 576
rect 5274 574 5276 576
rect 5294 574 5296 576
rect 5304 574 5306 576
rect 5324 574 5326 576
rect 5334 574 5336 576
rect 5356 574 5358 576
rect 5366 574 5368 576
rect 5376 574 5378 576
rect 5396 574 5398 576
rect 5406 574 5408 576
rect 5426 574 5428 576
rect 5436 574 5438 576
rect 5456 574 5458 576
rect 5466 574 5468 576
rect 5486 574 5488 576
rect 5496 574 5498 576
rect 5526 574 5528 576
rect 5556 574 5558 576
rect 5642 574 5644 576
rect 5672 574 5674 576
rect 5702 574 5704 576
rect 5712 574 5714 576
rect 5732 574 5734 576
rect 5742 574 5744 576
rect 5762 574 5764 576
rect 5772 574 5774 576
rect 5792 574 5794 576
rect 5802 574 5804 576
rect 5822 574 5824 576
rect 5832 574 5834 576
rect 5842 574 5844 576
rect 5864 574 5866 576
rect 5874 574 5876 576
rect 5894 574 5896 576
rect 5904 574 5906 576
rect 5924 574 5926 576
rect 5934 574 5936 576
rect 5956 574 5958 576
rect 5966 574 5968 576
rect 5976 574 5978 576
rect 5996 574 5998 576
rect 6006 574 6008 576
rect 6026 574 6028 576
rect 6036 574 6038 576
rect 6056 574 6058 576
rect 6066 574 6068 576
rect 6086 574 6088 576
rect 6096 574 6098 576
rect 6126 574 6128 576
rect 6156 574 6158 576
rect 6242 574 6244 576
rect 6272 574 6274 576
rect 6302 574 6304 576
rect 6312 574 6314 576
rect 6332 574 6334 576
rect 6342 574 6344 576
rect 6362 574 6364 576
rect 6372 574 6374 576
rect 6626 574 6628 576
rect 6636 574 6638 576
rect 6656 574 6658 576
rect 6666 574 6668 576
rect 6686 574 6688 576
rect 6696 574 6698 576
rect 6726 574 6728 576
rect 6756 574 6758 576
rect 1760 572 1762 574
rect 1766 572 1768 574
rect 1790 572 1792 574
rect 1796 572 1798 574
rect 1820 572 1822 574
rect 1826 572 1828 574
rect 1840 572 1842 574
rect 1866 572 1868 574
rect 1880 572 1882 574
rect 1886 572 1888 574
rect 1910 572 1912 574
rect 1916 572 1918 574
rect 1940 572 1942 574
rect 1946 572 1948 574
rect 1970 572 1972 574
rect 1976 572 1978 574
rect 3234 572 3236 574
rect 3240 572 3242 574
rect 3264 572 3266 574
rect 3270 572 3272 574
rect 3294 572 3296 574
rect 3300 572 3302 574
rect 3314 572 3316 574
rect 3330 572 3332 574
rect 3344 572 3346 574
rect 3360 572 3362 574
rect 3374 572 3376 574
rect 3624 572 3626 574
rect 3638 572 3640 574
rect 3654 572 3656 574
rect 3668 572 3670 574
rect 3684 572 3686 574
rect 3698 572 3700 574
rect 3704 572 3706 574
rect 3728 572 3730 574
rect 3734 572 3736 574
rect 3758 572 3760 574
rect 3764 572 3766 574
rect 3834 572 3836 574
rect 3840 572 3842 574
rect 3864 572 3866 574
rect 3870 572 3872 574
rect 3894 572 3896 574
rect 3900 572 3902 574
rect 3914 572 3916 574
rect 3930 572 3932 574
rect 3944 572 3946 574
rect 3960 572 3962 574
rect 3974 572 3976 574
rect 4224 572 4226 574
rect 4238 572 4240 574
rect 4254 572 4256 574
rect 4268 572 4270 574
rect 4284 572 4286 574
rect 4298 572 4300 574
rect 4304 572 4306 574
rect 4328 572 4330 574
rect 4334 572 4336 574
rect 4358 572 4360 574
rect 4364 572 4366 574
rect 4434 572 4436 574
rect 4440 572 4442 574
rect 4464 572 4466 574
rect 4470 572 4472 574
rect 4494 572 4496 574
rect 4500 572 4502 574
rect 4514 572 4516 574
rect 4530 572 4532 574
rect 4544 572 4546 574
rect 4560 572 4562 574
rect 4574 572 4576 574
rect 4590 572 4592 574
rect 4604 572 4606 574
rect 4620 572 4622 574
rect 4634 572 4636 574
rect 4640 572 4642 574
rect 4662 572 4664 574
rect 4676 572 4678 574
rect 4692 572 4694 574
rect 4706 572 4708 574
rect 4722 572 4724 574
rect 4736 572 4738 574
rect 4758 572 4760 574
rect 4764 572 4766 574
rect 4778 572 4780 574
rect 4794 572 4796 574
rect 4808 572 4810 574
rect 4824 572 4826 574
rect 4838 572 4840 574
rect 4854 572 4856 574
rect 4868 572 4870 574
rect 4884 572 4886 574
rect 4898 572 4900 574
rect 4904 572 4906 574
rect 4928 572 4930 574
rect 4934 572 4936 574
rect 4958 572 4960 574
rect 4964 572 4966 574
rect 5034 572 5036 574
rect 5040 572 5042 574
rect 5064 572 5066 574
rect 5070 572 5072 574
rect 5094 572 5096 574
rect 5100 572 5102 574
rect 5114 572 5116 574
rect 5130 572 5132 574
rect 5144 572 5146 574
rect 5160 572 5162 574
rect 5174 572 5176 574
rect 5190 572 5192 574
rect 5204 572 5206 574
rect 5220 572 5222 574
rect 5234 572 5236 574
rect 5240 572 5242 574
rect 5262 572 5264 574
rect 5276 572 5278 574
rect 5292 572 5294 574
rect 5306 572 5308 574
rect 5322 572 5324 574
rect 5336 572 5338 574
rect 5358 572 5360 574
rect 5364 572 5366 574
rect 5378 572 5380 574
rect 5394 572 5396 574
rect 5408 572 5410 574
rect 5424 572 5426 574
rect 5438 572 5440 574
rect 5454 572 5456 574
rect 5468 572 5470 574
rect 5484 572 5486 574
rect 5498 572 5500 574
rect 5504 572 5506 574
rect 5528 572 5530 574
rect 5534 572 5536 574
rect 5558 572 5560 574
rect 5564 572 5566 574
rect 5634 572 5636 574
rect 5640 572 5642 574
rect 5664 572 5666 574
rect 5670 572 5672 574
rect 5694 572 5696 574
rect 5700 572 5702 574
rect 5714 572 5716 574
rect 5730 572 5732 574
rect 5744 572 5746 574
rect 5760 572 5762 574
rect 5774 572 5776 574
rect 5790 572 5792 574
rect 5804 572 5806 574
rect 5820 572 5822 574
rect 5834 572 5836 574
rect 5840 572 5842 574
rect 5862 572 5864 574
rect 5876 572 5878 574
rect 5892 572 5894 574
rect 5906 572 5908 574
rect 5922 572 5924 574
rect 5936 572 5938 574
rect 5958 572 5960 574
rect 5964 572 5966 574
rect 5978 572 5980 574
rect 5994 572 5996 574
rect 6008 572 6010 574
rect 6024 572 6026 574
rect 6038 572 6040 574
rect 6054 572 6056 574
rect 6068 572 6070 574
rect 6084 572 6086 574
rect 6098 572 6100 574
rect 6104 572 6106 574
rect 6128 572 6130 574
rect 6134 572 6136 574
rect 6158 572 6160 574
rect 6164 572 6166 574
rect 6234 572 6236 574
rect 6240 572 6242 574
rect 6264 572 6266 574
rect 6270 572 6272 574
rect 6294 572 6296 574
rect 6300 572 6302 574
rect 6314 572 6316 574
rect 6330 572 6332 574
rect 6344 572 6346 574
rect 6360 572 6362 574
rect 6374 572 6376 574
rect 6624 572 6626 574
rect 6638 572 6640 574
rect 6654 572 6656 574
rect 6668 572 6670 574
rect 6684 572 6686 574
rect 6698 572 6700 574
rect 6704 572 6706 574
rect 6728 572 6730 574
rect 6734 572 6736 574
rect 6758 572 6760 574
rect 6764 572 6766 574
rect 1758 570 1760 572
rect 1788 570 1790 572
rect 1818 570 1820 572
rect 1828 570 1830 572
rect 1838 570 1840 572
rect 1888 570 1890 572
rect 1918 570 1920 572
rect 1948 570 1950 572
rect 1978 570 1980 572
rect 3232 570 3234 572
rect 3262 570 3264 572
rect 3292 570 3294 572
rect 3706 570 3708 572
rect 3736 570 3738 572
rect 3766 570 3768 572
rect 3832 570 3834 572
rect 3862 570 3864 572
rect 3892 570 3894 572
rect 4306 570 4308 572
rect 4336 570 4338 572
rect 4366 570 4368 572
rect 4432 570 4434 572
rect 4462 570 4464 572
rect 4492 570 4494 572
rect 4906 570 4908 572
rect 4936 570 4938 572
rect 4966 570 4968 572
rect 5032 570 5034 572
rect 5062 570 5064 572
rect 5092 570 5094 572
rect 5506 570 5508 572
rect 5536 570 5538 572
rect 5566 570 5568 572
rect 5632 570 5634 572
rect 5662 570 5664 572
rect 5692 570 5694 572
rect 6106 570 6108 572
rect 6136 570 6138 572
rect 6166 570 6168 572
rect 6232 570 6234 572
rect 6262 570 6264 572
rect 6292 570 6294 572
rect 6706 570 6708 572
rect 6736 570 6738 572
rect 6766 570 6768 572
rect 1758 564 1760 566
rect 1788 564 1790 566
rect 1858 564 1860 566
rect 1888 564 1890 566
rect 1918 564 1920 566
rect 1948 564 1950 566
rect 1978 564 1980 566
rect 3232 564 3234 566
rect 3262 564 3264 566
rect 3292 564 3294 566
rect 3322 564 3324 566
rect 3352 564 3354 566
rect 3382 564 3384 566
rect 3616 564 3618 566
rect 3646 564 3648 566
rect 3676 564 3678 566
rect 3706 564 3708 566
rect 3736 564 3738 566
rect 3766 564 3768 566
rect 3832 564 3834 566
rect 3862 564 3864 566
rect 3892 564 3894 566
rect 3922 564 3924 566
rect 3952 564 3954 566
rect 3982 564 3984 566
rect 4216 564 4218 566
rect 4246 564 4248 566
rect 4276 564 4278 566
rect 4306 564 4308 566
rect 4336 564 4338 566
rect 4366 564 4368 566
rect 4432 564 4434 566
rect 4462 564 4464 566
rect 4492 564 4494 566
rect 4522 564 4524 566
rect 4552 564 4554 566
rect 4582 564 4584 566
rect 4612 564 4614 566
rect 4684 564 4686 566
rect 4714 564 4716 566
rect 4786 564 4788 566
rect 4816 564 4818 566
rect 4846 564 4848 566
rect 4876 564 4878 566
rect 4906 564 4908 566
rect 4936 564 4938 566
rect 4966 564 4968 566
rect 5032 564 5034 566
rect 5062 564 5064 566
rect 5092 564 5094 566
rect 5122 564 5124 566
rect 5152 564 5154 566
rect 5182 564 5184 566
rect 5212 564 5214 566
rect 5284 564 5286 566
rect 5314 564 5316 566
rect 5386 564 5388 566
rect 5416 564 5418 566
rect 5446 564 5448 566
rect 5476 564 5478 566
rect 5506 564 5508 566
rect 5536 564 5538 566
rect 5566 564 5568 566
rect 5632 564 5634 566
rect 5662 564 5664 566
rect 5692 564 5694 566
rect 5722 564 5724 566
rect 5752 564 5754 566
rect 5782 564 5784 566
rect 5812 564 5814 566
rect 5884 564 5886 566
rect 5914 564 5916 566
rect 5986 564 5988 566
rect 6016 564 6018 566
rect 6046 564 6048 566
rect 6076 564 6078 566
rect 6106 564 6108 566
rect 6136 564 6138 566
rect 6166 564 6168 566
rect 6232 564 6234 566
rect 6262 564 6264 566
rect 6292 564 6294 566
rect 6322 564 6324 566
rect 6352 564 6354 566
rect 6382 564 6384 566
rect 6616 564 6618 566
rect 6646 564 6648 566
rect 6676 564 6678 566
rect 6706 564 6708 566
rect 6736 564 6738 566
rect 6766 564 6768 566
rect 1750 562 1752 564
rect 1756 562 1758 564
rect 1780 562 1782 564
rect 1786 562 1788 564
rect 1810 562 1812 564
rect 1856 562 1858 564
rect 1880 562 1882 564
rect 1886 562 1888 564
rect 1910 562 1912 564
rect 1916 562 1918 564
rect 1940 562 1942 564
rect 1946 562 1948 564
rect 1970 562 1972 564
rect 1976 562 1978 564
rect 3234 562 3236 564
rect 3240 562 3242 564
rect 3264 562 3266 564
rect 3270 562 3272 564
rect 3294 562 3296 564
rect 3300 562 3302 564
rect 3324 562 3326 564
rect 3330 562 3332 564
rect 3354 562 3356 564
rect 3360 562 3362 564
rect 3384 562 3386 564
rect 3614 562 3616 564
rect 3638 562 3640 564
rect 3644 562 3646 564
rect 3668 562 3670 564
rect 3674 562 3676 564
rect 3698 562 3700 564
rect 3704 562 3706 564
rect 3728 562 3730 564
rect 3734 562 3736 564
rect 3758 562 3760 564
rect 3764 562 3766 564
rect 3834 562 3836 564
rect 3840 562 3842 564
rect 3864 562 3866 564
rect 3870 562 3872 564
rect 3894 562 3896 564
rect 3900 562 3902 564
rect 3924 562 3926 564
rect 3930 562 3932 564
rect 3954 562 3956 564
rect 3960 562 3962 564
rect 3984 562 3986 564
rect 4214 562 4216 564
rect 4238 562 4240 564
rect 4244 562 4246 564
rect 4268 562 4270 564
rect 4274 562 4276 564
rect 4298 562 4300 564
rect 4304 562 4306 564
rect 4328 562 4330 564
rect 4334 562 4336 564
rect 4358 562 4360 564
rect 4364 562 4366 564
rect 4434 562 4436 564
rect 4440 562 4442 564
rect 4464 562 4466 564
rect 4470 562 4472 564
rect 4494 562 4496 564
rect 4500 562 4502 564
rect 4524 562 4526 564
rect 4530 562 4532 564
rect 4554 562 4556 564
rect 4560 562 4562 564
rect 4584 562 4586 564
rect 4590 562 4592 564
rect 4614 562 4616 564
rect 4620 562 4622 564
rect 4686 562 4688 564
rect 4692 562 4694 564
rect 4716 562 4718 564
rect 4722 562 4724 564
rect 4778 562 4780 564
rect 4784 562 4786 564
rect 4808 562 4810 564
rect 4814 562 4816 564
rect 4838 562 4840 564
rect 4844 562 4846 564
rect 4868 562 4870 564
rect 4874 562 4876 564
rect 4898 562 4900 564
rect 4904 562 4906 564
rect 4928 562 4930 564
rect 4934 562 4936 564
rect 4958 562 4960 564
rect 4964 562 4966 564
rect 5034 562 5036 564
rect 5040 562 5042 564
rect 5064 562 5066 564
rect 5070 562 5072 564
rect 5094 562 5096 564
rect 5100 562 5102 564
rect 5124 562 5126 564
rect 5130 562 5132 564
rect 5154 562 5156 564
rect 5160 562 5162 564
rect 5184 562 5186 564
rect 5190 562 5192 564
rect 5214 562 5216 564
rect 5220 562 5222 564
rect 5286 562 5288 564
rect 5292 562 5294 564
rect 5316 562 5318 564
rect 5322 562 5324 564
rect 5378 562 5380 564
rect 5384 562 5386 564
rect 5408 562 5410 564
rect 5414 562 5416 564
rect 5438 562 5440 564
rect 5444 562 5446 564
rect 5468 562 5470 564
rect 5474 562 5476 564
rect 5498 562 5500 564
rect 5504 562 5506 564
rect 5528 562 5530 564
rect 5534 562 5536 564
rect 5558 562 5560 564
rect 5564 562 5566 564
rect 5634 562 5636 564
rect 5640 562 5642 564
rect 5664 562 5666 564
rect 5670 562 5672 564
rect 5694 562 5696 564
rect 5700 562 5702 564
rect 5724 562 5726 564
rect 5730 562 5732 564
rect 5754 562 5756 564
rect 5760 562 5762 564
rect 5784 562 5786 564
rect 5790 562 5792 564
rect 5814 562 5816 564
rect 5820 562 5822 564
rect 5886 562 5888 564
rect 5892 562 5894 564
rect 5916 562 5918 564
rect 5922 562 5924 564
rect 5978 562 5980 564
rect 5984 562 5986 564
rect 6008 562 6010 564
rect 6014 562 6016 564
rect 6038 562 6040 564
rect 6044 562 6046 564
rect 6068 562 6070 564
rect 6074 562 6076 564
rect 6098 562 6100 564
rect 6104 562 6106 564
rect 6128 562 6130 564
rect 6134 562 6136 564
rect 6158 562 6160 564
rect 6164 562 6166 564
rect 6234 562 6236 564
rect 6240 562 6242 564
rect 6264 562 6266 564
rect 6270 562 6272 564
rect 6294 562 6296 564
rect 6300 562 6302 564
rect 6324 562 6326 564
rect 6330 562 6332 564
rect 6354 562 6356 564
rect 6360 562 6362 564
rect 6384 562 6386 564
rect 6614 562 6616 564
rect 6638 562 6640 564
rect 6644 562 6646 564
rect 6668 562 6670 564
rect 6674 562 6676 564
rect 6698 562 6700 564
rect 6704 562 6706 564
rect 6728 562 6730 564
rect 6734 562 6736 564
rect 6758 562 6760 564
rect 6764 562 6766 564
rect 1748 560 1750 562
rect 1778 560 1780 562
rect 1808 560 1810 562
rect 1878 560 1880 562
rect 1908 560 1910 562
rect 1938 560 1940 562
rect 1968 560 1970 562
rect 3242 560 3244 562
rect 3272 560 3274 562
rect 3302 560 3304 562
rect 3332 560 3334 562
rect 3362 560 3364 562
rect 3636 560 3638 562
rect 3666 560 3668 562
rect 3696 560 3698 562
rect 3726 560 3728 562
rect 3756 560 3758 562
rect 3842 560 3844 562
rect 3872 560 3874 562
rect 3902 560 3904 562
rect 3932 560 3934 562
rect 3962 560 3964 562
rect 4236 560 4238 562
rect 4266 560 4268 562
rect 4296 560 4298 562
rect 4326 560 4328 562
rect 4356 560 4358 562
rect 4442 560 4444 562
rect 4472 560 4474 562
rect 4502 560 4504 562
rect 4532 560 4534 562
rect 4562 560 4564 562
rect 4592 560 4594 562
rect 4622 560 4624 562
rect 4694 560 4696 562
rect 4724 560 4726 562
rect 4776 560 4778 562
rect 4806 560 4808 562
rect 4836 560 4838 562
rect 4866 560 4868 562
rect 4896 560 4898 562
rect 4926 560 4928 562
rect 4956 560 4958 562
rect 5042 560 5044 562
rect 5072 560 5074 562
rect 5102 560 5104 562
rect 5132 560 5134 562
rect 5162 560 5164 562
rect 5192 560 5194 562
rect 5222 560 5224 562
rect 5294 560 5296 562
rect 5324 560 5326 562
rect 5376 560 5378 562
rect 5406 560 5408 562
rect 5436 560 5438 562
rect 5466 560 5468 562
rect 5496 560 5498 562
rect 5526 560 5528 562
rect 5556 560 5558 562
rect 5642 560 5644 562
rect 5672 560 5674 562
rect 5702 560 5704 562
rect 5732 560 5734 562
rect 5762 560 5764 562
rect 5792 560 5794 562
rect 5822 560 5824 562
rect 5894 560 5896 562
rect 5924 560 5926 562
rect 5976 560 5978 562
rect 6006 560 6008 562
rect 6036 560 6038 562
rect 6066 560 6068 562
rect 6096 560 6098 562
rect 6126 560 6128 562
rect 6156 560 6158 562
rect 6242 560 6244 562
rect 6272 560 6274 562
rect 6302 560 6304 562
rect 6332 560 6334 562
rect 6362 560 6364 562
rect 6636 560 6638 562
rect 6666 560 6668 562
rect 6696 560 6698 562
rect 6726 560 6728 562
rect 6756 560 6758 562
rect 1748 554 1750 556
rect 1778 554 1780 556
rect 1838 554 1840 556
rect 1848 554 1850 556
rect 1878 554 1880 556
rect 1908 554 1910 556
rect 1938 554 1940 556
rect 1968 554 1970 556
rect 3242 554 3244 556
rect 3272 554 3274 556
rect 3302 554 3304 556
rect 3332 554 3334 556
rect 3362 554 3364 556
rect 3636 554 3638 556
rect 3666 554 3668 556
rect 3696 554 3698 556
rect 3726 554 3728 556
rect 3756 554 3758 556
rect 3842 554 3844 556
rect 3872 554 3874 556
rect 3902 554 3904 556
rect 3932 554 3934 556
rect 3962 554 3964 556
rect 4236 554 4238 556
rect 4266 554 4268 556
rect 4296 554 4298 556
rect 4326 554 4328 556
rect 4356 554 4358 556
rect 4442 554 4444 556
rect 4472 554 4474 556
rect 4502 554 4504 556
rect 4532 554 4534 556
rect 4562 554 4564 556
rect 4592 554 4594 556
rect 4622 554 4624 556
rect 4694 554 4696 556
rect 4724 554 4726 556
rect 4776 554 4778 556
rect 4806 554 4808 556
rect 4836 554 4838 556
rect 4866 554 4868 556
rect 4896 554 4898 556
rect 4926 554 4928 556
rect 4956 554 4958 556
rect 5042 554 5044 556
rect 5072 554 5074 556
rect 5102 554 5104 556
rect 5132 554 5134 556
rect 5162 554 5164 556
rect 5192 554 5194 556
rect 5222 554 5224 556
rect 5294 554 5296 556
rect 5324 554 5326 556
rect 5376 554 5378 556
rect 5406 554 5408 556
rect 5436 554 5438 556
rect 5466 554 5468 556
rect 5496 554 5498 556
rect 5526 554 5528 556
rect 5556 554 5558 556
rect 5642 554 5644 556
rect 5672 554 5674 556
rect 5702 554 5704 556
rect 5732 554 5734 556
rect 5762 554 5764 556
rect 5792 554 5794 556
rect 5822 554 5824 556
rect 5894 554 5896 556
rect 5924 554 5926 556
rect 5976 554 5978 556
rect 6006 554 6008 556
rect 6036 554 6038 556
rect 6066 554 6068 556
rect 6096 554 6098 556
rect 6126 554 6128 556
rect 6156 554 6158 556
rect 6242 554 6244 556
rect 6272 554 6274 556
rect 6302 554 6304 556
rect 6332 554 6334 556
rect 6362 554 6364 556
rect 6636 554 6638 556
rect 6666 554 6668 556
rect 6696 554 6698 556
rect 6726 554 6728 556
rect 6756 554 6758 556
rect 1740 552 1742 554
rect 1746 552 1748 554
rect 1770 552 1772 554
rect 1776 552 1778 554
rect 1800 552 1802 554
rect 1836 552 1838 554
rect 1850 552 1852 554
rect 1856 552 1858 554
rect 1880 552 1882 554
rect 1886 552 1888 554
rect 1910 552 1912 554
rect 1916 552 1918 554
rect 1940 552 1942 554
rect 1946 552 1948 554
rect 1970 552 1972 554
rect 1976 552 1978 554
rect 3234 552 3236 554
rect 3240 552 3242 554
rect 3264 552 3266 554
rect 3270 552 3272 554
rect 3294 552 3296 554
rect 3300 552 3302 554
rect 3324 552 3326 554
rect 3330 552 3332 554
rect 3354 552 3356 554
rect 3360 552 3362 554
rect 3384 552 3386 554
rect 3614 552 3616 554
rect 3638 552 3640 554
rect 3644 552 3646 554
rect 3668 552 3670 554
rect 3674 552 3676 554
rect 3698 552 3700 554
rect 3704 552 3706 554
rect 3728 552 3730 554
rect 3734 552 3736 554
rect 3758 552 3760 554
rect 3764 552 3766 554
rect 3834 552 3836 554
rect 3840 552 3842 554
rect 3864 552 3866 554
rect 3870 552 3872 554
rect 3894 552 3896 554
rect 3900 552 3902 554
rect 3924 552 3926 554
rect 3930 552 3932 554
rect 3954 552 3956 554
rect 3960 552 3962 554
rect 3984 552 3986 554
rect 4214 552 4216 554
rect 4238 552 4240 554
rect 4244 552 4246 554
rect 4268 552 4270 554
rect 4274 552 4276 554
rect 4298 552 4300 554
rect 4304 552 4306 554
rect 4328 552 4330 554
rect 4334 552 4336 554
rect 4358 552 4360 554
rect 4364 552 4366 554
rect 4434 552 4436 554
rect 4440 552 4442 554
rect 4464 552 4466 554
rect 4470 552 4472 554
rect 4494 552 4496 554
rect 4500 552 4502 554
rect 4524 552 4526 554
rect 4530 552 4532 554
rect 4554 552 4556 554
rect 4560 552 4562 554
rect 4584 552 4586 554
rect 4590 552 4592 554
rect 4614 552 4616 554
rect 4620 552 4622 554
rect 4686 552 4688 554
rect 4692 552 4694 554
rect 4716 552 4718 554
rect 4722 552 4724 554
rect 4778 552 4780 554
rect 4784 552 4786 554
rect 4808 552 4810 554
rect 4814 552 4816 554
rect 4838 552 4840 554
rect 4844 552 4846 554
rect 4868 552 4870 554
rect 4874 552 4876 554
rect 4898 552 4900 554
rect 4904 552 4906 554
rect 4928 552 4930 554
rect 4934 552 4936 554
rect 4958 552 4960 554
rect 4964 552 4966 554
rect 5034 552 5036 554
rect 5040 552 5042 554
rect 5064 552 5066 554
rect 5070 552 5072 554
rect 5094 552 5096 554
rect 5100 552 5102 554
rect 5124 552 5126 554
rect 5130 552 5132 554
rect 5154 552 5156 554
rect 5160 552 5162 554
rect 5184 552 5186 554
rect 5190 552 5192 554
rect 5214 552 5216 554
rect 5220 552 5222 554
rect 5286 552 5288 554
rect 5292 552 5294 554
rect 5316 552 5318 554
rect 5322 552 5324 554
rect 5378 552 5380 554
rect 5384 552 5386 554
rect 5408 552 5410 554
rect 5414 552 5416 554
rect 5438 552 5440 554
rect 5444 552 5446 554
rect 5468 552 5470 554
rect 5474 552 5476 554
rect 5498 552 5500 554
rect 5504 552 5506 554
rect 5528 552 5530 554
rect 5534 552 5536 554
rect 5558 552 5560 554
rect 5564 552 5566 554
rect 5634 552 5636 554
rect 5640 552 5642 554
rect 5664 552 5666 554
rect 5670 552 5672 554
rect 5694 552 5696 554
rect 5700 552 5702 554
rect 5724 552 5726 554
rect 5730 552 5732 554
rect 5754 552 5756 554
rect 5760 552 5762 554
rect 5784 552 5786 554
rect 5790 552 5792 554
rect 5814 552 5816 554
rect 5820 552 5822 554
rect 5886 552 5888 554
rect 5892 552 5894 554
rect 5916 552 5918 554
rect 5922 552 5924 554
rect 5978 552 5980 554
rect 5984 552 5986 554
rect 6008 552 6010 554
rect 6014 552 6016 554
rect 6038 552 6040 554
rect 6044 552 6046 554
rect 6068 552 6070 554
rect 6074 552 6076 554
rect 6098 552 6100 554
rect 6104 552 6106 554
rect 6128 552 6130 554
rect 6134 552 6136 554
rect 6158 552 6160 554
rect 6164 552 6166 554
rect 6234 552 6236 554
rect 6240 552 6242 554
rect 6264 552 6266 554
rect 6270 552 6272 554
rect 6294 552 6296 554
rect 6300 552 6302 554
rect 6324 552 6326 554
rect 6330 552 6332 554
rect 6354 552 6356 554
rect 6360 552 6362 554
rect 6384 552 6386 554
rect 6614 552 6616 554
rect 6638 552 6640 554
rect 6644 552 6646 554
rect 6668 552 6670 554
rect 6674 552 6676 554
rect 6698 552 6700 554
rect 6704 552 6706 554
rect 6728 552 6730 554
rect 6734 552 6736 554
rect 6758 552 6760 554
rect 6764 552 6766 554
rect 1738 550 1740 552
rect 1768 550 1770 552
rect 1798 550 1800 552
rect 1858 550 1860 552
rect 1888 550 1890 552
rect 1918 550 1920 552
rect 1948 550 1950 552
rect 1978 550 1980 552
rect 3232 550 3234 552
rect 3262 550 3264 552
rect 3292 550 3294 552
rect 3322 550 3324 552
rect 3352 550 3354 552
rect 3382 550 3384 552
rect 3616 550 3618 552
rect 3646 550 3648 552
rect 3676 550 3678 552
rect 3706 550 3708 552
rect 3736 550 3738 552
rect 3766 550 3768 552
rect 3832 550 3834 552
rect 3862 550 3864 552
rect 3892 550 3894 552
rect 3922 550 3924 552
rect 3952 550 3954 552
rect 3982 550 3984 552
rect 4216 550 4218 552
rect 4246 550 4248 552
rect 4276 550 4278 552
rect 4306 550 4308 552
rect 4336 550 4338 552
rect 4366 550 4368 552
rect 4432 550 4434 552
rect 4462 550 4464 552
rect 4492 550 4494 552
rect 4522 550 4524 552
rect 4552 550 4554 552
rect 4582 550 4584 552
rect 4612 550 4614 552
rect 4684 550 4686 552
rect 4714 550 4716 552
rect 4786 550 4788 552
rect 4816 550 4818 552
rect 4846 550 4848 552
rect 4876 550 4878 552
rect 4906 550 4908 552
rect 4936 550 4938 552
rect 4966 550 4968 552
rect 5032 550 5034 552
rect 5062 550 5064 552
rect 5092 550 5094 552
rect 5122 550 5124 552
rect 5152 550 5154 552
rect 5182 550 5184 552
rect 5212 550 5214 552
rect 5284 550 5286 552
rect 5314 550 5316 552
rect 5386 550 5388 552
rect 5416 550 5418 552
rect 5446 550 5448 552
rect 5476 550 5478 552
rect 5506 550 5508 552
rect 5536 550 5538 552
rect 5566 550 5568 552
rect 5632 550 5634 552
rect 5662 550 5664 552
rect 5692 550 5694 552
rect 5722 550 5724 552
rect 5752 550 5754 552
rect 5782 550 5784 552
rect 5812 550 5814 552
rect 5884 550 5886 552
rect 5914 550 5916 552
rect 5986 550 5988 552
rect 6016 550 6018 552
rect 6046 550 6048 552
rect 6076 550 6078 552
rect 6106 550 6108 552
rect 6136 550 6138 552
rect 6166 550 6168 552
rect 6232 550 6234 552
rect 6262 550 6264 552
rect 6292 550 6294 552
rect 6322 550 6324 552
rect 6352 550 6354 552
rect 6382 550 6384 552
rect 6616 550 6618 552
rect 6646 550 6648 552
rect 6676 550 6678 552
rect 6706 550 6708 552
rect 6736 550 6738 552
rect 6766 550 6768 552
rect 1738 544 1740 546
rect 1768 544 1770 546
rect 1828 544 1830 546
rect 1858 544 1860 546
rect 1888 544 1890 546
rect 1918 544 1920 546
rect 1948 544 1950 546
rect 1978 544 1980 546
rect 3232 544 3234 546
rect 3262 544 3264 546
rect 3292 544 3294 546
rect 3322 544 3324 546
rect 3352 544 3354 546
rect 3382 544 3384 546
rect 3616 544 3618 546
rect 3646 544 3648 546
rect 3676 544 3678 546
rect 3706 544 3708 546
rect 3736 544 3738 546
rect 3766 544 3768 546
rect 3832 544 3834 546
rect 3862 544 3864 546
rect 3892 544 3894 546
rect 3922 544 3924 546
rect 3952 544 3954 546
rect 3982 544 3984 546
rect 4216 544 4218 546
rect 4246 544 4248 546
rect 4276 544 4278 546
rect 4306 544 4308 546
rect 4336 544 4338 546
rect 4366 544 4368 546
rect 4432 544 4434 546
rect 4462 544 4464 546
rect 4492 544 4494 546
rect 4522 544 4524 546
rect 4552 544 4554 546
rect 4582 544 4584 546
rect 4612 544 4614 546
rect 4684 544 4686 546
rect 4714 544 4716 546
rect 4786 544 4788 546
rect 4816 544 4818 546
rect 4846 544 4848 546
rect 4876 544 4878 546
rect 4906 544 4908 546
rect 4936 544 4938 546
rect 4966 544 4968 546
rect 5032 544 5034 546
rect 5062 544 5064 546
rect 5092 544 5094 546
rect 5122 544 5124 546
rect 5152 544 5154 546
rect 5182 544 5184 546
rect 5212 544 5214 546
rect 5284 544 5286 546
rect 5314 544 5316 546
rect 5386 544 5388 546
rect 5416 544 5418 546
rect 5446 544 5448 546
rect 5476 544 5478 546
rect 5506 544 5508 546
rect 5536 544 5538 546
rect 5566 544 5568 546
rect 5632 544 5634 546
rect 5662 544 5664 546
rect 5692 544 5694 546
rect 5722 544 5724 546
rect 5752 544 5754 546
rect 5782 544 5784 546
rect 5812 544 5814 546
rect 5884 544 5886 546
rect 5914 544 5916 546
rect 5986 544 5988 546
rect 6016 544 6018 546
rect 6046 544 6048 546
rect 6076 544 6078 546
rect 6106 544 6108 546
rect 6136 544 6138 546
rect 6166 544 6168 546
rect 6232 544 6234 546
rect 6262 544 6264 546
rect 6292 544 6294 546
rect 6322 544 6324 546
rect 6352 544 6354 546
rect 6382 544 6384 546
rect 6616 544 6618 546
rect 6646 544 6648 546
rect 6676 544 6678 546
rect 6706 544 6708 546
rect 6736 544 6738 546
rect 6766 544 6768 546
rect 1730 542 1732 544
rect 1736 542 1738 544
rect 1760 542 1762 544
rect 1766 542 1768 544
rect 1790 542 1792 544
rect 1826 542 1828 544
rect 1850 542 1852 544
rect 1856 542 1858 544
rect 1880 542 1882 544
rect 1886 542 1888 544
rect 1910 542 1912 544
rect 1916 542 1918 544
rect 1940 542 1942 544
rect 1946 542 1948 544
rect 1970 542 1972 544
rect 1976 542 1978 544
rect 2580 543 2590 544
rect 3180 543 3190 544
rect 1728 540 1730 542
rect 1758 540 1760 542
rect 1788 540 1790 542
rect 1848 540 1850 542
rect 1878 540 1880 542
rect 1908 540 1910 542
rect 1938 540 1940 542
rect 1968 540 1970 542
rect 2580 541 2592 543
rect 3180 541 3192 543
rect 3234 542 3236 544
rect 3240 542 3242 544
rect 3264 542 3266 544
rect 3270 542 3272 544
rect 3294 542 3296 544
rect 3300 542 3302 544
rect 3324 542 3326 544
rect 3330 542 3332 544
rect 3354 542 3356 544
rect 3360 542 3362 544
rect 3384 542 3386 544
rect 3614 542 3616 544
rect 3638 542 3640 544
rect 3644 542 3646 544
rect 3668 542 3670 544
rect 3674 542 3676 544
rect 3698 542 3700 544
rect 3704 542 3706 544
rect 3728 542 3730 544
rect 3734 542 3736 544
rect 3758 542 3760 544
rect 3764 542 3766 544
rect 3834 542 3836 544
rect 3840 542 3842 544
rect 3864 542 3866 544
rect 3870 542 3872 544
rect 3894 542 3896 544
rect 3900 542 3902 544
rect 3924 542 3926 544
rect 3930 542 3932 544
rect 3954 542 3956 544
rect 3960 542 3962 544
rect 3984 542 3986 544
rect 4214 542 4216 544
rect 4238 542 4240 544
rect 4244 542 4246 544
rect 4268 542 4270 544
rect 4274 542 4276 544
rect 4298 542 4300 544
rect 4304 542 4306 544
rect 4328 542 4330 544
rect 4334 542 4336 544
rect 4358 542 4360 544
rect 4364 542 4366 544
rect 4434 542 4436 544
rect 4440 542 4442 544
rect 4464 542 4466 544
rect 4470 542 4472 544
rect 4494 542 4496 544
rect 4500 542 4502 544
rect 4524 542 4526 544
rect 4530 542 4532 544
rect 4554 542 4556 544
rect 4560 542 4562 544
rect 4584 542 4586 544
rect 4590 542 4592 544
rect 4614 542 4616 544
rect 4620 542 4622 544
rect 4686 542 4688 544
rect 4692 542 4694 544
rect 4716 542 4718 544
rect 4722 542 4724 544
rect 4778 542 4780 544
rect 4784 542 4786 544
rect 4808 542 4810 544
rect 4814 542 4816 544
rect 4838 542 4840 544
rect 4844 542 4846 544
rect 4868 542 4870 544
rect 4874 542 4876 544
rect 4898 542 4900 544
rect 4904 542 4906 544
rect 4928 542 4930 544
rect 4934 542 4936 544
rect 4958 542 4960 544
rect 4964 542 4966 544
rect 5034 542 5036 544
rect 5040 542 5042 544
rect 5064 542 5066 544
rect 5070 542 5072 544
rect 5094 542 5096 544
rect 5100 542 5102 544
rect 5124 542 5126 544
rect 5130 542 5132 544
rect 5154 542 5156 544
rect 5160 542 5162 544
rect 5184 542 5186 544
rect 5190 542 5192 544
rect 5214 542 5216 544
rect 5220 542 5222 544
rect 5286 542 5288 544
rect 5292 542 5294 544
rect 5316 542 5318 544
rect 5322 542 5324 544
rect 5378 542 5380 544
rect 5384 542 5386 544
rect 5408 542 5410 544
rect 5414 542 5416 544
rect 5438 542 5440 544
rect 5444 542 5446 544
rect 5468 542 5470 544
rect 5474 542 5476 544
rect 5498 542 5500 544
rect 5504 542 5506 544
rect 5528 542 5530 544
rect 5534 542 5536 544
rect 5558 542 5560 544
rect 5564 542 5566 544
rect 5634 542 5636 544
rect 5640 542 5642 544
rect 5664 542 5666 544
rect 5670 542 5672 544
rect 5694 542 5696 544
rect 5700 542 5702 544
rect 5724 542 5726 544
rect 5730 542 5732 544
rect 5754 542 5756 544
rect 5760 542 5762 544
rect 5784 542 5786 544
rect 5790 542 5792 544
rect 5814 542 5816 544
rect 5820 542 5822 544
rect 5886 542 5888 544
rect 5892 542 5894 544
rect 5916 542 5918 544
rect 5922 542 5924 544
rect 5978 542 5980 544
rect 5984 542 5986 544
rect 6008 542 6010 544
rect 6014 542 6016 544
rect 6038 542 6040 544
rect 6044 542 6046 544
rect 6068 542 6070 544
rect 6074 542 6076 544
rect 6098 542 6100 544
rect 6104 542 6106 544
rect 6128 542 6130 544
rect 6134 542 6136 544
rect 6158 542 6160 544
rect 6164 542 6166 544
rect 6234 542 6236 544
rect 6240 542 6242 544
rect 6264 542 6266 544
rect 6270 542 6272 544
rect 6294 542 6296 544
rect 6300 542 6302 544
rect 6324 542 6326 544
rect 6330 542 6332 544
rect 6354 542 6356 544
rect 6360 542 6362 544
rect 6384 542 6386 544
rect 6614 542 6616 544
rect 6638 542 6640 544
rect 6644 542 6646 544
rect 6668 542 6670 544
rect 6674 542 6676 544
rect 6698 542 6700 544
rect 6704 542 6706 544
rect 6728 542 6730 544
rect 6734 542 6736 544
rect 6758 542 6760 544
rect 6764 542 6766 544
rect 2588 539 2590 541
rect 3188 539 3190 541
rect 3242 540 3244 542
rect 3272 540 3274 542
rect 3302 540 3304 542
rect 3332 540 3334 542
rect 3362 540 3364 542
rect 3636 540 3638 542
rect 3666 540 3668 542
rect 3696 540 3698 542
rect 3726 540 3728 542
rect 3756 540 3758 542
rect 3842 540 3844 542
rect 3872 540 3874 542
rect 3902 540 3904 542
rect 3932 540 3934 542
rect 3962 540 3964 542
rect 4236 540 4238 542
rect 4266 540 4268 542
rect 4296 540 4298 542
rect 4326 540 4328 542
rect 4356 540 4358 542
rect 4442 540 4444 542
rect 4472 540 4474 542
rect 4502 540 4504 542
rect 4532 540 4534 542
rect 4562 540 4564 542
rect 4592 540 4594 542
rect 4622 540 4624 542
rect 4694 540 4696 542
rect 4724 540 4726 542
rect 4776 540 4778 542
rect 4806 540 4808 542
rect 4836 540 4838 542
rect 4866 540 4868 542
rect 4896 540 4898 542
rect 4926 540 4928 542
rect 4956 540 4958 542
rect 5042 540 5044 542
rect 5072 540 5074 542
rect 5102 540 5104 542
rect 5132 540 5134 542
rect 5162 540 5164 542
rect 5192 540 5194 542
rect 5222 540 5224 542
rect 5294 540 5296 542
rect 5324 540 5326 542
rect 5376 540 5378 542
rect 5406 540 5408 542
rect 5436 540 5438 542
rect 5466 540 5468 542
rect 5496 540 5498 542
rect 5526 540 5528 542
rect 5556 540 5558 542
rect 5642 540 5644 542
rect 5672 540 5674 542
rect 5702 540 5704 542
rect 5732 540 5734 542
rect 5762 540 5764 542
rect 5792 540 5794 542
rect 5822 540 5824 542
rect 5894 540 5896 542
rect 5924 540 5926 542
rect 5976 540 5978 542
rect 6006 540 6008 542
rect 6036 540 6038 542
rect 6066 540 6068 542
rect 6096 540 6098 542
rect 6126 540 6128 542
rect 6156 540 6158 542
rect 6242 540 6244 542
rect 6272 540 6274 542
rect 6302 540 6304 542
rect 6332 540 6334 542
rect 6362 540 6364 542
rect 6636 540 6638 542
rect 6666 540 6668 542
rect 6696 540 6698 542
rect 6726 540 6728 542
rect 6756 540 6758 542
rect 2588 536 2590 538
rect 3188 536 3190 538
rect 1728 534 1730 536
rect 1758 534 1760 536
rect 1808 534 1810 536
rect 1818 534 1820 536
rect 1848 534 1850 536
rect 1878 534 1880 536
rect 1908 534 1910 536
rect 1938 534 1940 536
rect 1968 534 1970 536
rect 1720 532 1722 534
rect 1726 532 1728 534
rect 1750 532 1752 534
rect 1756 532 1758 534
rect 1780 532 1782 534
rect 1718 530 1720 532
rect 1748 530 1750 532
rect 1778 530 1780 532
rect 1806 531 1808 534
rect 1820 531 1822 534
rect 1826 532 1828 534
rect 1850 532 1852 534
rect 1856 532 1858 534
rect 1880 532 1882 534
rect 1886 532 1888 534
rect 1910 532 1912 534
rect 1916 532 1918 534
rect 1940 532 1942 534
rect 1946 532 1948 534
rect 1970 532 1972 534
rect 1976 532 1978 534
rect 2158 533 2160 535
rect 2164 533 2166 535
rect 2392 533 2394 535
rect 2482 533 2484 535
rect 2488 533 2490 535
rect 2578 534 2580 535
rect 2586 534 2588 536
rect 2578 533 2590 534
rect 2758 533 2760 535
rect 2764 533 2766 535
rect 2992 533 2994 535
rect 3082 533 3084 535
rect 3088 533 3090 535
rect 3178 534 3180 535
rect 3186 534 3188 536
rect 3242 534 3244 536
rect 3272 534 3274 536
rect 3302 534 3304 536
rect 3332 534 3334 536
rect 3362 534 3364 536
rect 3636 534 3638 536
rect 3666 534 3668 536
rect 3696 534 3698 536
rect 3726 534 3728 536
rect 3756 534 3758 536
rect 3842 534 3844 536
rect 3872 534 3874 536
rect 3902 534 3904 536
rect 3932 534 3934 536
rect 3962 534 3964 536
rect 4236 534 4238 536
rect 4266 534 4268 536
rect 4296 534 4298 536
rect 4326 534 4328 536
rect 4356 534 4358 536
rect 4442 534 4444 536
rect 4472 534 4474 536
rect 4502 534 4504 536
rect 4532 534 4534 536
rect 4562 534 4564 536
rect 4592 534 4594 536
rect 4622 534 4624 536
rect 4694 534 4696 536
rect 4724 534 4726 536
rect 4776 534 4778 536
rect 4806 534 4808 536
rect 4836 534 4838 536
rect 4866 534 4868 536
rect 4896 534 4898 536
rect 4926 534 4928 536
rect 4956 534 4958 536
rect 5042 534 5044 536
rect 5072 534 5074 536
rect 5102 534 5104 536
rect 5132 534 5134 536
rect 5162 534 5164 536
rect 5192 534 5194 536
rect 5222 534 5224 536
rect 5294 534 5296 536
rect 5324 534 5326 536
rect 5376 534 5378 536
rect 5406 534 5408 536
rect 5436 534 5438 536
rect 5466 534 5468 536
rect 5496 534 5498 536
rect 5526 534 5528 536
rect 5556 534 5558 536
rect 5642 534 5644 536
rect 5672 534 5674 536
rect 5702 534 5704 536
rect 5732 534 5734 536
rect 5762 534 5764 536
rect 5792 534 5794 536
rect 5822 534 5824 536
rect 5894 534 5896 536
rect 5924 534 5926 536
rect 5976 534 5978 536
rect 6006 534 6008 536
rect 6036 534 6038 536
rect 6066 534 6068 536
rect 6096 534 6098 536
rect 6126 534 6128 536
rect 6156 534 6158 536
rect 6242 534 6244 536
rect 6272 534 6274 536
rect 6302 534 6304 536
rect 6332 534 6334 536
rect 6362 534 6364 536
rect 6636 534 6638 536
rect 6666 534 6668 536
rect 6696 534 6698 536
rect 6726 534 6728 536
rect 6756 534 6758 536
rect 3178 533 3190 534
rect 1808 529 1810 531
rect 1818 529 1820 531
rect 1828 530 1830 532
rect 1858 530 1860 532
rect 1888 530 1890 532
rect 1918 530 1920 532
rect 1948 530 1950 532
rect 1978 530 1980 532
rect 2580 531 2592 533
rect 3180 531 3192 533
rect 3234 532 3236 534
rect 3240 532 3242 534
rect 3264 532 3266 534
rect 3270 532 3272 534
rect 3294 532 3296 534
rect 3300 532 3302 534
rect 3324 532 3326 534
rect 3330 532 3332 534
rect 3354 532 3356 534
rect 3360 532 3362 534
rect 3384 532 3386 534
rect 3614 532 3616 534
rect 3638 532 3640 534
rect 3644 532 3646 534
rect 3668 532 3670 534
rect 3674 532 3676 534
rect 3698 532 3700 534
rect 3704 532 3706 534
rect 3728 532 3730 534
rect 3734 532 3736 534
rect 3758 532 3760 534
rect 3764 532 3766 534
rect 3834 532 3836 534
rect 3840 532 3842 534
rect 3864 532 3866 534
rect 3870 532 3872 534
rect 3894 532 3896 534
rect 3900 532 3902 534
rect 3924 532 3926 534
rect 3930 532 3932 534
rect 3954 532 3956 534
rect 3960 532 3962 534
rect 3984 532 3986 534
rect 4214 532 4216 534
rect 4238 532 4240 534
rect 4244 532 4246 534
rect 4268 532 4270 534
rect 4274 532 4276 534
rect 4298 532 4300 534
rect 4304 532 4306 534
rect 4328 532 4330 534
rect 4334 532 4336 534
rect 4358 532 4360 534
rect 4364 532 4366 534
rect 4434 532 4436 534
rect 4440 532 4442 534
rect 4464 532 4466 534
rect 4470 532 4472 534
rect 4494 532 4496 534
rect 4500 532 4502 534
rect 4524 532 4526 534
rect 4530 532 4532 534
rect 4554 532 4556 534
rect 4560 532 4562 534
rect 4584 532 4586 534
rect 4590 532 4592 534
rect 4614 532 4616 534
rect 4620 532 4622 534
rect 4686 532 4688 534
rect 4692 532 4694 534
rect 4716 532 4718 534
rect 4722 532 4724 534
rect 4778 532 4780 534
rect 4784 532 4786 534
rect 4808 532 4810 534
rect 4814 532 4816 534
rect 4838 532 4840 534
rect 4844 532 4846 534
rect 4868 532 4870 534
rect 4874 532 4876 534
rect 4898 532 4900 534
rect 4904 532 4906 534
rect 4928 532 4930 534
rect 4934 532 4936 534
rect 4958 532 4960 534
rect 4964 532 4966 534
rect 5034 532 5036 534
rect 5040 532 5042 534
rect 5064 532 5066 534
rect 5070 532 5072 534
rect 5094 532 5096 534
rect 5100 532 5102 534
rect 5124 532 5126 534
rect 5130 532 5132 534
rect 5154 532 5156 534
rect 5160 532 5162 534
rect 5184 532 5186 534
rect 5190 532 5192 534
rect 5214 532 5216 534
rect 5220 532 5222 534
rect 5286 532 5288 534
rect 5292 532 5294 534
rect 5316 532 5318 534
rect 5322 532 5324 534
rect 5378 532 5380 534
rect 5384 532 5386 534
rect 5408 532 5410 534
rect 5414 532 5416 534
rect 5438 532 5440 534
rect 5444 532 5446 534
rect 5468 532 5470 534
rect 5474 532 5476 534
rect 5498 532 5500 534
rect 5504 532 5506 534
rect 5528 532 5530 534
rect 5534 532 5536 534
rect 5558 532 5560 534
rect 5564 532 5566 534
rect 5634 532 5636 534
rect 5640 532 5642 534
rect 5664 532 5666 534
rect 5670 532 5672 534
rect 5694 532 5696 534
rect 5700 532 5702 534
rect 5724 532 5726 534
rect 5730 532 5732 534
rect 5754 532 5756 534
rect 5760 532 5762 534
rect 5784 532 5786 534
rect 5790 532 5792 534
rect 5814 532 5816 534
rect 5820 532 5822 534
rect 5886 532 5888 534
rect 5892 532 5894 534
rect 5916 532 5918 534
rect 5922 532 5924 534
rect 5978 532 5980 534
rect 5984 532 5986 534
rect 6008 532 6010 534
rect 6014 532 6016 534
rect 6038 532 6040 534
rect 6044 532 6046 534
rect 6068 532 6070 534
rect 6074 532 6076 534
rect 6098 532 6100 534
rect 6104 532 6106 534
rect 6128 532 6130 534
rect 6134 532 6136 534
rect 6158 532 6160 534
rect 6164 532 6166 534
rect 6234 532 6236 534
rect 6240 532 6242 534
rect 6264 532 6266 534
rect 6270 532 6272 534
rect 6294 532 6296 534
rect 6300 532 6302 534
rect 6324 532 6326 534
rect 6330 532 6332 534
rect 6354 532 6356 534
rect 6360 532 6362 534
rect 6384 532 6386 534
rect 6614 532 6616 534
rect 6638 532 6640 534
rect 6644 532 6646 534
rect 6668 532 6670 534
rect 6674 532 6676 534
rect 6698 532 6700 534
rect 6704 532 6706 534
rect 6728 532 6730 534
rect 6734 532 6736 534
rect 6758 532 6760 534
rect 6764 532 6766 534
rect 6958 533 6960 535
rect 6964 533 6966 535
rect 7192 533 7194 535
rect 2588 529 2590 531
rect 3188 529 3190 531
rect 3232 530 3234 532
rect 3262 530 3264 532
rect 3292 530 3294 532
rect 3322 530 3324 532
rect 3352 530 3354 532
rect 3382 530 3384 532
rect 3616 530 3618 532
rect 3646 530 3648 532
rect 3676 530 3678 532
rect 3706 530 3708 532
rect 3736 530 3738 532
rect 3766 530 3768 532
rect 3832 530 3834 532
rect 3862 530 3864 532
rect 3892 530 3894 532
rect 3922 530 3924 532
rect 3952 530 3954 532
rect 3982 530 3984 532
rect 4216 530 4218 532
rect 4246 530 4248 532
rect 4276 530 4278 532
rect 4306 530 4308 532
rect 4336 530 4338 532
rect 4366 530 4368 532
rect 4432 530 4434 532
rect 4462 530 4464 532
rect 4492 530 4494 532
rect 4522 530 4524 532
rect 4552 530 4554 532
rect 4582 530 4584 532
rect 4612 530 4614 532
rect 4684 530 4686 532
rect 4714 530 4716 532
rect 4786 530 4788 532
rect 4816 530 4818 532
rect 4846 530 4848 532
rect 4876 530 4878 532
rect 4906 530 4908 532
rect 4936 530 4938 532
rect 4966 530 4968 532
rect 5032 530 5034 532
rect 5062 530 5064 532
rect 5092 530 5094 532
rect 5122 530 5124 532
rect 5152 530 5154 532
rect 5182 530 5184 532
rect 5212 530 5214 532
rect 5284 530 5286 532
rect 5314 530 5316 532
rect 5386 530 5388 532
rect 5416 530 5418 532
rect 5446 530 5448 532
rect 5476 530 5478 532
rect 5506 530 5508 532
rect 5536 530 5538 532
rect 5566 530 5568 532
rect 5632 530 5634 532
rect 5662 530 5664 532
rect 5692 530 5694 532
rect 5722 530 5724 532
rect 5752 530 5754 532
rect 5782 530 5784 532
rect 5812 530 5814 532
rect 5884 530 5886 532
rect 5914 530 5916 532
rect 5986 530 5988 532
rect 6016 530 6018 532
rect 6046 530 6048 532
rect 6076 530 6078 532
rect 6106 530 6108 532
rect 6136 530 6138 532
rect 6166 530 6168 532
rect 6232 530 6234 532
rect 6262 530 6264 532
rect 6292 530 6294 532
rect 6322 530 6324 532
rect 6352 530 6354 532
rect 6382 530 6384 532
rect 6616 530 6618 532
rect 6646 530 6648 532
rect 6676 530 6678 532
rect 6706 530 6708 532
rect 6736 530 6738 532
rect 6766 530 6768 532
rect 2588 526 2590 528
rect 3188 526 3190 528
rect 1718 524 1720 526
rect 1748 524 1750 526
rect 1710 522 1712 524
rect 1716 522 1718 524
rect 1740 522 1742 524
rect 1746 522 1748 524
rect 1770 522 1772 524
rect 1808 523 1810 525
rect 1818 523 1820 525
rect 1828 524 1830 526
rect 1858 524 1860 526
rect 1888 524 1890 526
rect 1918 524 1920 526
rect 1948 524 1950 526
rect 1978 524 1980 526
rect 2586 524 2588 526
rect 3186 524 3188 526
rect 1708 520 1710 522
rect 1738 520 1740 522
rect 1768 520 1770 522
rect 1806 521 1808 523
rect 1820 521 1822 523
rect 1826 522 1828 524
rect 1850 522 1852 524
rect 1856 522 1858 524
rect 1880 522 1882 524
rect 1886 522 1888 524
rect 1910 522 1912 524
rect 1916 522 1918 524
rect 1940 522 1942 524
rect 1946 522 1948 524
rect 1970 522 1972 524
rect 1976 522 1978 524
rect 1848 520 1850 522
rect 1878 520 1880 522
rect 1908 520 1910 522
rect 1938 520 1940 522
rect 1968 520 1970 522
rect 2580 521 2582 523
rect 3180 521 3182 523
rect 2216 518 2218 520
rect 2482 519 2484 521
rect 2488 519 2490 521
rect 2578 519 2580 521
rect 2218 516 2220 518
rect 2480 517 2482 519
rect 2490 517 2492 519
rect 2816 518 2818 520
rect 3082 519 3084 521
rect 3088 519 3090 521
rect 3178 519 3180 521
rect 2818 516 2820 518
rect 3080 517 3082 519
rect 3090 517 3092 519
rect 7016 518 7018 520
rect 7018 516 7020 518
rect 1708 514 1710 516
rect 1738 514 1740 516
rect 1798 514 1800 516
rect 1848 514 1850 516
rect 1878 514 1880 516
rect 1908 514 1910 516
rect 1938 514 1940 516
rect 1968 514 1970 516
rect 2208 514 2220 516
rect 2808 514 2820 516
rect 4986 514 4996 516
rect 5586 514 5596 516
rect 7008 514 7020 516
rect 1700 512 1702 514
rect 1706 512 1708 514
rect 1730 512 1732 514
rect 1736 512 1738 514
rect 1760 512 1762 514
rect 1796 512 1798 514
rect 1820 512 1822 514
rect 1826 512 1828 514
rect 1850 512 1852 514
rect 1856 512 1858 514
rect 1880 512 1882 514
rect 1886 512 1888 514
rect 1910 512 1912 514
rect 1916 512 1918 514
rect 1940 512 1942 514
rect 1946 512 1948 514
rect 1970 512 1972 514
rect 1976 512 1978 514
rect 2216 512 2218 514
rect 2816 512 2818 514
rect 4984 512 4996 514
rect 5584 512 5596 514
rect 7016 512 7018 514
rect 1698 510 1700 512
rect 1728 510 1730 512
rect 1758 510 1760 512
rect 1818 510 1820 512
rect 1828 510 1830 512
rect 1858 510 1860 512
rect 1888 510 1890 512
rect 1918 510 1920 512
rect 1948 510 1950 512
rect 1978 510 1980 512
rect 2216 508 2218 510
rect 2816 508 2818 510
rect 4986 508 4988 512
rect 5586 508 5588 512
rect 6186 508 6188 510
rect 7016 508 7018 510
rect 2214 506 2216 508
rect 2814 506 2816 508
rect 4988 506 4990 508
rect 5588 506 5590 508
rect 6188 506 6190 508
rect 7014 506 7016 508
rect 1690 502 1692 504
rect 1706 502 1708 504
rect 1720 502 1722 504
rect 1736 502 1738 504
rect 1750 502 1752 504
rect 1796 502 1798 504
rect 1810 502 1812 504
rect 1836 502 1838 504
rect 1850 502 1852 504
rect 1866 502 1868 504
rect 1880 502 1882 504
rect 1896 502 1898 504
rect 1910 502 1912 504
rect 1926 502 1928 504
rect 1940 502 1942 504
rect 1956 502 1958 504
rect 1970 502 1972 504
rect 1986 502 1988 504
rect 2590 502 2592 504
rect 3190 502 3192 504
rect 1688 500 1690 502
rect 1708 500 1710 502
rect 1718 500 1720 502
rect 1738 500 1740 502
rect 1748 500 1750 502
rect 1798 500 1800 502
rect 1808 500 1810 502
rect 1838 500 1840 502
rect 1848 500 1850 502
rect 1868 500 1870 502
rect 1878 500 1880 502
rect 1898 500 1900 502
rect 1908 500 1910 502
rect 1928 500 1930 502
rect 1938 500 1940 502
rect 1958 500 1960 502
rect 1968 500 1970 502
rect 1988 500 1990 502
rect 2588 500 2590 502
rect 3188 500 3190 502
rect 1688 494 1690 496
rect 1698 494 1700 496
rect 1708 494 1710 496
rect 1718 494 1720 496
rect 1728 494 1730 496
rect 1738 494 1740 496
rect 1748 494 1750 496
rect 1788 494 1790 496
rect 1798 494 1800 496
rect 1808 494 1810 496
rect 1818 494 1820 496
rect 1828 494 1830 496
rect 1838 494 1840 496
rect 1848 494 1850 496
rect 1858 494 1860 496
rect 1868 494 1870 496
rect 1888 494 1890 496
rect 1690 492 1692 494
rect 1696 492 1698 494
rect 1710 492 1712 494
rect 1716 492 1718 494
rect 1730 492 1732 494
rect 1736 492 1738 494
rect 1750 492 1752 494
rect 1786 492 1788 494
rect 1800 492 1802 494
rect 1806 492 1808 494
rect 1820 492 1822 494
rect 1826 492 1828 494
rect 1840 492 1842 494
rect 1846 492 1848 494
rect 1860 492 1862 494
rect 1866 492 1868 494
rect 1890 492 1892 494
rect 1778 484 1780 486
rect 1750 482 1752 484
rect 1776 482 1778 484
rect 1890 482 1892 484
rect 1748 480 1750 482
rect 1888 480 1890 482
rect 1768 474 1770 476
rect 1740 472 1742 474
rect 1766 472 1768 474
rect 1880 472 1882 474
rect 1738 470 1740 472
rect 1878 470 1880 472
rect 2106 468 2108 470
rect 2126 468 2128 470
rect 2136 468 2138 470
rect 2156 468 2158 470
rect 2166 468 2168 470
rect 2186 468 2188 470
rect 2196 468 2198 470
rect 2216 468 2218 470
rect 2226 468 2228 470
rect 2234 468 2236 476
rect 2382 468 2384 470
rect 2392 468 2394 470
rect 2412 468 2414 470
rect 2422 468 2424 470
rect 2442 468 2444 470
rect 2452 468 2454 470
rect 2472 468 2474 470
rect 2482 468 2484 470
rect 2706 468 2708 470
rect 2726 468 2728 470
rect 2736 468 2738 470
rect 2756 468 2758 470
rect 2766 468 2768 470
rect 2786 468 2788 470
rect 2796 468 2798 470
rect 2816 468 2818 470
rect 2826 468 2828 470
rect 2834 468 2836 476
rect 2982 468 2984 470
rect 2992 468 2994 470
rect 3012 468 3014 470
rect 3022 468 3024 470
rect 3042 468 3044 470
rect 3052 468 3054 470
rect 3072 468 3074 470
rect 3082 468 3084 470
rect 6906 468 6908 470
rect 6926 468 6928 470
rect 6936 468 6938 470
rect 6956 468 6958 470
rect 6966 468 6968 470
rect 6986 468 6988 470
rect 6996 468 6998 470
rect 7016 468 7018 470
rect 7026 468 7028 470
rect 7034 468 7036 476
rect 7182 468 7184 470
rect 7192 468 7194 470
rect 2052 466 2054 468
rect 2108 466 2110 468
rect 2124 466 2126 468
rect 2138 466 2140 468
rect 2154 466 2156 468
rect 2168 466 2170 468
rect 2184 466 2186 468
rect 2198 466 2200 468
rect 2214 466 2216 468
rect 2228 466 2230 468
rect 2232 466 2236 468
rect 2380 466 2382 468
rect 2394 466 2396 468
rect 2410 466 2412 468
rect 2424 466 2426 468
rect 2440 466 2442 468
rect 2454 466 2456 468
rect 2470 466 2472 468
rect 2484 466 2486 468
rect 2652 466 2654 468
rect 2708 466 2710 468
rect 2724 466 2726 468
rect 2738 466 2740 468
rect 2754 466 2756 468
rect 2768 466 2770 468
rect 2784 466 2786 468
rect 2798 466 2800 468
rect 2814 466 2816 468
rect 2828 466 2830 468
rect 2832 466 2836 468
rect 2980 466 2982 468
rect 2994 466 2996 468
rect 3010 466 3012 468
rect 3024 466 3026 468
rect 3040 466 3042 468
rect 3054 466 3056 468
rect 3070 466 3072 468
rect 3084 466 3086 468
rect 3718 466 3720 468
rect 4304 466 4306 468
rect 5656 466 5658 468
rect 5676 466 5678 468
rect 6122 466 6124 468
rect 6142 466 6144 468
rect 6852 466 6854 468
rect 6908 466 6910 468
rect 6924 466 6926 468
rect 6938 466 6940 468
rect 6954 466 6956 468
rect 6968 466 6970 468
rect 6984 466 6986 468
rect 6998 466 7000 468
rect 7014 466 7016 468
rect 7028 466 7030 468
rect 7032 466 7036 468
rect 7180 466 7182 468
rect 7194 466 7196 468
rect 1758 464 1760 466
rect 2050 464 2052 466
rect 2234 464 2236 466
rect 2650 464 2652 466
rect 2834 464 2836 466
rect 3716 464 3718 466
rect 4302 464 4304 466
rect 5654 464 5656 466
rect 5678 464 5680 466
rect 6120 464 6122 466
rect 6144 464 6146 466
rect 6850 464 6852 466
rect 7034 464 7036 466
rect 1730 462 1732 464
rect 1756 462 1758 464
rect 1870 462 1872 464
rect 1728 460 1730 462
rect 1868 460 1870 462
rect 4440 460 4442 462
rect 4450 460 4452 462
rect 4460 460 4462 462
rect 4480 460 4482 462
rect 4490 460 4492 462
rect 4510 460 4512 462
rect 4520 460 4522 462
rect 4540 460 4542 462
rect 4550 460 4552 462
rect 4570 460 4572 462
rect 4580 460 4582 462
rect 4600 460 4602 462
rect 4610 460 4612 462
rect 4630 460 4632 462
rect 4640 460 4642 462
rect 4660 460 4662 462
rect 4670 460 4672 462
rect 4690 460 4692 462
rect 4700 460 4702 462
rect 4720 460 4722 462
rect 4730 460 4732 462
rect 4750 460 4752 462
rect 4760 460 4762 462
rect 4780 460 4782 462
rect 4790 460 4792 462
rect 4810 460 4812 462
rect 4820 460 4822 462
rect 4840 460 4842 462
rect 4850 460 4852 462
rect 4870 460 4872 462
rect 4880 460 4882 462
rect 4900 460 4902 462
rect 4910 460 4912 462
rect 4930 460 4932 462
rect 4940 460 4942 462
rect 4960 460 4962 462
rect 5040 460 5042 462
rect 5050 460 5052 462
rect 5060 460 5062 462
rect 5080 460 5082 462
rect 5090 460 5092 462
rect 5110 460 5112 462
rect 5120 460 5122 462
rect 5140 460 5142 462
rect 5150 460 5152 462
rect 5170 460 5172 462
rect 5180 460 5182 462
rect 5200 460 5202 462
rect 5210 460 5212 462
rect 5230 460 5232 462
rect 5240 460 5242 462
rect 5260 460 5262 462
rect 5270 460 5272 462
rect 5290 460 5292 462
rect 5300 460 5302 462
rect 5320 460 5322 462
rect 5330 460 5332 462
rect 5350 460 5352 462
rect 5360 460 5362 462
rect 5380 460 5382 462
rect 5390 460 5392 462
rect 5410 460 5412 462
rect 5420 460 5422 462
rect 5440 460 5442 462
rect 5450 460 5452 462
rect 5470 460 5472 462
rect 5480 460 5482 462
rect 5500 460 5502 462
rect 5510 460 5512 462
rect 5530 460 5532 462
rect 5540 460 5542 462
rect 5560 460 5562 462
rect 6238 461 6240 463
rect 6248 461 6250 463
rect 6258 461 6260 463
rect 6278 461 6280 463
rect 6288 461 6290 463
rect 6308 461 6310 463
rect 6318 461 6320 463
rect 6338 461 6340 463
rect 6348 461 6350 463
rect 6368 461 6370 463
rect 6378 461 6380 463
rect 6398 461 6400 463
rect 6408 461 6410 463
rect 6428 461 6430 463
rect 6438 461 6440 463
rect 6458 461 6460 463
rect 6468 461 6470 463
rect 6488 461 6490 463
rect 6498 461 6500 463
rect 6518 461 6520 463
rect 6528 461 6530 463
rect 6548 461 6550 463
rect 6558 461 6560 463
rect 6578 461 6580 463
rect 6588 461 6590 463
rect 6608 461 6610 463
rect 6618 461 6620 463
rect 6638 461 6640 463
rect 6648 461 6650 463
rect 6668 461 6670 463
rect 6678 461 6680 463
rect 6698 461 6700 463
rect 6708 461 6710 463
rect 6728 461 6730 463
rect 6738 461 6740 463
rect 6758 461 6760 463
rect 4442 458 4444 460
rect 4448 458 4450 460
rect 4462 458 4464 460
rect 4478 458 4480 460
rect 4492 458 4494 460
rect 4508 458 4510 460
rect 4522 458 4524 460
rect 4538 458 4540 460
rect 4552 458 4554 460
rect 4568 458 4570 460
rect 4582 458 4584 460
rect 4598 458 4600 460
rect 4612 458 4614 460
rect 4628 458 4630 460
rect 4642 458 4644 460
rect 4658 458 4660 460
rect 4672 458 4674 460
rect 4688 458 4690 460
rect 4702 458 4704 460
rect 4718 458 4720 460
rect 4732 458 4734 460
rect 4748 458 4750 460
rect 4762 458 4764 460
rect 4778 458 4780 460
rect 4792 458 4794 460
rect 4808 458 4810 460
rect 4822 458 4824 460
rect 4838 458 4840 460
rect 4852 458 4854 460
rect 4868 458 4870 460
rect 4882 458 4884 460
rect 4898 458 4900 460
rect 4912 458 4914 460
rect 4928 458 4930 460
rect 4942 458 4944 460
rect 4958 458 4960 460
rect 5042 458 5044 460
rect 5048 458 5050 460
rect 5062 458 5064 460
rect 5078 458 5080 460
rect 5092 458 5094 460
rect 5108 458 5110 460
rect 5122 458 5124 460
rect 5138 458 5140 460
rect 5152 458 5154 460
rect 5168 458 5170 460
rect 5182 458 5184 460
rect 5198 458 5200 460
rect 5212 458 5214 460
rect 5228 458 5230 460
rect 5242 458 5244 460
rect 5258 458 5260 460
rect 5272 458 5274 460
rect 5288 458 5290 460
rect 5302 458 5304 460
rect 5318 458 5320 460
rect 5332 458 5334 460
rect 5348 458 5350 460
rect 5362 458 5364 460
rect 5378 458 5380 460
rect 5392 458 5394 460
rect 5408 458 5410 460
rect 5422 458 5424 460
rect 5438 458 5440 460
rect 5452 458 5454 460
rect 5468 458 5470 460
rect 5482 458 5484 460
rect 5498 458 5500 460
rect 5512 458 5514 460
rect 5528 458 5530 460
rect 5542 458 5544 460
rect 5558 458 5560 460
rect 6240 459 6242 461
rect 6246 459 6248 461
rect 6260 459 6262 461
rect 6276 459 6278 461
rect 6290 459 6292 461
rect 6306 459 6308 461
rect 6320 459 6322 461
rect 6336 459 6338 461
rect 6350 459 6352 461
rect 6366 459 6368 461
rect 6380 459 6382 461
rect 6396 459 6398 461
rect 6410 459 6412 461
rect 6426 459 6428 461
rect 6440 459 6442 461
rect 6456 459 6458 461
rect 6470 459 6472 461
rect 6486 459 6488 461
rect 6500 459 6502 461
rect 6516 459 6518 461
rect 6530 459 6532 461
rect 6546 459 6548 461
rect 6560 459 6562 461
rect 6576 459 6578 461
rect 6590 459 6592 461
rect 6606 459 6608 461
rect 6620 459 6622 461
rect 6636 459 6638 461
rect 6650 459 6652 461
rect 6666 459 6668 461
rect 6680 459 6682 461
rect 6696 459 6698 461
rect 6710 459 6712 461
rect 6726 459 6728 461
rect 6740 459 6742 461
rect 6756 459 6758 461
rect 1748 454 1750 456
rect 1720 452 1722 454
rect 1746 452 1748 454
rect 1860 452 1862 454
rect 1718 450 1720 452
rect 1858 450 1860 452
rect 4470 450 4472 452
rect 4500 450 4502 452
rect 4530 450 4532 452
rect 4560 450 4562 452
rect 4590 450 4592 452
rect 4620 450 4622 452
rect 4650 450 4652 452
rect 4680 450 4682 452
rect 4710 450 4712 452
rect 4740 450 4742 452
rect 4770 450 4772 452
rect 4800 450 4802 452
rect 4830 450 4832 452
rect 4860 450 4862 452
rect 4890 450 4892 452
rect 4920 450 4922 452
rect 4950 450 4952 452
rect 5070 450 5072 452
rect 5100 450 5102 452
rect 5130 450 5132 452
rect 5160 450 5162 452
rect 5190 450 5192 452
rect 5220 450 5222 452
rect 5250 450 5252 452
rect 5280 450 5282 452
rect 5310 450 5312 452
rect 5340 450 5342 452
rect 5370 450 5372 452
rect 5400 450 5402 452
rect 5430 450 5432 452
rect 5460 450 5462 452
rect 5490 450 5492 452
rect 5520 450 5522 452
rect 5550 450 5552 452
rect 6268 451 6270 453
rect 6298 451 6300 453
rect 6328 451 6330 453
rect 6358 451 6360 453
rect 6388 451 6390 453
rect 6418 451 6420 453
rect 6448 451 6450 453
rect 6478 451 6480 453
rect 6508 451 6510 453
rect 6538 451 6540 453
rect 6568 451 6570 453
rect 6598 451 6600 453
rect 6628 451 6630 453
rect 6658 451 6660 453
rect 6688 451 6690 453
rect 6718 451 6720 453
rect 6748 451 6750 453
rect 4462 448 4464 450
rect 4468 448 4470 450
rect 4492 448 4494 450
rect 4498 448 4500 450
rect 4522 448 4524 450
rect 4528 448 4530 450
rect 4552 448 4554 450
rect 4558 448 4560 450
rect 4582 448 4584 450
rect 4588 448 4590 450
rect 4612 448 4614 450
rect 4618 448 4620 450
rect 4642 448 4644 450
rect 4648 448 4650 450
rect 4672 448 4674 450
rect 4678 448 4680 450
rect 4702 448 4704 450
rect 4708 448 4710 450
rect 4732 448 4734 450
rect 4738 448 4740 450
rect 4762 448 4764 450
rect 4768 448 4770 450
rect 4792 448 4794 450
rect 4798 448 4800 450
rect 4822 448 4824 450
rect 4828 448 4830 450
rect 4852 448 4854 450
rect 4858 448 4860 450
rect 4882 448 4884 450
rect 4888 448 4890 450
rect 4912 448 4914 450
rect 4918 448 4920 450
rect 4942 448 4944 450
rect 4948 448 4950 450
rect 5062 448 5064 450
rect 5068 448 5070 450
rect 5092 448 5094 450
rect 5098 448 5100 450
rect 5122 448 5124 450
rect 5128 448 5130 450
rect 5152 448 5154 450
rect 5158 448 5160 450
rect 5182 448 5184 450
rect 5188 448 5190 450
rect 5212 448 5214 450
rect 5218 448 5220 450
rect 5242 448 5244 450
rect 5248 448 5250 450
rect 5272 448 5274 450
rect 5278 448 5280 450
rect 5302 448 5304 450
rect 5308 448 5310 450
rect 5332 448 5334 450
rect 5338 448 5340 450
rect 5362 448 5364 450
rect 5368 448 5370 450
rect 5392 448 5394 450
rect 5398 448 5400 450
rect 5422 448 5424 450
rect 5428 448 5430 450
rect 5452 448 5454 450
rect 5458 448 5460 450
rect 5482 448 5484 450
rect 5488 448 5490 450
rect 5512 448 5514 450
rect 5518 448 5520 450
rect 5542 448 5544 450
rect 5548 448 5550 450
rect 6260 449 6262 451
rect 6266 449 6268 451
rect 6290 449 6292 451
rect 6296 449 6298 451
rect 6320 449 6322 451
rect 6326 449 6328 451
rect 6350 449 6352 451
rect 6356 449 6358 451
rect 6380 449 6382 451
rect 6386 449 6388 451
rect 6410 449 6412 451
rect 6416 449 6418 451
rect 6440 449 6442 451
rect 6446 449 6448 451
rect 6470 449 6472 451
rect 6476 449 6478 451
rect 6500 449 6502 451
rect 6506 449 6508 451
rect 6530 449 6532 451
rect 6536 449 6538 451
rect 6560 449 6562 451
rect 6566 449 6568 451
rect 6590 449 6592 451
rect 6596 449 6598 451
rect 6620 449 6622 451
rect 6626 449 6628 451
rect 6650 449 6652 451
rect 6656 449 6658 451
rect 6680 449 6682 451
rect 6686 449 6688 451
rect 6710 449 6712 451
rect 6716 449 6718 451
rect 6740 449 6742 451
rect 6746 449 6748 451
rect 4460 446 4462 448
rect 4490 446 4492 448
rect 4520 446 4522 448
rect 4550 446 4552 448
rect 4580 446 4582 448
rect 4610 446 4612 448
rect 4640 446 4642 448
rect 4670 446 4672 448
rect 4700 446 4702 448
rect 4730 446 4732 448
rect 4760 446 4762 448
rect 4790 446 4792 448
rect 4820 446 4822 448
rect 4850 446 4852 448
rect 4880 446 4882 448
rect 4910 446 4912 448
rect 4940 446 4942 448
rect 5060 446 5062 448
rect 5090 446 5092 448
rect 5120 446 5122 448
rect 5150 446 5152 448
rect 5180 446 5182 448
rect 5210 446 5212 448
rect 5240 446 5242 448
rect 5270 446 5272 448
rect 5300 446 5302 448
rect 5330 446 5332 448
rect 5360 446 5362 448
rect 5390 446 5392 448
rect 5420 446 5422 448
rect 5450 446 5452 448
rect 5480 446 5482 448
rect 5510 446 5512 448
rect 5540 446 5542 448
rect 6258 447 6260 449
rect 6288 447 6290 449
rect 6318 447 6320 449
rect 6348 447 6350 449
rect 6378 447 6380 449
rect 6408 447 6410 449
rect 6438 447 6440 449
rect 6468 447 6470 449
rect 6498 447 6500 449
rect 6528 447 6530 449
rect 6558 447 6560 449
rect 6588 447 6590 449
rect 6618 447 6620 449
rect 6648 447 6650 449
rect 6678 447 6680 449
rect 6708 447 6710 449
rect 6738 447 6740 449
rect 1738 444 1740 446
rect 1710 442 1712 444
rect 1736 442 1738 444
rect 1850 442 1852 444
rect 1708 440 1710 442
rect 1848 440 1850 442
rect 4460 440 4462 442
rect 4490 440 4492 442
rect 4520 440 4522 442
rect 4550 440 4552 442
rect 4580 440 4582 442
rect 4610 440 4612 442
rect 4640 440 4642 442
rect 4670 440 4672 442
rect 4700 440 4702 442
rect 4730 440 4732 442
rect 4760 440 4762 442
rect 4790 440 4792 442
rect 4820 440 4822 442
rect 4850 440 4852 442
rect 4880 440 4882 442
rect 4910 440 4912 442
rect 4940 440 4942 442
rect 5060 440 5062 442
rect 5090 440 5092 442
rect 5120 440 5122 442
rect 5150 440 5152 442
rect 5180 440 5182 442
rect 5210 440 5212 442
rect 5240 440 5242 442
rect 5270 440 5272 442
rect 5300 440 5302 442
rect 5330 440 5332 442
rect 5360 440 5362 442
rect 5390 440 5392 442
rect 5420 440 5422 442
rect 5450 440 5452 442
rect 5480 440 5482 442
rect 5510 440 5512 442
rect 5540 440 5542 442
rect 6258 441 6260 443
rect 6288 441 6290 443
rect 6318 441 6320 443
rect 6348 441 6350 443
rect 6378 441 6380 443
rect 6408 441 6410 443
rect 6438 441 6440 443
rect 6468 441 6470 443
rect 6498 441 6500 443
rect 6528 441 6530 443
rect 6558 441 6560 443
rect 6588 441 6590 443
rect 6618 441 6620 443
rect 6648 441 6650 443
rect 6678 441 6680 443
rect 6708 441 6710 443
rect 6738 441 6740 443
rect 4462 438 4464 440
rect 4468 438 4470 440
rect 4492 438 4494 440
rect 4498 438 4500 440
rect 4522 438 4524 440
rect 4528 438 4530 440
rect 4552 438 4554 440
rect 4558 438 4560 440
rect 4582 438 4584 440
rect 4588 438 4590 440
rect 4612 438 4614 440
rect 4618 438 4620 440
rect 4642 438 4644 440
rect 4648 438 4650 440
rect 4672 438 4674 440
rect 4678 438 4680 440
rect 4702 438 4704 440
rect 4708 438 4710 440
rect 4732 438 4734 440
rect 4738 438 4740 440
rect 4762 438 4764 440
rect 4768 438 4770 440
rect 4792 438 4794 440
rect 4798 438 4800 440
rect 4822 438 4824 440
rect 4828 438 4830 440
rect 4852 438 4854 440
rect 4858 438 4860 440
rect 4882 438 4884 440
rect 4888 438 4890 440
rect 4912 438 4914 440
rect 4918 438 4920 440
rect 4942 438 4944 440
rect 4948 438 4950 440
rect 5062 438 5064 440
rect 5068 438 5070 440
rect 5092 438 5094 440
rect 5098 438 5100 440
rect 5122 438 5124 440
rect 5128 438 5130 440
rect 5152 438 5154 440
rect 5158 438 5160 440
rect 5182 438 5184 440
rect 5188 438 5190 440
rect 5212 438 5214 440
rect 5218 438 5220 440
rect 5242 438 5244 440
rect 5248 438 5250 440
rect 5272 438 5274 440
rect 5278 438 5280 440
rect 5302 438 5304 440
rect 5308 438 5310 440
rect 5332 438 5334 440
rect 5338 438 5340 440
rect 5362 438 5364 440
rect 5368 438 5370 440
rect 5392 438 5394 440
rect 5398 438 5400 440
rect 5422 438 5424 440
rect 5428 438 5430 440
rect 5452 438 5454 440
rect 5458 438 5460 440
rect 5482 438 5484 440
rect 5488 438 5490 440
rect 5512 438 5514 440
rect 5518 438 5520 440
rect 5542 438 5544 440
rect 5548 438 5550 440
rect 6260 439 6262 441
rect 6266 439 6268 441
rect 6290 439 6292 441
rect 6296 439 6298 441
rect 6320 439 6322 441
rect 6326 439 6328 441
rect 6350 439 6352 441
rect 6356 439 6358 441
rect 6380 439 6382 441
rect 6386 439 6388 441
rect 6410 439 6412 441
rect 6416 439 6418 441
rect 6440 439 6442 441
rect 6446 439 6448 441
rect 6470 439 6472 441
rect 6476 439 6478 441
rect 6500 439 6502 441
rect 6506 439 6508 441
rect 6530 439 6532 441
rect 6536 439 6538 441
rect 6560 439 6562 441
rect 6566 439 6568 441
rect 6590 439 6592 441
rect 6596 439 6598 441
rect 6620 439 6622 441
rect 6626 439 6628 441
rect 6650 439 6652 441
rect 6656 439 6658 441
rect 6680 439 6682 441
rect 6686 439 6688 441
rect 6710 439 6712 441
rect 6716 439 6718 441
rect 6740 439 6742 441
rect 6746 439 6748 441
rect 4470 436 4472 438
rect 4500 436 4502 438
rect 4530 436 4532 438
rect 4560 436 4562 438
rect 4590 436 4592 438
rect 4620 436 4622 438
rect 4650 436 4652 438
rect 4680 436 4682 438
rect 4710 436 4712 438
rect 4740 436 4742 438
rect 4770 436 4772 438
rect 4800 436 4802 438
rect 4830 436 4832 438
rect 4860 436 4862 438
rect 4890 436 4892 438
rect 4920 436 4922 438
rect 4950 436 4952 438
rect 5070 436 5072 438
rect 5100 436 5102 438
rect 5130 436 5132 438
rect 5160 436 5162 438
rect 5190 436 5192 438
rect 5220 436 5222 438
rect 5250 436 5252 438
rect 5280 436 5282 438
rect 5310 436 5312 438
rect 5340 436 5342 438
rect 5370 436 5372 438
rect 5400 436 5402 438
rect 5430 436 5432 438
rect 5460 436 5462 438
rect 5490 436 5492 438
rect 5520 436 5522 438
rect 5550 436 5552 438
rect 6268 437 6270 439
rect 6298 437 6300 439
rect 6328 437 6330 439
rect 6358 437 6360 439
rect 6388 437 6390 439
rect 6418 437 6420 439
rect 6448 437 6450 439
rect 6478 437 6480 439
rect 6508 437 6510 439
rect 6538 437 6540 439
rect 6568 437 6570 439
rect 6598 437 6600 439
rect 6628 437 6630 439
rect 6658 437 6660 439
rect 6688 437 6690 439
rect 6718 437 6720 439
rect 6748 437 6750 439
rect 1728 434 1730 436
rect 1700 432 1702 434
rect 1726 432 1728 434
rect 1840 432 1842 434
rect 1698 430 1700 432
rect 1838 430 1840 432
rect 4470 430 4472 432
rect 4500 430 4502 432
rect 4530 430 4532 432
rect 4560 430 4562 432
rect 4590 430 4592 432
rect 4620 430 4622 432
rect 4650 430 4652 432
rect 4680 430 4682 432
rect 4710 430 4712 432
rect 4740 430 4742 432
rect 4770 430 4772 432
rect 4800 430 4802 432
rect 4830 430 4832 432
rect 4860 430 4862 432
rect 4890 430 4892 432
rect 4920 430 4922 432
rect 4950 430 4952 432
rect 5070 430 5072 432
rect 5100 430 5102 432
rect 5130 430 5132 432
rect 5160 430 5162 432
rect 5190 430 5192 432
rect 5220 430 5222 432
rect 5250 430 5252 432
rect 5280 430 5282 432
rect 5310 430 5312 432
rect 5340 430 5342 432
rect 5370 430 5372 432
rect 5400 430 5402 432
rect 5430 430 5432 432
rect 5460 430 5462 432
rect 5490 430 5492 432
rect 5520 430 5522 432
rect 5550 430 5552 432
rect 6268 431 6270 433
rect 6298 431 6300 433
rect 6328 431 6330 433
rect 6358 431 6360 433
rect 6388 431 6390 433
rect 6418 431 6420 433
rect 6448 431 6450 433
rect 6478 431 6480 433
rect 6508 431 6510 433
rect 6538 431 6540 433
rect 6568 431 6570 433
rect 6598 431 6600 433
rect 6628 431 6630 433
rect 6658 431 6660 433
rect 6688 431 6690 433
rect 6718 431 6720 433
rect 6748 431 6750 433
rect 4462 428 4464 430
rect 4468 428 4470 430
rect 4492 428 4494 430
rect 4498 428 4500 430
rect 4522 428 4524 430
rect 4528 428 4530 430
rect 4552 428 4554 430
rect 4558 428 4560 430
rect 4582 428 4584 430
rect 4588 428 4590 430
rect 4612 428 4614 430
rect 4618 428 4620 430
rect 4642 428 4644 430
rect 4648 428 4650 430
rect 4672 428 4674 430
rect 4678 428 4680 430
rect 4702 428 4704 430
rect 4708 428 4710 430
rect 4732 428 4734 430
rect 4738 428 4740 430
rect 4762 428 4764 430
rect 4768 428 4770 430
rect 4792 428 4794 430
rect 4798 428 4800 430
rect 4822 428 4824 430
rect 4828 428 4830 430
rect 4852 428 4854 430
rect 4858 428 4860 430
rect 4882 428 4884 430
rect 4888 428 4890 430
rect 4912 428 4914 430
rect 4918 428 4920 430
rect 4942 428 4944 430
rect 4948 428 4950 430
rect 5062 428 5064 430
rect 5068 428 5070 430
rect 5092 428 5094 430
rect 5098 428 5100 430
rect 5122 428 5124 430
rect 5128 428 5130 430
rect 5152 428 5154 430
rect 5158 428 5160 430
rect 5182 428 5184 430
rect 5188 428 5190 430
rect 5212 428 5214 430
rect 5218 428 5220 430
rect 5242 428 5244 430
rect 5248 428 5250 430
rect 5272 428 5274 430
rect 5278 428 5280 430
rect 5302 428 5304 430
rect 5308 428 5310 430
rect 5332 428 5334 430
rect 5338 428 5340 430
rect 5362 428 5364 430
rect 5368 428 5370 430
rect 5392 428 5394 430
rect 5398 428 5400 430
rect 5422 428 5424 430
rect 5428 428 5430 430
rect 5452 428 5454 430
rect 5458 428 5460 430
rect 5482 428 5484 430
rect 5488 428 5490 430
rect 5512 428 5514 430
rect 5518 428 5520 430
rect 5542 428 5544 430
rect 5548 428 5550 430
rect 6260 429 6262 431
rect 6266 429 6268 431
rect 6290 429 6292 431
rect 6296 429 6298 431
rect 6320 429 6322 431
rect 6326 429 6328 431
rect 6350 429 6352 431
rect 6356 429 6358 431
rect 6380 429 6382 431
rect 6386 429 6388 431
rect 6410 429 6412 431
rect 6416 429 6418 431
rect 6440 429 6442 431
rect 6446 429 6448 431
rect 6470 429 6472 431
rect 6476 429 6478 431
rect 6500 429 6502 431
rect 6506 429 6508 431
rect 6530 429 6532 431
rect 6536 429 6538 431
rect 6560 429 6562 431
rect 6566 429 6568 431
rect 6590 429 6592 431
rect 6596 429 6598 431
rect 6620 429 6622 431
rect 6626 429 6628 431
rect 6650 429 6652 431
rect 6656 429 6658 431
rect 6680 429 6682 431
rect 6686 429 6688 431
rect 6710 429 6712 431
rect 6716 429 6718 431
rect 6740 429 6742 431
rect 6746 429 6748 431
rect 4460 426 4462 428
rect 4490 426 4492 428
rect 4520 426 4522 428
rect 4550 426 4552 428
rect 4580 426 4582 428
rect 4610 426 4612 428
rect 4640 426 4642 428
rect 4670 426 4672 428
rect 4700 426 4702 428
rect 4730 426 4732 428
rect 4760 426 4762 428
rect 4790 426 4792 428
rect 4820 426 4822 428
rect 4850 426 4852 428
rect 4880 426 4882 428
rect 4910 426 4912 428
rect 4940 426 4942 428
rect 5060 426 5062 428
rect 5090 426 5092 428
rect 5120 426 5122 428
rect 5150 426 5152 428
rect 5180 426 5182 428
rect 5210 426 5212 428
rect 5240 426 5242 428
rect 5270 426 5272 428
rect 5300 426 5302 428
rect 5330 426 5332 428
rect 5360 426 5362 428
rect 5390 426 5392 428
rect 5420 426 5422 428
rect 5450 426 5452 428
rect 5480 426 5482 428
rect 5510 426 5512 428
rect 5540 426 5542 428
rect 6258 427 6260 429
rect 6288 427 6290 429
rect 6318 427 6320 429
rect 6348 427 6350 429
rect 6378 427 6380 429
rect 6408 427 6410 429
rect 6438 427 6440 429
rect 6468 427 6470 429
rect 6498 427 6500 429
rect 6528 427 6530 429
rect 6558 427 6560 429
rect 6588 427 6590 429
rect 6618 427 6620 429
rect 6648 427 6650 429
rect 6678 427 6680 429
rect 6708 427 6710 429
rect 6738 427 6740 429
rect 1718 424 1720 426
rect 1690 422 1692 424
rect 1716 422 1718 424
rect 3306 422 3308 424
rect 3692 422 3694 424
rect 3906 422 3908 424
rect 4292 422 4294 424
rect 1688 420 1690 422
rect 3304 420 3306 422
rect 3694 420 3696 422
rect 3904 420 3906 422
rect 4294 420 4296 422
rect 4460 420 4462 422
rect 4490 420 4492 422
rect 4520 420 4522 422
rect 4550 420 4552 422
rect 4580 420 4582 422
rect 4610 420 4612 422
rect 4640 420 4642 422
rect 4670 420 4672 422
rect 4700 420 4702 422
rect 4730 420 4732 422
rect 4760 420 4762 422
rect 4790 420 4792 422
rect 4820 420 4822 422
rect 4850 420 4852 422
rect 4880 420 4882 422
rect 4910 420 4912 422
rect 4940 420 4942 422
rect 5060 420 5062 422
rect 5090 420 5092 422
rect 5120 420 5122 422
rect 5150 420 5152 422
rect 5180 420 5182 422
rect 5210 420 5212 422
rect 5240 420 5242 422
rect 5270 420 5272 422
rect 5300 420 5302 422
rect 5330 420 5332 422
rect 5360 420 5362 422
rect 5390 420 5392 422
rect 5420 420 5422 422
rect 5450 420 5452 422
rect 5480 420 5482 422
rect 5510 420 5512 422
rect 5540 420 5542 422
rect 5706 420 5708 422
rect 6092 420 6094 422
rect 6258 421 6260 423
rect 6288 421 6290 423
rect 6318 421 6320 423
rect 6348 421 6350 423
rect 6378 421 6380 423
rect 6408 421 6410 423
rect 6438 421 6440 423
rect 6468 421 6470 423
rect 6498 421 6500 423
rect 6528 421 6530 423
rect 6558 421 6560 423
rect 6588 421 6590 423
rect 6618 421 6620 423
rect 6648 421 6650 423
rect 6678 421 6680 423
rect 6708 421 6710 423
rect 6738 421 6740 423
rect 4462 418 4464 420
rect 4468 418 4470 420
rect 4492 418 4494 420
rect 4498 418 4500 420
rect 4522 418 4524 420
rect 4528 418 4530 420
rect 4552 418 4554 420
rect 4558 418 4560 420
rect 4582 418 4584 420
rect 4588 418 4590 420
rect 4612 418 4614 420
rect 4618 418 4620 420
rect 4642 418 4644 420
rect 4648 418 4650 420
rect 4672 418 4674 420
rect 4678 418 4680 420
rect 4702 418 4704 420
rect 4708 418 4710 420
rect 4732 418 4734 420
rect 4738 418 4740 420
rect 4762 418 4764 420
rect 4768 418 4770 420
rect 4792 418 4794 420
rect 4798 418 4800 420
rect 4822 418 4824 420
rect 4828 418 4830 420
rect 4852 418 4854 420
rect 4858 418 4860 420
rect 4882 418 4884 420
rect 4888 418 4890 420
rect 4912 418 4914 420
rect 4918 418 4920 420
rect 4942 418 4944 420
rect 4948 418 4950 420
rect 5062 418 5064 420
rect 5068 418 5070 420
rect 5092 418 5094 420
rect 5098 418 5100 420
rect 5122 418 5124 420
rect 5128 418 5130 420
rect 5152 418 5154 420
rect 5158 418 5160 420
rect 5182 418 5184 420
rect 5188 418 5190 420
rect 5212 418 5214 420
rect 5218 418 5220 420
rect 5242 418 5244 420
rect 5248 418 5250 420
rect 5272 418 5274 420
rect 5278 418 5280 420
rect 5302 418 5304 420
rect 5308 418 5310 420
rect 5332 418 5334 420
rect 5338 418 5340 420
rect 5362 418 5364 420
rect 5368 418 5370 420
rect 5392 418 5394 420
rect 5398 418 5400 420
rect 5422 418 5424 420
rect 5428 418 5430 420
rect 5452 418 5454 420
rect 5458 418 5460 420
rect 5482 418 5484 420
rect 5488 418 5490 420
rect 5512 418 5514 420
rect 5518 418 5520 420
rect 5542 418 5544 420
rect 5548 418 5550 420
rect 5704 418 5706 420
rect 6094 418 6096 420
rect 6260 419 6262 421
rect 6266 419 6268 421
rect 6290 419 6292 421
rect 6296 419 6298 421
rect 6320 419 6322 421
rect 6326 419 6328 421
rect 6350 419 6352 421
rect 6356 419 6358 421
rect 6380 419 6382 421
rect 6386 419 6388 421
rect 6410 419 6412 421
rect 6416 419 6418 421
rect 6440 419 6442 421
rect 6446 419 6448 421
rect 6470 419 6472 421
rect 6476 419 6478 421
rect 6500 419 6502 421
rect 6506 419 6508 421
rect 6530 419 6532 421
rect 6536 419 6538 421
rect 6560 419 6562 421
rect 6566 419 6568 421
rect 6590 419 6592 421
rect 6596 419 6598 421
rect 6620 419 6622 421
rect 6626 419 6628 421
rect 6650 419 6652 421
rect 6656 419 6658 421
rect 6680 419 6682 421
rect 6686 419 6688 421
rect 6710 419 6712 421
rect 6716 419 6718 421
rect 6740 419 6742 421
rect 6746 419 6748 421
rect 4470 416 4472 418
rect 4500 416 4502 418
rect 4530 416 4532 418
rect 4560 416 4562 418
rect 4590 416 4592 418
rect 4620 416 4622 418
rect 4650 416 4652 418
rect 4680 416 4682 418
rect 4710 416 4712 418
rect 4740 416 4742 418
rect 4770 416 4772 418
rect 4800 416 4802 418
rect 4830 416 4832 418
rect 4860 416 4862 418
rect 4890 416 4892 418
rect 4920 416 4922 418
rect 4950 416 4952 418
rect 5070 416 5072 418
rect 5100 416 5102 418
rect 5130 416 5132 418
rect 5160 416 5162 418
rect 5190 416 5192 418
rect 5220 416 5222 418
rect 5250 416 5252 418
rect 5280 416 5282 418
rect 5310 416 5312 418
rect 5340 416 5342 418
rect 5370 416 5372 418
rect 5400 416 5402 418
rect 5430 416 5432 418
rect 5460 416 5462 418
rect 5490 416 5492 418
rect 5520 416 5522 418
rect 5550 416 5552 418
rect 6268 417 6270 419
rect 6298 417 6300 419
rect 6328 417 6330 419
rect 6358 417 6360 419
rect 6388 417 6390 419
rect 6418 417 6420 419
rect 6448 417 6450 419
rect 6478 417 6480 419
rect 6508 417 6510 419
rect 6538 417 6540 419
rect 6568 417 6570 419
rect 6598 417 6600 419
rect 6628 417 6630 419
rect 6658 417 6660 419
rect 6688 417 6690 419
rect 6718 417 6720 419
rect 6748 417 6750 419
rect 1708 414 1710 416
rect 1838 414 1840 416
rect 1680 412 1682 414
rect 1706 412 1708 414
rect 1840 412 1842 414
rect 1678 410 1680 412
rect 4470 410 4472 412
rect 4500 410 4502 412
rect 4530 410 4532 412
rect 4560 410 4562 412
rect 4590 410 4592 412
rect 4620 410 4622 412
rect 4650 410 4652 412
rect 4680 410 4682 412
rect 4710 410 4712 412
rect 4740 410 4742 412
rect 4770 410 4772 412
rect 4800 410 4802 412
rect 4830 410 4832 412
rect 4860 410 4862 412
rect 4890 410 4892 412
rect 4920 410 4922 412
rect 4950 410 4952 412
rect 5070 410 5072 412
rect 5100 410 5102 412
rect 5130 410 5132 412
rect 5160 410 5162 412
rect 5190 410 5192 412
rect 5220 410 5222 412
rect 5250 410 5252 412
rect 5280 410 5282 412
rect 5310 410 5312 412
rect 5340 410 5342 412
rect 5370 410 5372 412
rect 5400 410 5402 412
rect 5430 410 5432 412
rect 5460 410 5462 412
rect 5490 410 5492 412
rect 5520 410 5522 412
rect 5550 410 5552 412
rect 6268 411 6270 413
rect 6298 411 6300 413
rect 6328 411 6330 413
rect 6358 411 6360 413
rect 6388 411 6390 413
rect 6418 411 6420 413
rect 6448 411 6450 413
rect 6478 411 6480 413
rect 6508 411 6510 413
rect 6538 411 6540 413
rect 6568 411 6570 413
rect 6598 411 6600 413
rect 6628 411 6630 413
rect 6658 411 6660 413
rect 6688 411 6690 413
rect 6718 411 6720 413
rect 6748 411 6750 413
rect 4462 408 4464 410
rect 4468 408 4470 410
rect 4492 408 4494 410
rect 4498 408 4500 410
rect 4522 408 4524 410
rect 4528 408 4530 410
rect 4552 408 4554 410
rect 4558 408 4560 410
rect 4582 408 4584 410
rect 4588 408 4590 410
rect 4612 408 4614 410
rect 4618 408 4620 410
rect 4642 408 4644 410
rect 4648 408 4650 410
rect 4672 408 4674 410
rect 4678 408 4680 410
rect 4702 408 4704 410
rect 4708 408 4710 410
rect 4732 408 4734 410
rect 4738 408 4740 410
rect 4762 408 4764 410
rect 4768 408 4770 410
rect 4792 408 4794 410
rect 4798 408 4800 410
rect 4822 408 4824 410
rect 4828 408 4830 410
rect 4852 408 4854 410
rect 4858 408 4860 410
rect 4882 408 4884 410
rect 4888 408 4890 410
rect 4912 408 4914 410
rect 4918 408 4920 410
rect 4942 408 4944 410
rect 4948 408 4950 410
rect 5062 408 5064 410
rect 5068 408 5070 410
rect 5092 408 5094 410
rect 5098 408 5100 410
rect 5122 408 5124 410
rect 5128 408 5130 410
rect 5152 408 5154 410
rect 5158 408 5160 410
rect 5182 408 5184 410
rect 5188 408 5190 410
rect 5212 408 5214 410
rect 5218 408 5220 410
rect 5242 408 5244 410
rect 5248 408 5250 410
rect 5272 408 5274 410
rect 5278 408 5280 410
rect 5302 408 5304 410
rect 5308 408 5310 410
rect 5332 408 5334 410
rect 5338 408 5340 410
rect 5362 408 5364 410
rect 5368 408 5370 410
rect 5392 408 5394 410
rect 5398 408 5400 410
rect 5422 408 5424 410
rect 5428 408 5430 410
rect 5452 408 5454 410
rect 5458 408 5460 410
rect 5482 408 5484 410
rect 5488 408 5490 410
rect 5512 408 5514 410
rect 5518 408 5520 410
rect 5542 408 5544 410
rect 5548 408 5550 410
rect 6260 409 6262 411
rect 6266 409 6268 411
rect 6290 409 6292 411
rect 6296 409 6298 411
rect 6320 409 6322 411
rect 6326 409 6328 411
rect 6350 409 6352 411
rect 6356 409 6358 411
rect 6380 409 6382 411
rect 6386 409 6388 411
rect 6410 409 6412 411
rect 6416 409 6418 411
rect 6440 409 6442 411
rect 6446 409 6448 411
rect 6470 409 6472 411
rect 6476 409 6478 411
rect 6500 409 6502 411
rect 6506 409 6508 411
rect 6530 409 6532 411
rect 6536 409 6538 411
rect 6560 409 6562 411
rect 6566 409 6568 411
rect 6590 409 6592 411
rect 6596 409 6598 411
rect 6620 409 6622 411
rect 6626 409 6628 411
rect 6650 409 6652 411
rect 6656 409 6658 411
rect 6680 409 6682 411
rect 6686 409 6688 411
rect 6710 409 6712 411
rect 6716 409 6718 411
rect 6740 409 6742 411
rect 6746 409 6748 411
rect 4460 406 4462 408
rect 4490 406 4492 408
rect 4520 406 4522 408
rect 4550 406 4552 408
rect 4580 406 4582 408
rect 4610 406 4612 408
rect 4640 406 4642 408
rect 4670 406 4672 408
rect 4700 406 4702 408
rect 4730 406 4732 408
rect 4760 406 4762 408
rect 4790 406 4792 408
rect 4820 406 4822 408
rect 4850 406 4852 408
rect 4880 406 4882 408
rect 4910 406 4912 408
rect 4940 406 4942 408
rect 5060 406 5062 408
rect 5090 406 5092 408
rect 5120 406 5122 408
rect 5150 406 5152 408
rect 5180 406 5182 408
rect 5210 406 5212 408
rect 5240 406 5242 408
rect 5270 406 5272 408
rect 5300 406 5302 408
rect 5330 406 5332 408
rect 5360 406 5362 408
rect 5390 406 5392 408
rect 5420 406 5422 408
rect 5450 406 5452 408
rect 5480 406 5482 408
rect 5510 406 5512 408
rect 5540 406 5542 408
rect 6258 407 6260 409
rect 6288 407 6290 409
rect 6318 407 6320 409
rect 6348 407 6350 409
rect 6378 407 6380 409
rect 6408 407 6410 409
rect 6438 407 6440 409
rect 6468 407 6470 409
rect 6498 407 6500 409
rect 6528 407 6530 409
rect 6558 407 6560 409
rect 6588 407 6590 409
rect 6618 407 6620 409
rect 6648 407 6650 409
rect 6678 407 6680 409
rect 6708 407 6710 409
rect 6738 407 6740 409
rect 1698 404 1700 406
rect 1670 402 1672 404
rect 1696 402 1698 404
rect 1840 402 1842 404
rect 1668 400 1670 402
rect 1838 400 1840 402
rect 4460 400 4462 402
rect 4490 400 4492 402
rect 4520 400 4522 402
rect 4550 400 4552 402
rect 4580 400 4582 402
rect 4610 400 4612 402
rect 4640 400 4642 402
rect 4670 400 4672 402
rect 4700 400 4702 402
rect 4730 400 4732 402
rect 4760 400 4762 402
rect 4790 400 4792 402
rect 4820 400 4822 402
rect 4850 400 4852 402
rect 4880 400 4882 402
rect 4910 400 4912 402
rect 4940 400 4942 402
rect 5060 400 5062 402
rect 5090 400 5092 402
rect 5120 400 5122 402
rect 5150 400 5152 402
rect 5180 400 5182 402
rect 5210 400 5212 402
rect 5240 400 5242 402
rect 5270 400 5272 402
rect 5300 400 5302 402
rect 5330 400 5332 402
rect 5360 400 5362 402
rect 5390 400 5392 402
rect 5420 400 5422 402
rect 5450 400 5452 402
rect 5480 400 5482 402
rect 5510 400 5512 402
rect 5540 400 5542 402
rect 6258 401 6260 403
rect 6288 401 6290 403
rect 6318 401 6320 403
rect 6348 401 6350 403
rect 6378 401 6380 403
rect 6408 401 6410 403
rect 6438 401 6440 403
rect 6468 401 6470 403
rect 6498 401 6500 403
rect 6528 401 6530 403
rect 6558 401 6560 403
rect 6588 401 6590 403
rect 6618 401 6620 403
rect 6648 401 6650 403
rect 6678 401 6680 403
rect 6708 401 6710 403
rect 6738 401 6740 403
rect 4462 398 4464 400
rect 4468 398 4470 400
rect 4492 398 4494 400
rect 4498 398 4500 400
rect 4522 398 4524 400
rect 4528 398 4530 400
rect 4552 398 4554 400
rect 4558 398 4560 400
rect 4582 398 4584 400
rect 4588 398 4590 400
rect 4612 398 4614 400
rect 4618 398 4620 400
rect 4642 398 4644 400
rect 4648 398 4650 400
rect 4672 398 4674 400
rect 4678 398 4680 400
rect 4702 398 4704 400
rect 4708 398 4710 400
rect 4732 398 4734 400
rect 4738 398 4740 400
rect 4762 398 4764 400
rect 4768 398 4770 400
rect 4792 398 4794 400
rect 4798 398 4800 400
rect 4822 398 4824 400
rect 4828 398 4830 400
rect 4852 398 4854 400
rect 4858 398 4860 400
rect 4882 398 4884 400
rect 4888 398 4890 400
rect 4912 398 4914 400
rect 4918 398 4920 400
rect 4942 398 4944 400
rect 4948 398 4950 400
rect 5062 398 5064 400
rect 5068 398 5070 400
rect 5092 398 5094 400
rect 5098 398 5100 400
rect 5122 398 5124 400
rect 5128 398 5130 400
rect 5152 398 5154 400
rect 5158 398 5160 400
rect 5182 398 5184 400
rect 5188 398 5190 400
rect 5212 398 5214 400
rect 5218 398 5220 400
rect 5242 398 5244 400
rect 5248 398 5250 400
rect 5272 398 5274 400
rect 5278 398 5280 400
rect 5302 398 5304 400
rect 5308 398 5310 400
rect 5332 398 5334 400
rect 5338 398 5340 400
rect 5362 398 5364 400
rect 5368 398 5370 400
rect 5392 398 5394 400
rect 5398 398 5400 400
rect 5422 398 5424 400
rect 5428 398 5430 400
rect 5452 398 5454 400
rect 5458 398 5460 400
rect 5482 398 5484 400
rect 5488 398 5490 400
rect 5512 398 5514 400
rect 5518 398 5520 400
rect 5542 398 5544 400
rect 5548 398 5550 400
rect 6260 399 6262 401
rect 6266 399 6268 401
rect 6290 399 6292 401
rect 6296 399 6298 401
rect 6320 399 6322 401
rect 6326 399 6328 401
rect 6350 399 6352 401
rect 6356 399 6358 401
rect 6380 399 6382 401
rect 6386 399 6388 401
rect 6410 399 6412 401
rect 6416 399 6418 401
rect 6440 399 6442 401
rect 6446 399 6448 401
rect 6470 399 6472 401
rect 6476 399 6478 401
rect 6500 399 6502 401
rect 6506 399 6508 401
rect 6530 399 6532 401
rect 6536 399 6538 401
rect 6560 399 6562 401
rect 6566 399 6568 401
rect 6590 399 6592 401
rect 6596 399 6598 401
rect 6620 399 6622 401
rect 6626 399 6628 401
rect 6650 399 6652 401
rect 6656 399 6658 401
rect 6680 399 6682 401
rect 6686 399 6688 401
rect 6710 399 6712 401
rect 6716 399 6718 401
rect 6740 399 6742 401
rect 6746 399 6748 401
rect 4470 396 4472 398
rect 4500 396 4502 398
rect 4530 396 4532 398
rect 4560 396 4562 398
rect 4590 396 4592 398
rect 4620 396 4622 398
rect 4650 396 4652 398
rect 4680 396 4682 398
rect 4710 396 4712 398
rect 4740 396 4742 398
rect 4770 396 4772 398
rect 4800 396 4802 398
rect 4830 396 4832 398
rect 4860 396 4862 398
rect 4890 396 4892 398
rect 4920 396 4922 398
rect 4950 396 4952 398
rect 5070 396 5072 398
rect 5100 396 5102 398
rect 5130 396 5132 398
rect 5160 396 5162 398
rect 5190 396 5192 398
rect 5220 396 5222 398
rect 5250 396 5252 398
rect 5280 396 5282 398
rect 5310 396 5312 398
rect 5340 396 5342 398
rect 5370 396 5372 398
rect 5400 396 5402 398
rect 5430 396 5432 398
rect 5460 396 5462 398
rect 5490 396 5492 398
rect 5520 396 5522 398
rect 5550 396 5552 398
rect 6268 397 6270 399
rect 6298 397 6300 399
rect 6328 397 6330 399
rect 6358 397 6360 399
rect 6388 397 6390 399
rect 6418 397 6420 399
rect 6448 397 6450 399
rect 6478 397 6480 399
rect 6508 397 6510 399
rect 6538 397 6540 399
rect 6568 397 6570 399
rect 6598 397 6600 399
rect 6628 397 6630 399
rect 6658 397 6660 399
rect 6688 397 6690 399
rect 6718 397 6720 399
rect 6748 397 6750 399
rect 1688 394 1690 396
rect 1660 392 1662 394
rect 1686 392 1688 394
rect 1830 392 1832 394
rect 1658 390 1660 392
rect 1828 390 1830 392
rect 4500 390 4502 392
rect 4920 390 4922 392
rect 4950 390 4952 392
rect 5100 390 5102 392
rect 5520 390 5522 392
rect 5550 390 5552 392
rect 6298 391 6300 393
rect 6718 391 6720 393
rect 6748 391 6750 393
rect 4498 388 4500 390
rect 4918 388 4920 390
rect 4942 388 4944 390
rect 4948 388 4950 390
rect 5098 388 5100 390
rect 5518 388 5520 390
rect 5542 388 5544 390
rect 5548 388 5550 390
rect 6296 389 6298 391
rect 6716 389 6718 391
rect 6740 389 6742 391
rect 6746 389 6748 391
rect 4940 386 4942 388
rect 5540 386 5542 388
rect 6738 387 6740 389
rect 1678 384 1680 386
rect 1650 382 1652 384
rect 1676 382 1678 384
rect 1820 382 1822 384
rect 1648 380 1650 382
rect 1818 380 1820 382
rect 4940 380 4942 382
rect 5540 380 5542 382
rect 6738 381 6740 383
rect 4498 378 4500 380
rect 4918 378 4920 380
rect 4942 378 4944 380
rect 4948 378 4950 380
rect 5098 378 5100 380
rect 5518 378 5520 380
rect 5542 378 5544 380
rect 5548 378 5550 380
rect 6296 379 6298 381
rect 6716 379 6718 381
rect 6740 379 6742 381
rect 6746 379 6748 381
rect 4500 376 4502 378
rect 4920 376 4922 378
rect 4950 376 4952 378
rect 5100 376 5102 378
rect 5520 376 5522 378
rect 5550 376 5552 378
rect 6298 377 6300 379
rect 6718 377 6720 379
rect 6748 377 6750 379
rect 1668 374 1670 376
rect 1640 372 1642 374
rect 1666 372 1668 374
rect 1810 372 1812 374
rect 1638 370 1640 372
rect 1808 370 1810 372
rect 4470 370 4472 372
rect 4500 370 4502 372
rect 4530 370 4532 372
rect 4560 370 4562 372
rect 4590 370 4592 372
rect 4620 370 4622 372
rect 4650 370 4652 372
rect 4680 370 4682 372
rect 4710 370 4712 372
rect 4740 370 4742 372
rect 4770 370 4772 372
rect 4800 370 4802 372
rect 4830 370 4832 372
rect 4860 370 4862 372
rect 4890 370 4892 372
rect 4920 370 4922 372
rect 4950 370 4952 372
rect 5070 370 5072 372
rect 5100 370 5102 372
rect 5130 370 5132 372
rect 5160 370 5162 372
rect 5190 370 5192 372
rect 5220 370 5222 372
rect 5250 370 5252 372
rect 5280 370 5282 372
rect 5310 370 5312 372
rect 5340 370 5342 372
rect 5370 370 5372 372
rect 5400 370 5402 372
rect 5430 370 5432 372
rect 5460 370 5462 372
rect 5490 370 5492 372
rect 5520 370 5522 372
rect 5550 370 5552 372
rect 6268 371 6270 373
rect 6298 371 6300 373
rect 6328 371 6330 373
rect 6358 371 6360 373
rect 6388 371 6390 373
rect 6418 371 6420 373
rect 6448 371 6450 373
rect 6478 371 6480 373
rect 6508 371 6510 373
rect 6538 371 6540 373
rect 6568 371 6570 373
rect 6598 371 6600 373
rect 6628 371 6630 373
rect 6658 371 6660 373
rect 6688 371 6690 373
rect 6718 371 6720 373
rect 6748 371 6750 373
rect 4462 368 4464 370
rect 4468 368 4470 370
rect 4492 368 4494 370
rect 4498 368 4500 370
rect 4522 368 4524 370
rect 4528 368 4530 370
rect 4552 368 4554 370
rect 4558 368 4560 370
rect 4582 368 4584 370
rect 4588 368 4590 370
rect 4612 368 4614 370
rect 4618 368 4620 370
rect 4642 368 4644 370
rect 4648 368 4650 370
rect 4672 368 4674 370
rect 4678 368 4680 370
rect 4702 368 4704 370
rect 4708 368 4710 370
rect 4732 368 4734 370
rect 4738 368 4740 370
rect 4762 368 4764 370
rect 4768 368 4770 370
rect 4792 368 4794 370
rect 4798 368 4800 370
rect 4822 368 4824 370
rect 4828 368 4830 370
rect 4852 368 4854 370
rect 4858 368 4860 370
rect 4882 368 4884 370
rect 4888 368 4890 370
rect 4912 368 4914 370
rect 4918 368 4920 370
rect 4942 368 4944 370
rect 4948 368 4950 370
rect 5062 368 5064 370
rect 5068 368 5070 370
rect 5092 368 5094 370
rect 5098 368 5100 370
rect 5122 368 5124 370
rect 5128 368 5130 370
rect 5152 368 5154 370
rect 5158 368 5160 370
rect 5182 368 5184 370
rect 5188 368 5190 370
rect 5212 368 5214 370
rect 5218 368 5220 370
rect 5242 368 5244 370
rect 5248 368 5250 370
rect 5272 368 5274 370
rect 5278 368 5280 370
rect 5302 368 5304 370
rect 5308 368 5310 370
rect 5332 368 5334 370
rect 5338 368 5340 370
rect 5362 368 5364 370
rect 5368 368 5370 370
rect 5392 368 5394 370
rect 5398 368 5400 370
rect 5422 368 5424 370
rect 5428 368 5430 370
rect 5452 368 5454 370
rect 5458 368 5460 370
rect 5482 368 5484 370
rect 5488 368 5490 370
rect 5512 368 5514 370
rect 5518 368 5520 370
rect 5542 368 5544 370
rect 5548 368 5550 370
rect 6260 369 6262 371
rect 6266 369 6268 371
rect 6290 369 6292 371
rect 6296 369 6298 371
rect 6320 369 6322 371
rect 6326 369 6328 371
rect 6350 369 6352 371
rect 6356 369 6358 371
rect 6380 369 6382 371
rect 6386 369 6388 371
rect 6410 369 6412 371
rect 6416 369 6418 371
rect 6440 369 6442 371
rect 6446 369 6448 371
rect 6470 369 6472 371
rect 6476 369 6478 371
rect 6500 369 6502 371
rect 6506 369 6508 371
rect 6530 369 6532 371
rect 6536 369 6538 371
rect 6560 369 6562 371
rect 6566 369 6568 371
rect 6590 369 6592 371
rect 6596 369 6598 371
rect 6620 369 6622 371
rect 6626 369 6628 371
rect 6650 369 6652 371
rect 6656 369 6658 371
rect 6680 369 6682 371
rect 6686 369 6688 371
rect 6710 369 6712 371
rect 6716 369 6718 371
rect 6740 369 6742 371
rect 6746 369 6748 371
rect 4460 366 4462 368
rect 4490 366 4492 368
rect 4520 366 4522 368
rect 4550 366 4552 368
rect 4580 366 4582 368
rect 4610 366 4612 368
rect 4640 366 4642 368
rect 4670 366 4672 368
rect 4700 366 4702 368
rect 4730 366 4732 368
rect 4760 366 4762 368
rect 4790 366 4792 368
rect 4820 366 4822 368
rect 4850 366 4852 368
rect 4880 366 4882 368
rect 4910 366 4912 368
rect 4940 366 4942 368
rect 5060 366 5062 368
rect 5090 366 5092 368
rect 5120 366 5122 368
rect 5150 366 5152 368
rect 5180 366 5182 368
rect 5210 366 5212 368
rect 5240 366 5242 368
rect 5270 366 5272 368
rect 5300 366 5302 368
rect 5330 366 5332 368
rect 5360 366 5362 368
rect 5390 366 5392 368
rect 5420 366 5422 368
rect 5450 366 5452 368
rect 5480 366 5482 368
rect 5510 366 5512 368
rect 5540 366 5542 368
rect 6258 367 6260 369
rect 6288 367 6290 369
rect 6318 367 6320 369
rect 6348 367 6350 369
rect 6378 367 6380 369
rect 6408 367 6410 369
rect 6438 367 6440 369
rect 6468 367 6470 369
rect 6498 367 6500 369
rect 6528 367 6530 369
rect 6558 367 6560 369
rect 6588 367 6590 369
rect 6618 367 6620 369
rect 6648 367 6650 369
rect 6678 367 6680 369
rect 6708 367 6710 369
rect 6738 367 6740 369
rect 1658 364 1660 366
rect 1630 362 1632 364
rect 1656 362 1658 364
rect 1800 362 1802 364
rect 1628 360 1630 362
rect 1798 360 1800 362
rect 4460 360 4462 362
rect 4490 360 4492 362
rect 4520 360 4522 362
rect 4550 360 4552 362
rect 4580 360 4582 362
rect 4610 360 4612 362
rect 4640 360 4642 362
rect 4670 360 4672 362
rect 4700 360 4702 362
rect 4730 360 4732 362
rect 4760 360 4762 362
rect 4790 360 4792 362
rect 4820 360 4822 362
rect 4850 360 4852 362
rect 4880 360 4882 362
rect 4910 360 4912 362
rect 4940 360 4942 362
rect 5060 360 5062 362
rect 5090 360 5092 362
rect 5120 360 5122 362
rect 5150 360 5152 362
rect 5180 360 5182 362
rect 5210 360 5212 362
rect 5240 360 5242 362
rect 5270 360 5272 362
rect 5300 360 5302 362
rect 5330 360 5332 362
rect 5360 360 5362 362
rect 5390 360 5392 362
rect 5420 360 5422 362
rect 5450 360 5452 362
rect 5480 360 5482 362
rect 5510 360 5512 362
rect 5540 360 5542 362
rect 6258 361 6260 363
rect 6288 361 6290 363
rect 6318 361 6320 363
rect 6348 361 6350 363
rect 6378 361 6380 363
rect 6408 361 6410 363
rect 6438 361 6440 363
rect 6468 361 6470 363
rect 6498 361 6500 363
rect 6528 361 6530 363
rect 6558 361 6560 363
rect 6588 361 6590 363
rect 6618 361 6620 363
rect 6648 361 6650 363
rect 6678 361 6680 363
rect 6708 361 6710 363
rect 6738 361 6740 363
rect 3304 358 3306 360
rect 3694 358 3696 360
rect 3904 358 3906 360
rect 4294 358 4296 360
rect 4462 358 4464 360
rect 4468 358 4470 360
rect 4492 358 4494 360
rect 4498 358 4500 360
rect 4522 358 4524 360
rect 4528 358 4530 360
rect 4552 358 4554 360
rect 4558 358 4560 360
rect 4582 358 4584 360
rect 4588 358 4590 360
rect 4612 358 4614 360
rect 4618 358 4620 360
rect 4642 358 4644 360
rect 4648 358 4650 360
rect 4672 358 4674 360
rect 4678 358 4680 360
rect 4702 358 4704 360
rect 4708 358 4710 360
rect 4732 358 4734 360
rect 4738 358 4740 360
rect 4762 358 4764 360
rect 4768 358 4770 360
rect 4792 358 4794 360
rect 4798 358 4800 360
rect 4822 358 4824 360
rect 4828 358 4830 360
rect 4852 358 4854 360
rect 4858 358 4860 360
rect 4882 358 4884 360
rect 4888 358 4890 360
rect 4912 358 4914 360
rect 4918 358 4920 360
rect 4942 358 4944 360
rect 4948 358 4950 360
rect 5062 358 5064 360
rect 5068 358 5070 360
rect 5092 358 5094 360
rect 5098 358 5100 360
rect 5122 358 5124 360
rect 5128 358 5130 360
rect 5152 358 5154 360
rect 5158 358 5160 360
rect 5182 358 5184 360
rect 5188 358 5190 360
rect 5212 358 5214 360
rect 5218 358 5220 360
rect 5242 358 5244 360
rect 5248 358 5250 360
rect 5272 358 5274 360
rect 5278 358 5280 360
rect 5302 358 5304 360
rect 5308 358 5310 360
rect 5332 358 5334 360
rect 5338 358 5340 360
rect 5362 358 5364 360
rect 5368 358 5370 360
rect 5392 358 5394 360
rect 5398 358 5400 360
rect 5422 358 5424 360
rect 5428 358 5430 360
rect 5452 358 5454 360
rect 5458 358 5460 360
rect 5482 358 5484 360
rect 5488 358 5490 360
rect 5512 358 5514 360
rect 5518 358 5520 360
rect 5542 358 5544 360
rect 5548 358 5550 360
rect 6260 359 6262 361
rect 6266 359 6268 361
rect 6290 359 6292 361
rect 6296 359 6298 361
rect 6320 359 6322 361
rect 6326 359 6328 361
rect 6350 359 6352 361
rect 6356 359 6358 361
rect 6380 359 6382 361
rect 6386 359 6388 361
rect 6410 359 6412 361
rect 6416 359 6418 361
rect 6440 359 6442 361
rect 6446 359 6448 361
rect 6470 359 6472 361
rect 6476 359 6478 361
rect 6500 359 6502 361
rect 6506 359 6508 361
rect 6530 359 6532 361
rect 6536 359 6538 361
rect 6560 359 6562 361
rect 6566 359 6568 361
rect 6590 359 6592 361
rect 6596 359 6598 361
rect 6620 359 6622 361
rect 6626 359 6628 361
rect 6650 359 6652 361
rect 6656 359 6658 361
rect 6680 359 6682 361
rect 6686 359 6688 361
rect 6710 359 6712 361
rect 6716 359 6718 361
rect 6740 359 6742 361
rect 6746 359 6748 361
rect 3306 356 3308 358
rect 3692 356 3694 358
rect 3906 356 3908 358
rect 4292 356 4294 358
rect 4470 356 4472 358
rect 4500 356 4502 358
rect 4530 356 4532 358
rect 4560 356 4562 358
rect 4590 356 4592 358
rect 4620 356 4622 358
rect 4650 356 4652 358
rect 4680 356 4682 358
rect 4710 356 4712 358
rect 4740 356 4742 358
rect 4770 356 4772 358
rect 4800 356 4802 358
rect 4830 356 4832 358
rect 4860 356 4862 358
rect 4890 356 4892 358
rect 4920 356 4922 358
rect 4950 356 4952 358
rect 5070 356 5072 358
rect 5100 356 5102 358
rect 5130 356 5132 358
rect 5160 356 5162 358
rect 5190 356 5192 358
rect 5220 356 5222 358
rect 5250 356 5252 358
rect 5280 356 5282 358
rect 5310 356 5312 358
rect 5340 356 5342 358
rect 5370 356 5372 358
rect 5400 356 5402 358
rect 5430 356 5432 358
rect 5460 356 5462 358
rect 5490 356 5492 358
rect 5520 356 5522 358
rect 5550 356 5552 358
rect 5704 356 5706 358
rect 6094 356 6096 358
rect 6268 357 6270 359
rect 6298 357 6300 359
rect 6328 357 6330 359
rect 6358 357 6360 359
rect 6388 357 6390 359
rect 6418 357 6420 359
rect 6448 357 6450 359
rect 6478 357 6480 359
rect 6508 357 6510 359
rect 6538 357 6540 359
rect 6568 357 6570 359
rect 6598 357 6600 359
rect 6628 357 6630 359
rect 6658 357 6660 359
rect 6688 357 6690 359
rect 6718 357 6720 359
rect 6748 357 6750 359
rect 1648 354 1650 356
rect 5706 354 5708 356
rect 6092 354 6094 356
rect 1620 352 1622 354
rect 1646 352 1648 354
rect 1790 352 1792 354
rect 1618 350 1620 352
rect 1788 350 1790 352
rect 4470 350 4472 352
rect 4500 350 4502 352
rect 4530 350 4532 352
rect 4560 350 4562 352
rect 4590 350 4592 352
rect 4620 350 4622 352
rect 4650 350 4652 352
rect 4680 350 4682 352
rect 4710 350 4712 352
rect 4740 350 4742 352
rect 4770 350 4772 352
rect 4800 350 4802 352
rect 4830 350 4832 352
rect 4860 350 4862 352
rect 4890 350 4892 352
rect 4920 350 4922 352
rect 4950 350 4952 352
rect 5070 350 5072 352
rect 5100 350 5102 352
rect 5130 350 5132 352
rect 5160 350 5162 352
rect 5190 350 5192 352
rect 5220 350 5222 352
rect 5250 350 5252 352
rect 5280 350 5282 352
rect 5310 350 5312 352
rect 5340 350 5342 352
rect 5370 350 5372 352
rect 5400 350 5402 352
rect 5430 350 5432 352
rect 5460 350 5462 352
rect 5490 350 5492 352
rect 5520 350 5522 352
rect 5550 350 5552 352
rect 6268 351 6270 353
rect 6298 351 6300 353
rect 6328 351 6330 353
rect 6358 351 6360 353
rect 6388 351 6390 353
rect 6418 351 6420 353
rect 6448 351 6450 353
rect 6478 351 6480 353
rect 6508 351 6510 353
rect 6538 351 6540 353
rect 6568 351 6570 353
rect 6598 351 6600 353
rect 6628 351 6630 353
rect 6658 351 6660 353
rect 6688 351 6690 353
rect 6718 351 6720 353
rect 6748 351 6750 353
rect 4462 348 4464 350
rect 4468 348 4470 350
rect 4492 348 4494 350
rect 4498 348 4500 350
rect 4522 348 4524 350
rect 4528 348 4530 350
rect 4552 348 4554 350
rect 4558 348 4560 350
rect 4582 348 4584 350
rect 4588 348 4590 350
rect 4612 348 4614 350
rect 4618 348 4620 350
rect 4642 348 4644 350
rect 4648 348 4650 350
rect 4672 348 4674 350
rect 4678 348 4680 350
rect 4702 348 4704 350
rect 4708 348 4710 350
rect 4732 348 4734 350
rect 4738 348 4740 350
rect 4762 348 4764 350
rect 4768 348 4770 350
rect 4792 348 4794 350
rect 4798 348 4800 350
rect 4822 348 4824 350
rect 4828 348 4830 350
rect 4852 348 4854 350
rect 4858 348 4860 350
rect 4882 348 4884 350
rect 4888 348 4890 350
rect 4912 348 4914 350
rect 4918 348 4920 350
rect 4942 348 4944 350
rect 4948 348 4950 350
rect 5062 348 5064 350
rect 5068 348 5070 350
rect 5092 348 5094 350
rect 5098 348 5100 350
rect 5122 348 5124 350
rect 5128 348 5130 350
rect 5152 348 5154 350
rect 5158 348 5160 350
rect 5182 348 5184 350
rect 5188 348 5190 350
rect 5212 348 5214 350
rect 5218 348 5220 350
rect 5242 348 5244 350
rect 5248 348 5250 350
rect 5272 348 5274 350
rect 5278 348 5280 350
rect 5302 348 5304 350
rect 5308 348 5310 350
rect 5332 348 5334 350
rect 5338 348 5340 350
rect 5362 348 5364 350
rect 5368 348 5370 350
rect 5392 348 5394 350
rect 5398 348 5400 350
rect 5422 348 5424 350
rect 5428 348 5430 350
rect 5452 348 5454 350
rect 5458 348 5460 350
rect 5482 348 5484 350
rect 5488 348 5490 350
rect 5512 348 5514 350
rect 5518 348 5520 350
rect 5542 348 5544 350
rect 5548 348 5550 350
rect 6260 349 6262 351
rect 6266 349 6268 351
rect 6290 349 6292 351
rect 6296 349 6298 351
rect 6320 349 6322 351
rect 6326 349 6328 351
rect 6350 349 6352 351
rect 6356 349 6358 351
rect 6380 349 6382 351
rect 6386 349 6388 351
rect 6410 349 6412 351
rect 6416 349 6418 351
rect 6440 349 6442 351
rect 6446 349 6448 351
rect 6470 349 6472 351
rect 6476 349 6478 351
rect 6500 349 6502 351
rect 6506 349 6508 351
rect 6530 349 6532 351
rect 6536 349 6538 351
rect 6560 349 6562 351
rect 6566 349 6568 351
rect 6590 349 6592 351
rect 6596 349 6598 351
rect 6620 349 6622 351
rect 6626 349 6628 351
rect 6650 349 6652 351
rect 6656 349 6658 351
rect 6680 349 6682 351
rect 6686 349 6688 351
rect 6710 349 6712 351
rect 6716 349 6718 351
rect 6740 349 6742 351
rect 6746 349 6748 351
rect 4460 346 4462 348
rect 4490 346 4492 348
rect 4520 346 4522 348
rect 4550 346 4552 348
rect 4580 346 4582 348
rect 4610 346 4612 348
rect 4640 346 4642 348
rect 4670 346 4672 348
rect 4700 346 4702 348
rect 4730 346 4732 348
rect 4760 346 4762 348
rect 4790 346 4792 348
rect 4820 346 4822 348
rect 4850 346 4852 348
rect 4880 346 4882 348
rect 4910 346 4912 348
rect 4940 346 4942 348
rect 5060 346 5062 348
rect 5090 346 5092 348
rect 5120 346 5122 348
rect 5150 346 5152 348
rect 5180 346 5182 348
rect 5210 346 5212 348
rect 5240 346 5242 348
rect 5270 346 5272 348
rect 5300 346 5302 348
rect 5330 346 5332 348
rect 5360 346 5362 348
rect 5390 346 5392 348
rect 5420 346 5422 348
rect 5450 346 5452 348
rect 5480 346 5482 348
rect 5510 346 5512 348
rect 5540 346 5542 348
rect 6258 347 6260 349
rect 6288 347 6290 349
rect 6318 347 6320 349
rect 6348 347 6350 349
rect 6378 347 6380 349
rect 6408 347 6410 349
rect 6438 347 6440 349
rect 6468 347 6470 349
rect 6498 347 6500 349
rect 6528 347 6530 349
rect 6558 347 6560 349
rect 6588 347 6590 349
rect 6618 347 6620 349
rect 6648 347 6650 349
rect 6678 347 6680 349
rect 6708 347 6710 349
rect 6738 347 6740 349
rect 1638 344 1640 346
rect 1610 342 1612 344
rect 1636 342 1638 344
rect 1780 342 1782 344
rect 1608 340 1610 342
rect 1778 340 1780 342
rect 4460 340 4462 342
rect 4490 340 4492 342
rect 4520 340 4522 342
rect 4550 340 4552 342
rect 4580 340 4582 342
rect 4610 340 4612 342
rect 4640 340 4642 342
rect 4670 340 4672 342
rect 4700 340 4702 342
rect 4730 340 4732 342
rect 4760 340 4762 342
rect 4790 340 4792 342
rect 4820 340 4822 342
rect 4850 340 4852 342
rect 4880 340 4882 342
rect 4910 340 4912 342
rect 4940 340 4942 342
rect 5060 340 5062 342
rect 5090 340 5092 342
rect 5120 340 5122 342
rect 5150 340 5152 342
rect 5180 340 5182 342
rect 5210 340 5212 342
rect 5240 340 5242 342
rect 5270 340 5272 342
rect 5300 340 5302 342
rect 5330 340 5332 342
rect 5360 340 5362 342
rect 5390 340 5392 342
rect 5420 340 5422 342
rect 5450 340 5452 342
rect 5480 340 5482 342
rect 5510 340 5512 342
rect 5540 340 5542 342
rect 6258 341 6260 343
rect 6288 341 6290 343
rect 6318 341 6320 343
rect 6348 341 6350 343
rect 6378 341 6380 343
rect 6408 341 6410 343
rect 6438 341 6440 343
rect 6468 341 6470 343
rect 6498 341 6500 343
rect 6528 341 6530 343
rect 6558 341 6560 343
rect 6588 341 6590 343
rect 6618 341 6620 343
rect 6648 341 6650 343
rect 6678 341 6680 343
rect 6708 341 6710 343
rect 6738 341 6740 343
rect 4462 338 4464 340
rect 4468 338 4470 340
rect 4492 338 4494 340
rect 4498 338 4500 340
rect 4522 338 4524 340
rect 4528 338 4530 340
rect 4552 338 4554 340
rect 4558 338 4560 340
rect 4582 338 4584 340
rect 4588 338 4590 340
rect 4612 338 4614 340
rect 4618 338 4620 340
rect 4642 338 4644 340
rect 4648 338 4650 340
rect 4672 338 4674 340
rect 4678 338 4680 340
rect 4702 338 4704 340
rect 4708 338 4710 340
rect 4732 338 4734 340
rect 4738 338 4740 340
rect 4762 338 4764 340
rect 4768 338 4770 340
rect 4792 338 4794 340
rect 4798 338 4800 340
rect 4822 338 4824 340
rect 4828 338 4830 340
rect 4852 338 4854 340
rect 4858 338 4860 340
rect 4882 338 4884 340
rect 4888 338 4890 340
rect 4912 338 4914 340
rect 4918 338 4920 340
rect 4942 338 4944 340
rect 4948 338 4950 340
rect 5062 338 5064 340
rect 5068 338 5070 340
rect 5092 338 5094 340
rect 5098 338 5100 340
rect 5122 338 5124 340
rect 5128 338 5130 340
rect 5152 338 5154 340
rect 5158 338 5160 340
rect 5182 338 5184 340
rect 5188 338 5190 340
rect 5212 338 5214 340
rect 5218 338 5220 340
rect 5242 338 5244 340
rect 5248 338 5250 340
rect 5272 338 5274 340
rect 5278 338 5280 340
rect 5302 338 5304 340
rect 5308 338 5310 340
rect 5332 338 5334 340
rect 5338 338 5340 340
rect 5362 338 5364 340
rect 5368 338 5370 340
rect 5392 338 5394 340
rect 5398 338 5400 340
rect 5422 338 5424 340
rect 5428 338 5430 340
rect 5452 338 5454 340
rect 5458 338 5460 340
rect 5482 338 5484 340
rect 5488 338 5490 340
rect 5512 338 5514 340
rect 5518 338 5520 340
rect 5542 338 5544 340
rect 5548 338 5550 340
rect 6260 339 6262 341
rect 6266 339 6268 341
rect 6290 339 6292 341
rect 6296 339 6298 341
rect 6320 339 6322 341
rect 6326 339 6328 341
rect 6350 339 6352 341
rect 6356 339 6358 341
rect 6380 339 6382 341
rect 6386 339 6388 341
rect 6410 339 6412 341
rect 6416 339 6418 341
rect 6440 339 6442 341
rect 6446 339 6448 341
rect 6470 339 6472 341
rect 6476 339 6478 341
rect 6500 339 6502 341
rect 6506 339 6508 341
rect 6530 339 6532 341
rect 6536 339 6538 341
rect 6560 339 6562 341
rect 6566 339 6568 341
rect 6590 339 6592 341
rect 6596 339 6598 341
rect 6620 339 6622 341
rect 6626 339 6628 341
rect 6650 339 6652 341
rect 6656 339 6658 341
rect 6680 339 6682 341
rect 6686 339 6688 341
rect 6710 339 6712 341
rect 6716 339 6718 341
rect 6740 339 6742 341
rect 6746 339 6748 341
rect 4470 336 4472 338
rect 4500 336 4502 338
rect 4530 336 4532 338
rect 4560 336 4562 338
rect 4590 336 4592 338
rect 4620 336 4622 338
rect 4650 336 4652 338
rect 4680 336 4682 338
rect 4710 336 4712 338
rect 4740 336 4742 338
rect 4770 336 4772 338
rect 4800 336 4802 338
rect 4830 336 4832 338
rect 4860 336 4862 338
rect 4890 336 4892 338
rect 4920 336 4922 338
rect 4950 336 4952 338
rect 5070 336 5072 338
rect 5100 336 5102 338
rect 5130 336 5132 338
rect 5160 336 5162 338
rect 5190 336 5192 338
rect 5220 336 5222 338
rect 5250 336 5252 338
rect 5280 336 5282 338
rect 5310 336 5312 338
rect 5340 336 5342 338
rect 5370 336 5372 338
rect 5400 336 5402 338
rect 5430 336 5432 338
rect 5460 336 5462 338
rect 5490 336 5492 338
rect 5520 336 5522 338
rect 5550 336 5552 338
rect 6268 337 6270 339
rect 6298 337 6300 339
rect 6328 337 6330 339
rect 6358 337 6360 339
rect 6388 337 6390 339
rect 6418 337 6420 339
rect 6448 337 6450 339
rect 6478 337 6480 339
rect 6508 337 6510 339
rect 6538 337 6540 339
rect 6568 337 6570 339
rect 6598 337 6600 339
rect 6628 337 6630 339
rect 6658 337 6660 339
rect 6688 337 6690 339
rect 6718 337 6720 339
rect 6748 337 6750 339
rect 1628 334 1630 336
rect 1600 332 1602 334
rect 1626 332 1628 334
rect 1770 332 1772 334
rect 1768 330 1770 332
rect 4470 330 4472 332
rect 4500 330 4502 332
rect 4530 330 4532 332
rect 4560 330 4562 332
rect 4590 330 4592 332
rect 4620 330 4622 332
rect 4650 330 4652 332
rect 4680 330 4682 332
rect 4710 330 4712 332
rect 4740 330 4742 332
rect 4770 330 4772 332
rect 4800 330 4802 332
rect 4830 330 4832 332
rect 4860 330 4862 332
rect 4890 330 4892 332
rect 4920 330 4922 332
rect 4950 330 4952 332
rect 5070 330 5072 332
rect 5100 330 5102 332
rect 5130 330 5132 332
rect 5160 330 5162 332
rect 5190 330 5192 332
rect 5220 330 5222 332
rect 5250 330 5252 332
rect 5280 330 5282 332
rect 5310 330 5312 332
rect 5340 330 5342 332
rect 5370 330 5372 332
rect 5400 330 5402 332
rect 5430 330 5432 332
rect 5460 330 5462 332
rect 5490 330 5492 332
rect 5520 330 5522 332
rect 5550 330 5552 332
rect 6268 331 6270 333
rect 6298 331 6300 333
rect 6328 331 6330 333
rect 6358 331 6360 333
rect 6388 331 6390 333
rect 6418 331 6420 333
rect 6448 331 6450 333
rect 6478 331 6480 333
rect 6508 331 6510 333
rect 6538 331 6540 333
rect 6568 331 6570 333
rect 6598 331 6600 333
rect 6628 331 6630 333
rect 6658 331 6660 333
rect 6688 331 6690 333
rect 6718 331 6720 333
rect 6748 331 6750 333
rect 4462 328 4464 330
rect 4468 328 4470 330
rect 4492 328 4494 330
rect 4498 328 4500 330
rect 4522 328 4524 330
rect 4528 328 4530 330
rect 4552 328 4554 330
rect 4558 328 4560 330
rect 4582 328 4584 330
rect 4588 328 4590 330
rect 4612 328 4614 330
rect 4618 328 4620 330
rect 4642 328 4644 330
rect 4648 328 4650 330
rect 4672 328 4674 330
rect 4678 328 4680 330
rect 4702 328 4704 330
rect 4708 328 4710 330
rect 4732 328 4734 330
rect 4738 328 4740 330
rect 4762 328 4764 330
rect 4768 328 4770 330
rect 4792 328 4794 330
rect 4798 328 4800 330
rect 4822 328 4824 330
rect 4828 328 4830 330
rect 4852 328 4854 330
rect 4858 328 4860 330
rect 4882 328 4884 330
rect 4888 328 4890 330
rect 4912 328 4914 330
rect 4918 328 4920 330
rect 4942 328 4944 330
rect 4948 328 4950 330
rect 5062 328 5064 330
rect 5068 328 5070 330
rect 5092 328 5094 330
rect 5098 328 5100 330
rect 5122 328 5124 330
rect 5128 328 5130 330
rect 5152 328 5154 330
rect 5158 328 5160 330
rect 5182 328 5184 330
rect 5188 328 5190 330
rect 5212 328 5214 330
rect 5218 328 5220 330
rect 5242 328 5244 330
rect 5248 328 5250 330
rect 5272 328 5274 330
rect 5278 328 5280 330
rect 5302 328 5304 330
rect 5308 328 5310 330
rect 5332 328 5334 330
rect 5338 328 5340 330
rect 5362 328 5364 330
rect 5368 328 5370 330
rect 5392 328 5394 330
rect 5398 328 5400 330
rect 5422 328 5424 330
rect 5428 328 5430 330
rect 5452 328 5454 330
rect 5458 328 5460 330
rect 5482 328 5484 330
rect 5488 328 5490 330
rect 5512 328 5514 330
rect 5518 328 5520 330
rect 5542 328 5544 330
rect 5548 328 5550 330
rect 6260 329 6262 331
rect 6266 329 6268 331
rect 6290 329 6292 331
rect 6296 329 6298 331
rect 6320 329 6322 331
rect 6326 329 6328 331
rect 6350 329 6352 331
rect 6356 329 6358 331
rect 6380 329 6382 331
rect 6386 329 6388 331
rect 6410 329 6412 331
rect 6416 329 6418 331
rect 6440 329 6442 331
rect 6446 329 6448 331
rect 6470 329 6472 331
rect 6476 329 6478 331
rect 6500 329 6502 331
rect 6506 329 6508 331
rect 6530 329 6532 331
rect 6536 329 6538 331
rect 6560 329 6562 331
rect 6566 329 6568 331
rect 6590 329 6592 331
rect 6596 329 6598 331
rect 6620 329 6622 331
rect 6626 329 6628 331
rect 6650 329 6652 331
rect 6656 329 6658 331
rect 6680 329 6682 331
rect 6686 329 6688 331
rect 6710 329 6712 331
rect 6716 329 6718 331
rect 6740 329 6742 331
rect 6746 329 6748 331
rect 4460 326 4462 328
rect 4490 326 4492 328
rect 4520 326 4522 328
rect 4550 326 4552 328
rect 4580 326 4582 328
rect 4610 326 4612 328
rect 4640 326 4642 328
rect 4670 326 4672 328
rect 4700 326 4702 328
rect 4730 326 4732 328
rect 4760 326 4762 328
rect 4790 326 4792 328
rect 4820 326 4822 328
rect 4850 326 4852 328
rect 4880 326 4882 328
rect 4910 326 4912 328
rect 4940 326 4942 328
rect 5060 326 5062 328
rect 5090 326 5092 328
rect 5120 326 5122 328
rect 5150 326 5152 328
rect 5180 326 5182 328
rect 5210 326 5212 328
rect 5240 326 5242 328
rect 5270 326 5272 328
rect 5300 326 5302 328
rect 5330 326 5332 328
rect 5360 326 5362 328
rect 5390 326 5392 328
rect 5420 326 5422 328
rect 5450 326 5452 328
rect 5480 326 5482 328
rect 5510 326 5512 328
rect 5540 326 5542 328
rect 6258 327 6260 329
rect 6288 327 6290 329
rect 6318 327 6320 329
rect 6348 327 6350 329
rect 6378 327 6380 329
rect 6408 327 6410 329
rect 6438 327 6440 329
rect 6468 327 6470 329
rect 6498 327 6500 329
rect 6528 327 6530 329
rect 6558 327 6560 329
rect 6588 327 6590 329
rect 6618 327 6620 329
rect 6648 327 6650 329
rect 6678 327 6680 329
rect 6708 327 6710 329
rect 6738 327 6740 329
rect 1618 324 1620 326
rect 1616 322 1618 324
rect 1760 322 1762 324
rect 1758 320 1760 322
rect 4460 320 4462 322
rect 4490 320 4492 322
rect 4520 320 4522 322
rect 4550 320 4552 322
rect 4580 320 4582 322
rect 4610 320 4612 322
rect 4640 320 4642 322
rect 4670 320 4672 322
rect 4700 320 4702 322
rect 4730 320 4732 322
rect 4760 320 4762 322
rect 4790 320 4792 322
rect 4820 320 4822 322
rect 4850 320 4852 322
rect 4880 320 4882 322
rect 4910 320 4912 322
rect 4940 320 4942 322
rect 5060 320 5062 322
rect 5090 320 5092 322
rect 5120 320 5122 322
rect 5150 320 5152 322
rect 5180 320 5182 322
rect 5210 320 5212 322
rect 5240 320 5242 322
rect 5270 320 5272 322
rect 5300 320 5302 322
rect 5330 320 5332 322
rect 5360 320 5362 322
rect 5390 320 5392 322
rect 5420 320 5422 322
rect 5450 320 5452 322
rect 5480 320 5482 322
rect 5510 320 5512 322
rect 5540 320 5542 322
rect 6258 321 6260 323
rect 6288 321 6290 323
rect 6318 321 6320 323
rect 6348 321 6350 323
rect 6378 321 6380 323
rect 6408 321 6410 323
rect 6438 321 6440 323
rect 6468 321 6470 323
rect 6498 321 6500 323
rect 6528 321 6530 323
rect 6558 321 6560 323
rect 6588 321 6590 323
rect 6618 321 6620 323
rect 6648 321 6650 323
rect 6678 321 6680 323
rect 6708 321 6710 323
rect 6738 321 6740 323
rect 4462 318 4464 320
rect 4468 318 4470 320
rect 4492 318 4494 320
rect 4498 318 4500 320
rect 4522 318 4524 320
rect 4528 318 4530 320
rect 4552 318 4554 320
rect 4558 318 4560 320
rect 4582 318 4584 320
rect 4588 318 4590 320
rect 4612 318 4614 320
rect 4618 318 4620 320
rect 4642 318 4644 320
rect 4648 318 4650 320
rect 4672 318 4674 320
rect 4678 318 4680 320
rect 4702 318 4704 320
rect 4708 318 4710 320
rect 4732 318 4734 320
rect 4738 318 4740 320
rect 4762 318 4764 320
rect 4768 318 4770 320
rect 4792 318 4794 320
rect 4798 318 4800 320
rect 4822 318 4824 320
rect 4828 318 4830 320
rect 4852 318 4854 320
rect 4858 318 4860 320
rect 4882 318 4884 320
rect 4888 318 4890 320
rect 4912 318 4914 320
rect 4918 318 4920 320
rect 4942 318 4944 320
rect 4948 318 4950 320
rect 5062 318 5064 320
rect 5068 318 5070 320
rect 5092 318 5094 320
rect 5098 318 5100 320
rect 5122 318 5124 320
rect 5128 318 5130 320
rect 5152 318 5154 320
rect 5158 318 5160 320
rect 5182 318 5184 320
rect 5188 318 5190 320
rect 5212 318 5214 320
rect 5218 318 5220 320
rect 5242 318 5244 320
rect 5248 318 5250 320
rect 5272 318 5274 320
rect 5278 318 5280 320
rect 5302 318 5304 320
rect 5308 318 5310 320
rect 5332 318 5334 320
rect 5338 318 5340 320
rect 5362 318 5364 320
rect 5368 318 5370 320
rect 5392 318 5394 320
rect 5398 318 5400 320
rect 5422 318 5424 320
rect 5428 318 5430 320
rect 5452 318 5454 320
rect 5458 318 5460 320
rect 5482 318 5484 320
rect 5488 318 5490 320
rect 5512 318 5514 320
rect 5518 318 5520 320
rect 5542 318 5544 320
rect 5548 318 5550 320
rect 6260 319 6262 321
rect 6266 319 6268 321
rect 6290 319 6292 321
rect 6296 319 6298 321
rect 6320 319 6322 321
rect 6326 319 6328 321
rect 6350 319 6352 321
rect 6356 319 6358 321
rect 6380 319 6382 321
rect 6386 319 6388 321
rect 6410 319 6412 321
rect 6416 319 6418 321
rect 6440 319 6442 321
rect 6446 319 6448 321
rect 6470 319 6472 321
rect 6476 319 6478 321
rect 6500 319 6502 321
rect 6506 319 6508 321
rect 6530 319 6532 321
rect 6536 319 6538 321
rect 6560 319 6562 321
rect 6566 319 6568 321
rect 6590 319 6592 321
rect 6596 319 6598 321
rect 6620 319 6622 321
rect 6626 319 6628 321
rect 6650 319 6652 321
rect 6656 319 6658 321
rect 6680 319 6682 321
rect 6686 319 6688 321
rect 6710 319 6712 321
rect 6716 319 6718 321
rect 6740 319 6742 321
rect 6746 319 6748 321
rect 4470 316 4472 318
rect 4500 316 4502 318
rect 4530 316 4532 318
rect 4560 316 4562 318
rect 4590 316 4592 318
rect 4620 316 4622 318
rect 4650 316 4652 318
rect 4680 316 4682 318
rect 4710 316 4712 318
rect 4740 316 4742 318
rect 4770 316 4772 318
rect 4800 316 4802 318
rect 4830 316 4832 318
rect 4860 316 4862 318
rect 4890 316 4892 318
rect 4920 316 4922 318
rect 4950 316 4952 318
rect 5070 316 5072 318
rect 5100 316 5102 318
rect 5130 316 5132 318
rect 5160 316 5162 318
rect 5190 316 5192 318
rect 5220 316 5222 318
rect 5250 316 5252 318
rect 5280 316 5282 318
rect 5310 316 5312 318
rect 5340 316 5342 318
rect 5370 316 5372 318
rect 5400 316 5402 318
rect 5430 316 5432 318
rect 5460 316 5462 318
rect 5490 316 5492 318
rect 5520 316 5522 318
rect 5550 316 5552 318
rect 6268 317 6270 319
rect 6298 317 6300 319
rect 6328 317 6330 319
rect 6358 317 6360 319
rect 6388 317 6390 319
rect 6418 317 6420 319
rect 6448 317 6450 319
rect 6478 317 6480 319
rect 6508 317 6510 319
rect 6538 317 6540 319
rect 6568 317 6570 319
rect 6598 317 6600 319
rect 6628 317 6630 319
rect 6658 317 6660 319
rect 6688 317 6690 319
rect 6718 317 6720 319
rect 6748 317 6750 319
rect 1608 314 1610 316
rect 1606 312 1608 314
rect 1750 312 1752 314
rect 1748 310 1750 312
rect 4470 310 4472 312
rect 4920 310 4922 312
rect 4950 310 4952 312
rect 5070 310 5072 312
rect 5520 310 5522 312
rect 5550 310 5552 312
rect 6268 311 6270 313
rect 6718 311 6720 313
rect 6748 311 6750 313
rect 4462 308 4464 310
rect 4468 308 4470 310
rect 4912 308 4914 310
rect 4918 308 4920 310
rect 4942 308 4944 310
rect 4948 308 4950 310
rect 5062 308 5064 310
rect 5068 308 5070 310
rect 5512 308 5514 310
rect 5518 308 5520 310
rect 5542 308 5544 310
rect 5548 308 5550 310
rect 6260 309 6262 311
rect 6266 309 6268 311
rect 6710 309 6712 311
rect 6716 309 6718 311
rect 6740 309 6742 311
rect 6746 309 6748 311
rect 4460 306 4462 308
rect 4910 306 4912 308
rect 4940 306 4942 308
rect 5060 306 5062 308
rect 5510 306 5512 308
rect 5540 306 5542 308
rect 6258 307 6260 309
rect 6708 307 6710 309
rect 6738 307 6740 309
rect 1740 302 1742 304
rect 1738 300 1740 302
rect 4460 300 4462 302
rect 4910 300 4912 302
rect 4940 300 4942 302
rect 5060 300 5062 302
rect 5510 300 5512 302
rect 5540 300 5542 302
rect 6258 301 6260 303
rect 6708 301 6710 303
rect 6738 301 6740 303
rect 4462 298 4464 300
rect 4468 298 4470 300
rect 4912 298 4914 300
rect 4918 298 4920 300
rect 4942 298 4944 300
rect 4948 298 4950 300
rect 5062 298 5064 300
rect 5068 298 5070 300
rect 5512 298 5514 300
rect 5518 298 5520 300
rect 5542 298 5544 300
rect 5548 298 5550 300
rect 6260 299 6262 301
rect 6266 299 6268 301
rect 6710 299 6712 301
rect 6716 299 6718 301
rect 6740 299 6742 301
rect 6746 299 6748 301
rect 4470 296 4472 298
rect 4920 296 4922 298
rect 4950 296 4952 298
rect 5070 296 5072 298
rect 5520 296 5522 298
rect 5550 296 5552 298
rect 6268 297 6270 299
rect 6718 297 6720 299
rect 6748 297 6750 299
rect 1730 292 1732 294
rect 1728 290 1730 292
rect 3306 290 3308 292
rect 3692 290 3694 292
rect 3906 290 3908 292
rect 4292 290 4294 292
rect 4470 290 4472 292
rect 4500 290 4502 292
rect 4530 290 4532 292
rect 4560 290 4562 292
rect 4590 290 4592 292
rect 4620 290 4622 292
rect 4650 290 4652 292
rect 4680 290 4682 292
rect 4710 290 4712 292
rect 4740 290 4742 292
rect 4770 290 4772 292
rect 4800 290 4802 292
rect 4830 290 4832 292
rect 4860 290 4862 292
rect 4890 290 4892 292
rect 4920 290 4922 292
rect 4950 290 4952 292
rect 5070 290 5072 292
rect 5100 290 5102 292
rect 5130 290 5132 292
rect 5160 290 5162 292
rect 5190 290 5192 292
rect 5220 290 5222 292
rect 5250 290 5252 292
rect 5280 290 5282 292
rect 5310 290 5312 292
rect 5340 290 5342 292
rect 5370 290 5372 292
rect 5400 290 5402 292
rect 5430 290 5432 292
rect 5460 290 5462 292
rect 5490 290 5492 292
rect 5520 290 5522 292
rect 5550 290 5552 292
rect 6268 291 6270 293
rect 6298 291 6300 293
rect 6328 291 6330 293
rect 6358 291 6360 293
rect 6388 291 6390 293
rect 6418 291 6420 293
rect 6448 291 6450 293
rect 6478 291 6480 293
rect 6508 291 6510 293
rect 6538 291 6540 293
rect 6568 291 6570 293
rect 6598 291 6600 293
rect 6628 291 6630 293
rect 6658 291 6660 293
rect 6688 291 6690 293
rect 6718 291 6720 293
rect 6748 291 6750 293
rect 3304 288 3306 290
rect 3694 288 3696 290
rect 3904 288 3906 290
rect 4294 288 4296 290
rect 4462 288 4464 290
rect 4468 288 4470 290
rect 4492 288 4494 290
rect 4498 288 4500 290
rect 4522 288 4524 290
rect 4528 288 4530 290
rect 4552 288 4554 290
rect 4558 288 4560 290
rect 4582 288 4584 290
rect 4588 288 4590 290
rect 4612 288 4614 290
rect 4618 288 4620 290
rect 4642 288 4644 290
rect 4648 288 4650 290
rect 4672 288 4674 290
rect 4678 288 4680 290
rect 4702 288 4704 290
rect 4708 288 4710 290
rect 4732 288 4734 290
rect 4738 288 4740 290
rect 4762 288 4764 290
rect 4768 288 4770 290
rect 4792 288 4794 290
rect 4798 288 4800 290
rect 4822 288 4824 290
rect 4828 288 4830 290
rect 4852 288 4854 290
rect 4858 288 4860 290
rect 4882 288 4884 290
rect 4888 288 4890 290
rect 4912 288 4914 290
rect 4918 288 4920 290
rect 4942 288 4944 290
rect 4948 288 4950 290
rect 5062 288 5064 290
rect 5068 288 5070 290
rect 5092 288 5094 290
rect 5098 288 5100 290
rect 5122 288 5124 290
rect 5128 288 5130 290
rect 5152 288 5154 290
rect 5158 288 5160 290
rect 5182 288 5184 290
rect 5188 288 5190 290
rect 5212 288 5214 290
rect 5218 288 5220 290
rect 5242 288 5244 290
rect 5248 288 5250 290
rect 5272 288 5274 290
rect 5278 288 5280 290
rect 5302 288 5304 290
rect 5308 288 5310 290
rect 5332 288 5334 290
rect 5338 288 5340 290
rect 5362 288 5364 290
rect 5368 288 5370 290
rect 5392 288 5394 290
rect 5398 288 5400 290
rect 5422 288 5424 290
rect 5428 288 5430 290
rect 5452 288 5454 290
rect 5458 288 5460 290
rect 5482 288 5484 290
rect 5488 288 5490 290
rect 5512 288 5514 290
rect 5518 288 5520 290
rect 5542 288 5544 290
rect 5548 288 5550 290
rect 5706 288 5708 290
rect 6092 288 6094 290
rect 6260 289 6262 291
rect 6266 289 6268 291
rect 6290 289 6292 291
rect 6296 289 6298 291
rect 6320 289 6322 291
rect 6326 289 6328 291
rect 6350 289 6352 291
rect 6356 289 6358 291
rect 6380 289 6382 291
rect 6386 289 6388 291
rect 6410 289 6412 291
rect 6416 289 6418 291
rect 6440 289 6442 291
rect 6446 289 6448 291
rect 6470 289 6472 291
rect 6476 289 6478 291
rect 6500 289 6502 291
rect 6506 289 6508 291
rect 6530 289 6532 291
rect 6536 289 6538 291
rect 6560 289 6562 291
rect 6566 289 6568 291
rect 6590 289 6592 291
rect 6596 289 6598 291
rect 6620 289 6622 291
rect 6626 289 6628 291
rect 6650 289 6652 291
rect 6656 289 6658 291
rect 6680 289 6682 291
rect 6686 289 6688 291
rect 6710 289 6712 291
rect 6716 289 6718 291
rect 6740 289 6742 291
rect 6746 289 6748 291
rect 4460 286 4462 288
rect 4490 286 4492 288
rect 4520 286 4522 288
rect 4550 286 4552 288
rect 4580 286 4582 288
rect 4610 286 4612 288
rect 4640 286 4642 288
rect 4670 286 4672 288
rect 4700 286 4702 288
rect 4730 286 4732 288
rect 4760 286 4762 288
rect 4790 286 4792 288
rect 4820 286 4822 288
rect 4850 286 4852 288
rect 4880 286 4882 288
rect 4910 286 4912 288
rect 4940 286 4942 288
rect 5060 286 5062 288
rect 5090 286 5092 288
rect 5120 286 5122 288
rect 5150 286 5152 288
rect 5180 286 5182 288
rect 5210 286 5212 288
rect 5240 286 5242 288
rect 5270 286 5272 288
rect 5300 286 5302 288
rect 5330 286 5332 288
rect 5360 286 5362 288
rect 5390 286 5392 288
rect 5420 286 5422 288
rect 5450 286 5452 288
rect 5480 286 5482 288
rect 5510 286 5512 288
rect 5540 286 5542 288
rect 5704 286 5706 288
rect 6094 286 6096 288
rect 6258 287 6260 289
rect 6288 287 6290 289
rect 6318 287 6320 289
rect 6348 287 6350 289
rect 6378 287 6380 289
rect 6408 287 6410 289
rect 6438 287 6440 289
rect 6468 287 6470 289
rect 6498 287 6500 289
rect 6528 287 6530 289
rect 6558 287 6560 289
rect 6588 287 6590 289
rect 6618 287 6620 289
rect 6648 287 6650 289
rect 6678 287 6680 289
rect 6708 287 6710 289
rect 6738 287 6740 289
rect 1720 282 1722 284
rect 1718 280 1720 282
rect 4460 280 4462 282
rect 4490 280 4492 282
rect 4520 280 4522 282
rect 4550 280 4552 282
rect 4580 280 4582 282
rect 4610 280 4612 282
rect 4640 280 4642 282
rect 4670 280 4672 282
rect 4700 280 4702 282
rect 4730 280 4732 282
rect 4760 280 4762 282
rect 4790 280 4792 282
rect 4820 280 4822 282
rect 4850 280 4852 282
rect 4880 280 4882 282
rect 4910 280 4912 282
rect 4940 280 4942 282
rect 5060 280 5062 282
rect 5090 280 5092 282
rect 5120 280 5122 282
rect 5150 280 5152 282
rect 5180 280 5182 282
rect 5210 280 5212 282
rect 5240 280 5242 282
rect 5270 280 5272 282
rect 5300 280 5302 282
rect 5330 280 5332 282
rect 5360 280 5362 282
rect 5390 280 5392 282
rect 5420 280 5422 282
rect 5450 280 5452 282
rect 5480 280 5482 282
rect 5510 280 5512 282
rect 5540 280 5542 282
rect 6258 281 6260 283
rect 6288 281 6290 283
rect 6318 281 6320 283
rect 6348 281 6350 283
rect 6378 281 6380 283
rect 6408 281 6410 283
rect 6438 281 6440 283
rect 6468 281 6470 283
rect 6498 281 6500 283
rect 6528 281 6530 283
rect 6558 281 6560 283
rect 6588 281 6590 283
rect 6618 281 6620 283
rect 6648 281 6650 283
rect 6678 281 6680 283
rect 6708 281 6710 283
rect 6738 281 6740 283
rect 4462 278 4464 280
rect 4468 278 4470 280
rect 4492 278 4494 280
rect 4498 278 4500 280
rect 4522 278 4524 280
rect 4528 278 4530 280
rect 4552 278 4554 280
rect 4558 278 4560 280
rect 4582 278 4584 280
rect 4588 278 4590 280
rect 4612 278 4614 280
rect 4618 278 4620 280
rect 4642 278 4644 280
rect 4648 278 4650 280
rect 4672 278 4674 280
rect 4678 278 4680 280
rect 4702 278 4704 280
rect 4708 278 4710 280
rect 4732 278 4734 280
rect 4738 278 4740 280
rect 4762 278 4764 280
rect 4768 278 4770 280
rect 4792 278 4794 280
rect 4798 278 4800 280
rect 4822 278 4824 280
rect 4828 278 4830 280
rect 4852 278 4854 280
rect 4858 278 4860 280
rect 4882 278 4884 280
rect 4888 278 4890 280
rect 4912 278 4914 280
rect 4918 278 4920 280
rect 4942 278 4944 280
rect 4948 278 4950 280
rect 5062 278 5064 280
rect 5068 278 5070 280
rect 5092 278 5094 280
rect 5098 278 5100 280
rect 5122 278 5124 280
rect 5128 278 5130 280
rect 5152 278 5154 280
rect 5158 278 5160 280
rect 5182 278 5184 280
rect 5188 278 5190 280
rect 5212 278 5214 280
rect 5218 278 5220 280
rect 5242 278 5244 280
rect 5248 278 5250 280
rect 5272 278 5274 280
rect 5278 278 5280 280
rect 5302 278 5304 280
rect 5308 278 5310 280
rect 5332 278 5334 280
rect 5338 278 5340 280
rect 5362 278 5364 280
rect 5368 278 5370 280
rect 5392 278 5394 280
rect 5398 278 5400 280
rect 5422 278 5424 280
rect 5428 278 5430 280
rect 5452 278 5454 280
rect 5458 278 5460 280
rect 5482 278 5484 280
rect 5488 278 5490 280
rect 5512 278 5514 280
rect 5518 278 5520 280
rect 5542 278 5544 280
rect 5548 278 5550 280
rect 6260 279 6262 281
rect 6266 279 6268 281
rect 6290 279 6292 281
rect 6296 279 6298 281
rect 6320 279 6322 281
rect 6326 279 6328 281
rect 6350 279 6352 281
rect 6356 279 6358 281
rect 6380 279 6382 281
rect 6386 279 6388 281
rect 6410 279 6412 281
rect 6416 279 6418 281
rect 6440 279 6442 281
rect 6446 279 6448 281
rect 6470 279 6472 281
rect 6476 279 6478 281
rect 6500 279 6502 281
rect 6506 279 6508 281
rect 6530 279 6532 281
rect 6536 279 6538 281
rect 6560 279 6562 281
rect 6566 279 6568 281
rect 6590 279 6592 281
rect 6596 279 6598 281
rect 6620 279 6622 281
rect 6626 279 6628 281
rect 6650 279 6652 281
rect 6656 279 6658 281
rect 6680 279 6682 281
rect 6686 279 6688 281
rect 6710 279 6712 281
rect 6716 279 6718 281
rect 6740 279 6742 281
rect 6746 279 6748 281
rect 4470 276 4472 278
rect 4500 276 4502 278
rect 4530 276 4532 278
rect 4560 276 4562 278
rect 4590 276 4592 278
rect 4620 276 4622 278
rect 4650 276 4652 278
rect 4680 276 4682 278
rect 4710 276 4712 278
rect 4740 276 4742 278
rect 4770 276 4772 278
rect 4800 276 4802 278
rect 4830 276 4832 278
rect 4860 276 4862 278
rect 4890 276 4892 278
rect 4920 276 4922 278
rect 4950 276 4952 278
rect 5070 276 5072 278
rect 5100 276 5102 278
rect 5130 276 5132 278
rect 5160 276 5162 278
rect 5190 276 5192 278
rect 5220 276 5222 278
rect 5250 276 5252 278
rect 5280 276 5282 278
rect 5310 276 5312 278
rect 5340 276 5342 278
rect 5370 276 5372 278
rect 5400 276 5402 278
rect 5430 276 5432 278
rect 5460 276 5462 278
rect 5490 276 5492 278
rect 5520 276 5522 278
rect 5550 276 5552 278
rect 6268 277 6270 279
rect 6298 277 6300 279
rect 6328 277 6330 279
rect 6358 277 6360 279
rect 6388 277 6390 279
rect 6418 277 6420 279
rect 6448 277 6450 279
rect 6478 277 6480 279
rect 6508 277 6510 279
rect 6538 277 6540 279
rect 6568 277 6570 279
rect 6598 277 6600 279
rect 6628 277 6630 279
rect 6658 277 6660 279
rect 6688 277 6690 279
rect 6718 277 6720 279
rect 6748 277 6750 279
rect 1710 272 1712 274
rect 1708 270 1710 272
rect 4470 270 4472 272
rect 4500 270 4502 272
rect 4530 270 4532 272
rect 4560 270 4562 272
rect 4590 270 4592 272
rect 4620 270 4622 272
rect 4650 270 4652 272
rect 4680 270 4682 272
rect 4710 270 4712 272
rect 4740 270 4742 272
rect 4770 270 4772 272
rect 4800 270 4802 272
rect 4830 270 4832 272
rect 4860 270 4862 272
rect 4890 270 4892 272
rect 4920 270 4922 272
rect 4950 270 4952 272
rect 5070 270 5072 272
rect 5100 270 5102 272
rect 5130 270 5132 272
rect 5160 270 5162 272
rect 5190 270 5192 272
rect 5220 270 5222 272
rect 5250 270 5252 272
rect 5280 270 5282 272
rect 5310 270 5312 272
rect 5340 270 5342 272
rect 5370 270 5372 272
rect 5400 270 5402 272
rect 5430 270 5432 272
rect 5460 270 5462 272
rect 5490 270 5492 272
rect 5520 270 5522 272
rect 5550 270 5552 272
rect 6268 271 6270 273
rect 6298 271 6300 273
rect 6328 271 6330 273
rect 6358 271 6360 273
rect 6388 271 6390 273
rect 6418 271 6420 273
rect 6448 271 6450 273
rect 6478 271 6480 273
rect 6508 271 6510 273
rect 6538 271 6540 273
rect 6568 271 6570 273
rect 6598 271 6600 273
rect 6628 271 6630 273
rect 6658 271 6660 273
rect 6688 271 6690 273
rect 6718 271 6720 273
rect 6748 271 6750 273
rect 4462 268 4464 270
rect 4468 268 4470 270
rect 4492 268 4494 270
rect 4498 268 4500 270
rect 4522 268 4524 270
rect 4528 268 4530 270
rect 4552 268 4554 270
rect 4558 268 4560 270
rect 4582 268 4584 270
rect 4588 268 4590 270
rect 4612 268 4614 270
rect 4618 268 4620 270
rect 4642 268 4644 270
rect 4648 268 4650 270
rect 4672 268 4674 270
rect 4678 268 4680 270
rect 4702 268 4704 270
rect 4708 268 4710 270
rect 4732 268 4734 270
rect 4738 268 4740 270
rect 4762 268 4764 270
rect 4768 268 4770 270
rect 4792 268 4794 270
rect 4798 268 4800 270
rect 4822 268 4824 270
rect 4828 268 4830 270
rect 4852 268 4854 270
rect 4858 268 4860 270
rect 4882 268 4884 270
rect 4888 268 4890 270
rect 4912 268 4914 270
rect 4918 268 4920 270
rect 4942 268 4944 270
rect 4948 268 4950 270
rect 5062 268 5064 270
rect 5068 268 5070 270
rect 5092 268 5094 270
rect 5098 268 5100 270
rect 5122 268 5124 270
rect 5128 268 5130 270
rect 5152 268 5154 270
rect 5158 268 5160 270
rect 5182 268 5184 270
rect 5188 268 5190 270
rect 5212 268 5214 270
rect 5218 268 5220 270
rect 5242 268 5244 270
rect 5248 268 5250 270
rect 5272 268 5274 270
rect 5278 268 5280 270
rect 5302 268 5304 270
rect 5308 268 5310 270
rect 5332 268 5334 270
rect 5338 268 5340 270
rect 5362 268 5364 270
rect 5368 268 5370 270
rect 5392 268 5394 270
rect 5398 268 5400 270
rect 5422 268 5424 270
rect 5428 268 5430 270
rect 5452 268 5454 270
rect 5458 268 5460 270
rect 5482 268 5484 270
rect 5488 268 5490 270
rect 5512 268 5514 270
rect 5518 268 5520 270
rect 5542 268 5544 270
rect 5548 268 5550 270
rect 6260 269 6262 271
rect 6266 269 6268 271
rect 6290 269 6292 271
rect 6296 269 6298 271
rect 6320 269 6322 271
rect 6326 269 6328 271
rect 6350 269 6352 271
rect 6356 269 6358 271
rect 6380 269 6382 271
rect 6386 269 6388 271
rect 6410 269 6412 271
rect 6416 269 6418 271
rect 6440 269 6442 271
rect 6446 269 6448 271
rect 6470 269 6472 271
rect 6476 269 6478 271
rect 6500 269 6502 271
rect 6506 269 6508 271
rect 6530 269 6532 271
rect 6536 269 6538 271
rect 6560 269 6562 271
rect 6566 269 6568 271
rect 6590 269 6592 271
rect 6596 269 6598 271
rect 6620 269 6622 271
rect 6626 269 6628 271
rect 6650 269 6652 271
rect 6656 269 6658 271
rect 6680 269 6682 271
rect 6686 269 6688 271
rect 6710 269 6712 271
rect 6716 269 6718 271
rect 6740 269 6742 271
rect 6746 269 6748 271
rect 4460 266 4462 268
rect 4490 266 4492 268
rect 4520 266 4522 268
rect 4550 266 4552 268
rect 4580 266 4582 268
rect 4610 266 4612 268
rect 4640 266 4642 268
rect 4670 266 4672 268
rect 4700 266 4702 268
rect 4730 266 4732 268
rect 4760 266 4762 268
rect 4790 266 4792 268
rect 4820 266 4822 268
rect 4850 266 4852 268
rect 4880 266 4882 268
rect 4910 266 4912 268
rect 4940 266 4942 268
rect 5060 266 5062 268
rect 5090 266 5092 268
rect 5120 266 5122 268
rect 5150 266 5152 268
rect 5180 266 5182 268
rect 5210 266 5212 268
rect 5240 266 5242 268
rect 5270 266 5272 268
rect 5300 266 5302 268
rect 5330 266 5332 268
rect 5360 266 5362 268
rect 5390 266 5392 268
rect 5420 266 5422 268
rect 5450 266 5452 268
rect 5480 266 5482 268
rect 5510 266 5512 268
rect 5540 266 5542 268
rect 6258 267 6260 269
rect 6288 267 6290 269
rect 6318 267 6320 269
rect 6348 267 6350 269
rect 6378 267 6380 269
rect 6408 267 6410 269
rect 6438 267 6440 269
rect 6468 267 6470 269
rect 6498 267 6500 269
rect 6528 267 6530 269
rect 6558 267 6560 269
rect 6588 267 6590 269
rect 6618 267 6620 269
rect 6648 267 6650 269
rect 6678 267 6680 269
rect 6708 267 6710 269
rect 6738 267 6740 269
rect 1700 262 1702 264
rect 1698 260 1700 262
rect 4460 260 4462 262
rect 4490 260 4492 262
rect 4520 260 4522 262
rect 4550 260 4552 262
rect 4580 260 4582 262
rect 4610 260 4612 262
rect 4640 260 4642 262
rect 4670 260 4672 262
rect 4700 260 4702 262
rect 4730 260 4732 262
rect 4760 260 4762 262
rect 4790 260 4792 262
rect 4820 260 4822 262
rect 4850 260 4852 262
rect 4880 260 4882 262
rect 4910 260 4912 262
rect 4940 260 4942 262
rect 5060 260 5062 262
rect 5090 260 5092 262
rect 5120 260 5122 262
rect 5150 260 5152 262
rect 5180 260 5182 262
rect 5210 260 5212 262
rect 5240 260 5242 262
rect 5270 260 5272 262
rect 5300 260 5302 262
rect 5330 260 5332 262
rect 5360 260 5362 262
rect 5390 260 5392 262
rect 5420 260 5422 262
rect 5450 260 5452 262
rect 5480 260 5482 262
rect 5510 260 5512 262
rect 5540 260 5542 262
rect 6258 261 6260 263
rect 6288 261 6290 263
rect 6318 261 6320 263
rect 6348 261 6350 263
rect 6378 261 6380 263
rect 6408 261 6410 263
rect 6438 261 6440 263
rect 6468 261 6470 263
rect 6498 261 6500 263
rect 6528 261 6530 263
rect 6558 261 6560 263
rect 6588 261 6590 263
rect 6618 261 6620 263
rect 6648 261 6650 263
rect 6678 261 6680 263
rect 6708 261 6710 263
rect 6738 261 6740 263
rect 4462 258 4464 260
rect 4468 258 4470 260
rect 4492 258 4494 260
rect 4498 258 4500 260
rect 4522 258 4524 260
rect 4528 258 4530 260
rect 4552 258 4554 260
rect 4558 258 4560 260
rect 4582 258 4584 260
rect 4588 258 4590 260
rect 4612 258 4614 260
rect 4618 258 4620 260
rect 4642 258 4644 260
rect 4648 258 4650 260
rect 4672 258 4674 260
rect 4678 258 4680 260
rect 4702 258 4704 260
rect 4708 258 4710 260
rect 4732 258 4734 260
rect 4738 258 4740 260
rect 4762 258 4764 260
rect 4768 258 4770 260
rect 4792 258 4794 260
rect 4798 258 4800 260
rect 4822 258 4824 260
rect 4828 258 4830 260
rect 4852 258 4854 260
rect 4858 258 4860 260
rect 4882 258 4884 260
rect 4888 258 4890 260
rect 4912 258 4914 260
rect 4918 258 4920 260
rect 4942 258 4944 260
rect 4948 258 4950 260
rect 5062 258 5064 260
rect 5068 258 5070 260
rect 5092 258 5094 260
rect 5098 258 5100 260
rect 5122 258 5124 260
rect 5128 258 5130 260
rect 5152 258 5154 260
rect 5158 258 5160 260
rect 5182 258 5184 260
rect 5188 258 5190 260
rect 5212 258 5214 260
rect 5218 258 5220 260
rect 5242 258 5244 260
rect 5248 258 5250 260
rect 5272 258 5274 260
rect 5278 258 5280 260
rect 5302 258 5304 260
rect 5308 258 5310 260
rect 5332 258 5334 260
rect 5338 258 5340 260
rect 5362 258 5364 260
rect 5368 258 5370 260
rect 5392 258 5394 260
rect 5398 258 5400 260
rect 5422 258 5424 260
rect 5428 258 5430 260
rect 5452 258 5454 260
rect 5458 258 5460 260
rect 5482 258 5484 260
rect 5488 258 5490 260
rect 5512 258 5514 260
rect 5518 258 5520 260
rect 5542 258 5544 260
rect 5548 258 5550 260
rect 6260 259 6262 261
rect 6266 259 6268 261
rect 6290 259 6292 261
rect 6296 259 6298 261
rect 6320 259 6322 261
rect 6326 259 6328 261
rect 6350 259 6352 261
rect 6356 259 6358 261
rect 6380 259 6382 261
rect 6386 259 6388 261
rect 6410 259 6412 261
rect 6416 259 6418 261
rect 6440 259 6442 261
rect 6446 259 6448 261
rect 6470 259 6472 261
rect 6476 259 6478 261
rect 6500 259 6502 261
rect 6506 259 6508 261
rect 6530 259 6532 261
rect 6536 259 6538 261
rect 6560 259 6562 261
rect 6566 259 6568 261
rect 6590 259 6592 261
rect 6596 259 6598 261
rect 6620 259 6622 261
rect 6626 259 6628 261
rect 6650 259 6652 261
rect 6656 259 6658 261
rect 6680 259 6682 261
rect 6686 259 6688 261
rect 6710 259 6712 261
rect 6716 259 6718 261
rect 6740 259 6742 261
rect 6746 259 6748 261
rect 4470 256 4472 258
rect 4500 256 4502 258
rect 4530 256 4532 258
rect 4560 256 4562 258
rect 4590 256 4592 258
rect 4620 256 4622 258
rect 4650 256 4652 258
rect 4680 256 4682 258
rect 4710 256 4712 258
rect 4740 256 4742 258
rect 4770 256 4772 258
rect 4800 256 4802 258
rect 4830 256 4832 258
rect 4860 256 4862 258
rect 4890 256 4892 258
rect 4920 256 4922 258
rect 4950 256 4952 258
rect 5070 256 5072 258
rect 5100 256 5102 258
rect 5130 256 5132 258
rect 5160 256 5162 258
rect 5190 256 5192 258
rect 5220 256 5222 258
rect 5250 256 5252 258
rect 5280 256 5282 258
rect 5310 256 5312 258
rect 5340 256 5342 258
rect 5370 256 5372 258
rect 5400 256 5402 258
rect 5430 256 5432 258
rect 5460 256 5462 258
rect 5490 256 5492 258
rect 5520 256 5522 258
rect 5550 256 5552 258
rect 6268 257 6270 259
rect 6298 257 6300 259
rect 6328 257 6330 259
rect 6358 257 6360 259
rect 6388 257 6390 259
rect 6418 257 6420 259
rect 6448 257 6450 259
rect 6478 257 6480 259
rect 6508 257 6510 259
rect 6538 257 6540 259
rect 6568 257 6570 259
rect 6598 257 6600 259
rect 6628 257 6630 259
rect 6658 257 6660 259
rect 6688 257 6690 259
rect 6718 257 6720 259
rect 6748 257 6750 259
rect 1690 252 1692 254
rect 1688 250 1690 252
rect 4470 250 4472 252
rect 4500 250 4502 252
rect 4530 250 4532 252
rect 4560 250 4562 252
rect 4590 250 4592 252
rect 4620 250 4622 252
rect 4650 250 4652 252
rect 4680 250 4682 252
rect 4710 250 4712 252
rect 4740 250 4742 252
rect 4770 250 4772 252
rect 4800 250 4802 252
rect 4830 250 4832 252
rect 4860 250 4862 252
rect 4890 250 4892 252
rect 4920 250 4922 252
rect 4950 250 4952 252
rect 5070 250 5072 252
rect 5100 250 5102 252
rect 5130 250 5132 252
rect 5160 250 5162 252
rect 5190 250 5192 252
rect 5220 250 5222 252
rect 5250 250 5252 252
rect 5280 250 5282 252
rect 5310 250 5312 252
rect 5340 250 5342 252
rect 5370 250 5372 252
rect 5400 250 5402 252
rect 5430 250 5432 252
rect 5460 250 5462 252
rect 5490 250 5492 252
rect 5520 250 5522 252
rect 5550 250 5552 252
rect 6268 251 6270 253
rect 6298 251 6300 253
rect 6328 251 6330 253
rect 6358 251 6360 253
rect 6388 251 6390 253
rect 6418 251 6420 253
rect 6448 251 6450 253
rect 6478 251 6480 253
rect 6508 251 6510 253
rect 6538 251 6540 253
rect 6568 251 6570 253
rect 6598 251 6600 253
rect 6628 251 6630 253
rect 6658 251 6660 253
rect 6688 251 6690 253
rect 6718 251 6720 253
rect 6748 251 6750 253
rect 4462 248 4464 250
rect 4468 248 4470 250
rect 4492 248 4494 250
rect 4498 248 4500 250
rect 4522 248 4524 250
rect 4528 248 4530 250
rect 4552 248 4554 250
rect 4558 248 4560 250
rect 4582 248 4584 250
rect 4588 248 4590 250
rect 4612 248 4614 250
rect 4618 248 4620 250
rect 4642 248 4644 250
rect 4648 248 4650 250
rect 4672 248 4674 250
rect 4678 248 4680 250
rect 4702 248 4704 250
rect 4708 248 4710 250
rect 4732 248 4734 250
rect 4738 248 4740 250
rect 4762 248 4764 250
rect 4768 248 4770 250
rect 4792 248 4794 250
rect 4798 248 4800 250
rect 4822 248 4824 250
rect 4828 248 4830 250
rect 4852 248 4854 250
rect 4858 248 4860 250
rect 4882 248 4884 250
rect 4888 248 4890 250
rect 4912 248 4914 250
rect 4918 248 4920 250
rect 4942 248 4944 250
rect 4948 248 4950 250
rect 5062 248 5064 250
rect 5068 248 5070 250
rect 5092 248 5094 250
rect 5098 248 5100 250
rect 5122 248 5124 250
rect 5128 248 5130 250
rect 5152 248 5154 250
rect 5158 248 5160 250
rect 5182 248 5184 250
rect 5188 248 5190 250
rect 5212 248 5214 250
rect 5218 248 5220 250
rect 5242 248 5244 250
rect 5248 248 5250 250
rect 5272 248 5274 250
rect 5278 248 5280 250
rect 5302 248 5304 250
rect 5308 248 5310 250
rect 5332 248 5334 250
rect 5338 248 5340 250
rect 5362 248 5364 250
rect 5368 248 5370 250
rect 5392 248 5394 250
rect 5398 248 5400 250
rect 5422 248 5424 250
rect 5428 248 5430 250
rect 5452 248 5454 250
rect 5458 248 5460 250
rect 5482 248 5484 250
rect 5488 248 5490 250
rect 5512 248 5514 250
rect 5518 248 5520 250
rect 5542 248 5544 250
rect 5548 248 5550 250
rect 6260 249 6262 251
rect 6266 249 6268 251
rect 6290 249 6292 251
rect 6296 249 6298 251
rect 6320 249 6322 251
rect 6326 249 6328 251
rect 6350 249 6352 251
rect 6356 249 6358 251
rect 6380 249 6382 251
rect 6386 249 6388 251
rect 6410 249 6412 251
rect 6416 249 6418 251
rect 6440 249 6442 251
rect 6446 249 6448 251
rect 6470 249 6472 251
rect 6476 249 6478 251
rect 6500 249 6502 251
rect 6506 249 6508 251
rect 6530 249 6532 251
rect 6536 249 6538 251
rect 6560 249 6562 251
rect 6566 249 6568 251
rect 6590 249 6592 251
rect 6596 249 6598 251
rect 6620 249 6622 251
rect 6626 249 6628 251
rect 6650 249 6652 251
rect 6656 249 6658 251
rect 6680 249 6682 251
rect 6686 249 6688 251
rect 6710 249 6712 251
rect 6716 249 6718 251
rect 6740 249 6742 251
rect 6746 249 6748 251
rect 4460 246 4462 248
rect 4490 246 4492 248
rect 4520 246 4522 248
rect 4550 246 4552 248
rect 4580 246 4582 248
rect 4610 246 4612 248
rect 4640 246 4642 248
rect 4670 246 4672 248
rect 4700 246 4702 248
rect 4730 246 4732 248
rect 4760 246 4762 248
rect 4790 246 4792 248
rect 4820 246 4822 248
rect 4850 246 4852 248
rect 4880 246 4882 248
rect 4910 246 4912 248
rect 4940 246 4942 248
rect 5060 246 5062 248
rect 5090 246 5092 248
rect 5120 246 5122 248
rect 5150 246 5152 248
rect 5180 246 5182 248
rect 5210 246 5212 248
rect 5240 246 5242 248
rect 5270 246 5272 248
rect 5300 246 5302 248
rect 5330 246 5332 248
rect 5360 246 5362 248
rect 5390 246 5392 248
rect 5420 246 5422 248
rect 5450 246 5452 248
rect 5480 246 5482 248
rect 5510 246 5512 248
rect 5540 246 5542 248
rect 6258 247 6260 249
rect 6288 247 6290 249
rect 6318 247 6320 249
rect 6348 247 6350 249
rect 6378 247 6380 249
rect 6408 247 6410 249
rect 6438 247 6440 249
rect 6468 247 6470 249
rect 6498 247 6500 249
rect 6528 247 6530 249
rect 6558 247 6560 249
rect 6588 247 6590 249
rect 6618 247 6620 249
rect 6648 247 6650 249
rect 6678 247 6680 249
rect 6708 247 6710 249
rect 6738 247 6740 249
rect 1680 242 1682 244
rect 1678 240 1680 242
rect 4460 240 4462 242
rect 4490 240 4492 242
rect 4910 240 4912 242
rect 4940 240 4942 242
rect 5060 240 5062 242
rect 5090 240 5092 242
rect 5510 240 5512 242
rect 5540 240 5542 242
rect 6258 241 6260 243
rect 6288 241 6290 243
rect 6708 241 6710 243
rect 6738 241 6740 243
rect 4462 238 4464 240
rect 4488 238 4490 240
rect 4908 238 4910 240
rect 4942 238 4944 240
rect 4948 238 4950 240
rect 5062 238 5064 240
rect 5088 238 5090 240
rect 5508 238 5510 240
rect 5542 238 5544 240
rect 5548 238 5550 240
rect 6260 239 6262 241
rect 6286 239 6288 241
rect 6706 239 6708 241
rect 6740 239 6742 241
rect 6746 239 6748 241
rect 4950 236 4952 238
rect 5550 236 5552 238
rect 6748 237 6750 239
rect 1670 232 1672 234
rect 1668 230 1670 232
rect 4950 230 4952 232
rect 5550 230 5552 232
rect 6748 231 6750 233
rect 3304 228 3306 230
rect 3694 228 3696 230
rect 3904 228 3906 230
rect 4294 228 4296 230
rect 4462 228 4464 230
rect 4488 228 4490 230
rect 4908 228 4910 230
rect 4942 228 4944 230
rect 4948 228 4950 230
rect 5062 228 5064 230
rect 5088 228 5090 230
rect 5508 228 5510 230
rect 5542 228 5544 230
rect 5548 228 5550 230
rect 6260 229 6262 231
rect 6286 229 6288 231
rect 6706 229 6708 231
rect 6740 229 6742 231
rect 6746 229 6748 231
rect 3306 226 3308 228
rect 3692 226 3694 228
rect 3906 226 3908 228
rect 4292 226 4294 228
rect 4460 226 4462 228
rect 4490 226 4492 228
rect 4910 226 4912 228
rect 4940 226 4942 228
rect 5060 226 5062 228
rect 5090 226 5092 228
rect 5510 226 5512 228
rect 5540 226 5542 228
rect 5704 226 5706 228
rect 6094 226 6096 228
rect 6258 227 6260 229
rect 6288 227 6290 229
rect 6708 227 6710 229
rect 6738 227 6740 229
rect 5706 224 5708 226
rect 6092 224 6094 226
rect 1660 222 1662 224
rect 1658 220 1660 222
rect 4460 220 4462 222
rect 4490 220 4492 222
rect 4520 220 4522 222
rect 4550 220 4552 222
rect 4580 220 4582 222
rect 4610 220 4612 222
rect 4640 220 4642 222
rect 4670 220 4672 222
rect 4700 220 4702 222
rect 4730 220 4732 222
rect 4760 220 4762 222
rect 4790 220 4792 222
rect 4820 220 4822 222
rect 4850 220 4852 222
rect 4880 220 4882 222
rect 4910 220 4912 222
rect 4940 220 4942 222
rect 5060 220 5062 222
rect 5090 220 5092 222
rect 5120 220 5122 222
rect 5150 220 5152 222
rect 5180 220 5182 222
rect 5210 220 5212 222
rect 5240 220 5242 222
rect 5270 220 5272 222
rect 5300 220 5302 222
rect 5330 220 5332 222
rect 5360 220 5362 222
rect 5390 220 5392 222
rect 5420 220 5422 222
rect 5450 220 5452 222
rect 5480 220 5482 222
rect 5510 220 5512 222
rect 5540 220 5542 222
rect 6258 221 6260 223
rect 6288 221 6290 223
rect 6318 221 6320 223
rect 6348 221 6350 223
rect 6378 221 6380 223
rect 6408 221 6410 223
rect 6438 221 6440 223
rect 6468 221 6470 223
rect 6498 221 6500 223
rect 6528 221 6530 223
rect 6558 221 6560 223
rect 6588 221 6590 223
rect 6618 221 6620 223
rect 6648 221 6650 223
rect 6678 221 6680 223
rect 6708 221 6710 223
rect 6738 221 6740 223
rect 4462 218 4464 220
rect 4468 218 4470 220
rect 4492 218 4494 220
rect 4498 218 4500 220
rect 4522 218 4524 220
rect 4528 218 4530 220
rect 4552 218 4554 220
rect 4558 218 4560 220
rect 4582 218 4584 220
rect 4588 218 4590 220
rect 4612 218 4614 220
rect 4618 218 4620 220
rect 4642 218 4644 220
rect 4648 218 4650 220
rect 4672 218 4674 220
rect 4678 218 4680 220
rect 4702 218 4704 220
rect 4708 218 4710 220
rect 4732 218 4734 220
rect 4738 218 4740 220
rect 4762 218 4764 220
rect 4768 218 4770 220
rect 4792 218 4794 220
rect 4798 218 4800 220
rect 4822 218 4824 220
rect 4828 218 4830 220
rect 4852 218 4854 220
rect 4858 218 4860 220
rect 4882 218 4884 220
rect 4888 218 4890 220
rect 4912 218 4914 220
rect 4918 218 4920 220
rect 4942 218 4944 220
rect 4948 218 4950 220
rect 5062 218 5064 220
rect 5068 218 5070 220
rect 5092 218 5094 220
rect 5098 218 5100 220
rect 5122 218 5124 220
rect 5128 218 5130 220
rect 5152 218 5154 220
rect 5158 218 5160 220
rect 5182 218 5184 220
rect 5188 218 5190 220
rect 5212 218 5214 220
rect 5218 218 5220 220
rect 5242 218 5244 220
rect 5248 218 5250 220
rect 5272 218 5274 220
rect 5278 218 5280 220
rect 5302 218 5304 220
rect 5308 218 5310 220
rect 5332 218 5334 220
rect 5338 218 5340 220
rect 5362 218 5364 220
rect 5368 218 5370 220
rect 5392 218 5394 220
rect 5398 218 5400 220
rect 5422 218 5424 220
rect 5428 218 5430 220
rect 5452 218 5454 220
rect 5458 218 5460 220
rect 5482 218 5484 220
rect 5488 218 5490 220
rect 5512 218 5514 220
rect 5518 218 5520 220
rect 5542 218 5544 220
rect 5548 218 5550 220
rect 6260 219 6262 221
rect 6266 219 6268 221
rect 6290 219 6292 221
rect 6296 219 6298 221
rect 6320 219 6322 221
rect 6326 219 6328 221
rect 6350 219 6352 221
rect 6356 219 6358 221
rect 6380 219 6382 221
rect 6386 219 6388 221
rect 6410 219 6412 221
rect 6416 219 6418 221
rect 6440 219 6442 221
rect 6446 219 6448 221
rect 6470 219 6472 221
rect 6476 219 6478 221
rect 6500 219 6502 221
rect 6506 219 6508 221
rect 6530 219 6532 221
rect 6536 219 6538 221
rect 6560 219 6562 221
rect 6566 219 6568 221
rect 6590 219 6592 221
rect 6596 219 6598 221
rect 6620 219 6622 221
rect 6626 219 6628 221
rect 6650 219 6652 221
rect 6656 219 6658 221
rect 6680 219 6682 221
rect 6686 219 6688 221
rect 6710 219 6712 221
rect 6716 219 6718 221
rect 6740 219 6742 221
rect 6746 219 6748 221
rect 4470 216 4472 218
rect 4500 216 4502 218
rect 4530 216 4532 218
rect 4560 216 4562 218
rect 4590 216 4592 218
rect 4620 216 4622 218
rect 4650 216 4652 218
rect 4680 216 4682 218
rect 4710 216 4712 218
rect 4740 216 4742 218
rect 4770 216 4772 218
rect 4800 216 4802 218
rect 4830 216 4832 218
rect 4860 216 4862 218
rect 4890 216 4892 218
rect 4920 216 4922 218
rect 4950 216 4952 218
rect 5070 216 5072 218
rect 5100 216 5102 218
rect 5130 216 5132 218
rect 5160 216 5162 218
rect 5190 216 5192 218
rect 5220 216 5222 218
rect 5250 216 5252 218
rect 5280 216 5282 218
rect 5310 216 5312 218
rect 5340 216 5342 218
rect 5370 216 5372 218
rect 5400 216 5402 218
rect 5430 216 5432 218
rect 5460 216 5462 218
rect 5490 216 5492 218
rect 5520 216 5522 218
rect 5550 216 5552 218
rect 6268 217 6270 219
rect 6298 217 6300 219
rect 6328 217 6330 219
rect 6358 217 6360 219
rect 6388 217 6390 219
rect 6418 217 6420 219
rect 6448 217 6450 219
rect 6478 217 6480 219
rect 6508 217 6510 219
rect 6538 217 6540 219
rect 6568 217 6570 219
rect 6598 217 6600 219
rect 6628 217 6630 219
rect 6658 217 6660 219
rect 6688 217 6690 219
rect 6718 217 6720 219
rect 6748 217 6750 219
rect 1650 212 1652 214
rect 1648 210 1650 212
rect 4470 210 4472 212
rect 4500 210 4502 212
rect 4530 210 4532 212
rect 4560 210 4562 212
rect 4590 210 4592 212
rect 4620 210 4622 212
rect 4650 210 4652 212
rect 4680 210 4682 212
rect 4710 210 4712 212
rect 4740 210 4742 212
rect 4770 210 4772 212
rect 4800 210 4802 212
rect 4830 210 4832 212
rect 4860 210 4862 212
rect 4890 210 4892 212
rect 4920 210 4922 212
rect 4950 210 4952 212
rect 5070 210 5072 212
rect 5100 210 5102 212
rect 5130 210 5132 212
rect 5160 210 5162 212
rect 5190 210 5192 212
rect 5220 210 5222 212
rect 5250 210 5252 212
rect 5280 210 5282 212
rect 5310 210 5312 212
rect 5340 210 5342 212
rect 5370 210 5372 212
rect 5400 210 5402 212
rect 5430 210 5432 212
rect 5460 210 5462 212
rect 5490 210 5492 212
rect 5520 210 5522 212
rect 5550 210 5552 212
rect 6268 211 6270 213
rect 6298 211 6300 213
rect 6328 211 6330 213
rect 6358 211 6360 213
rect 6388 211 6390 213
rect 6418 211 6420 213
rect 6448 211 6450 213
rect 6478 211 6480 213
rect 6508 211 6510 213
rect 6538 211 6540 213
rect 6568 211 6570 213
rect 6598 211 6600 213
rect 6628 211 6630 213
rect 6658 211 6660 213
rect 6688 211 6690 213
rect 6718 211 6720 213
rect 6748 211 6750 213
rect 4462 208 4464 210
rect 4468 208 4470 210
rect 4492 208 4494 210
rect 4498 208 4500 210
rect 4522 208 4524 210
rect 4528 208 4530 210
rect 4552 208 4554 210
rect 4558 208 4560 210
rect 4582 208 4584 210
rect 4588 208 4590 210
rect 4612 208 4614 210
rect 4618 208 4620 210
rect 4642 208 4644 210
rect 4648 208 4650 210
rect 4672 208 4674 210
rect 4678 208 4680 210
rect 4702 208 4704 210
rect 4708 208 4710 210
rect 4732 208 4734 210
rect 4738 208 4740 210
rect 4762 208 4764 210
rect 4768 208 4770 210
rect 4792 208 4794 210
rect 4798 208 4800 210
rect 4822 208 4824 210
rect 4828 208 4830 210
rect 4852 208 4854 210
rect 4858 208 4860 210
rect 4882 208 4884 210
rect 4888 208 4890 210
rect 4912 208 4914 210
rect 4918 208 4920 210
rect 4942 208 4944 210
rect 4948 208 4950 210
rect 5062 208 5064 210
rect 5068 208 5070 210
rect 5092 208 5094 210
rect 5098 208 5100 210
rect 5122 208 5124 210
rect 5128 208 5130 210
rect 5152 208 5154 210
rect 5158 208 5160 210
rect 5182 208 5184 210
rect 5188 208 5190 210
rect 5212 208 5214 210
rect 5218 208 5220 210
rect 5242 208 5244 210
rect 5248 208 5250 210
rect 5272 208 5274 210
rect 5278 208 5280 210
rect 5302 208 5304 210
rect 5308 208 5310 210
rect 5332 208 5334 210
rect 5338 208 5340 210
rect 5362 208 5364 210
rect 5368 208 5370 210
rect 5392 208 5394 210
rect 5398 208 5400 210
rect 5422 208 5424 210
rect 5428 208 5430 210
rect 5452 208 5454 210
rect 5458 208 5460 210
rect 5482 208 5484 210
rect 5488 208 5490 210
rect 5512 208 5514 210
rect 5518 208 5520 210
rect 5542 208 5544 210
rect 5548 208 5550 210
rect 6260 209 6262 211
rect 6266 209 6268 211
rect 6290 209 6292 211
rect 6296 209 6298 211
rect 6320 209 6322 211
rect 6326 209 6328 211
rect 6350 209 6352 211
rect 6356 209 6358 211
rect 6380 209 6382 211
rect 6386 209 6388 211
rect 6410 209 6412 211
rect 6416 209 6418 211
rect 6440 209 6442 211
rect 6446 209 6448 211
rect 6470 209 6472 211
rect 6476 209 6478 211
rect 6500 209 6502 211
rect 6506 209 6508 211
rect 6530 209 6532 211
rect 6536 209 6538 211
rect 6560 209 6562 211
rect 6566 209 6568 211
rect 6590 209 6592 211
rect 6596 209 6598 211
rect 6620 209 6622 211
rect 6626 209 6628 211
rect 6650 209 6652 211
rect 6656 209 6658 211
rect 6680 209 6682 211
rect 6686 209 6688 211
rect 6710 209 6712 211
rect 6716 209 6718 211
rect 6740 209 6742 211
rect 6746 209 6748 211
rect 4460 206 4462 208
rect 4490 206 4492 208
rect 4520 206 4522 208
rect 4550 206 4552 208
rect 4580 206 4582 208
rect 4610 206 4612 208
rect 4640 206 4642 208
rect 4670 206 4672 208
rect 4700 206 4702 208
rect 4730 206 4732 208
rect 4760 206 4762 208
rect 4790 206 4792 208
rect 4820 206 4822 208
rect 4850 206 4852 208
rect 4880 206 4882 208
rect 4910 206 4912 208
rect 4940 206 4942 208
rect 5060 206 5062 208
rect 5090 206 5092 208
rect 5120 206 5122 208
rect 5150 206 5152 208
rect 5180 206 5182 208
rect 5210 206 5212 208
rect 5240 206 5242 208
rect 5270 206 5272 208
rect 5300 206 5302 208
rect 5330 206 5332 208
rect 5360 206 5362 208
rect 5390 206 5392 208
rect 5420 206 5422 208
rect 5450 206 5452 208
rect 5480 206 5482 208
rect 5510 206 5512 208
rect 5540 206 5542 208
rect 6258 207 6260 209
rect 6288 207 6290 209
rect 6318 207 6320 209
rect 6348 207 6350 209
rect 6378 207 6380 209
rect 6408 207 6410 209
rect 6438 207 6440 209
rect 6468 207 6470 209
rect 6498 207 6500 209
rect 6528 207 6530 209
rect 6558 207 6560 209
rect 6588 207 6590 209
rect 6618 207 6620 209
rect 6648 207 6650 209
rect 6678 207 6680 209
rect 6708 207 6710 209
rect 6738 207 6740 209
rect 1640 202 1642 204
rect 1638 200 1640 202
rect 4460 200 4462 202
rect 4490 200 4492 202
rect 4520 200 4522 202
rect 4550 200 4552 202
rect 4580 200 4582 202
rect 4610 200 4612 202
rect 4640 200 4642 202
rect 4670 200 4672 202
rect 4700 200 4702 202
rect 4730 200 4732 202
rect 4760 200 4762 202
rect 4790 200 4792 202
rect 4820 200 4822 202
rect 4850 200 4852 202
rect 4880 200 4882 202
rect 4910 200 4912 202
rect 4940 200 4942 202
rect 5060 200 5062 202
rect 5090 200 5092 202
rect 5120 200 5122 202
rect 5150 200 5152 202
rect 5180 200 5182 202
rect 5210 200 5212 202
rect 5240 200 5242 202
rect 5270 200 5272 202
rect 5300 200 5302 202
rect 5330 200 5332 202
rect 5360 200 5362 202
rect 5390 200 5392 202
rect 5420 200 5422 202
rect 5450 200 5452 202
rect 5480 200 5482 202
rect 5510 200 5512 202
rect 5540 200 5542 202
rect 6258 201 6260 203
rect 6288 201 6290 203
rect 6318 201 6320 203
rect 6348 201 6350 203
rect 6378 201 6380 203
rect 6408 201 6410 203
rect 6438 201 6440 203
rect 6468 201 6470 203
rect 6498 201 6500 203
rect 6528 201 6530 203
rect 6558 201 6560 203
rect 6588 201 6590 203
rect 6618 201 6620 203
rect 6648 201 6650 203
rect 6678 201 6680 203
rect 6708 201 6710 203
rect 6738 201 6740 203
rect 4462 198 4464 200
rect 4468 198 4470 200
rect 4492 198 4494 200
rect 4498 198 4500 200
rect 4522 198 4524 200
rect 4528 198 4530 200
rect 4552 198 4554 200
rect 4558 198 4560 200
rect 4582 198 4584 200
rect 4588 198 4590 200
rect 4612 198 4614 200
rect 4618 198 4620 200
rect 4642 198 4644 200
rect 4648 198 4650 200
rect 4672 198 4674 200
rect 4678 198 4680 200
rect 4702 198 4704 200
rect 4708 198 4710 200
rect 4732 198 4734 200
rect 4738 198 4740 200
rect 4762 198 4764 200
rect 4768 198 4770 200
rect 4792 198 4794 200
rect 4798 198 4800 200
rect 4822 198 4824 200
rect 4828 198 4830 200
rect 4852 198 4854 200
rect 4858 198 4860 200
rect 4882 198 4884 200
rect 4888 198 4890 200
rect 4912 198 4914 200
rect 4918 198 4920 200
rect 4942 198 4944 200
rect 4948 198 4950 200
rect 5062 198 5064 200
rect 5068 198 5070 200
rect 5092 198 5094 200
rect 5098 198 5100 200
rect 5122 198 5124 200
rect 5128 198 5130 200
rect 5152 198 5154 200
rect 5158 198 5160 200
rect 5182 198 5184 200
rect 5188 198 5190 200
rect 5212 198 5214 200
rect 5218 198 5220 200
rect 5242 198 5244 200
rect 5248 198 5250 200
rect 5272 198 5274 200
rect 5278 198 5280 200
rect 5302 198 5304 200
rect 5308 198 5310 200
rect 5332 198 5334 200
rect 5338 198 5340 200
rect 5362 198 5364 200
rect 5368 198 5370 200
rect 5392 198 5394 200
rect 5398 198 5400 200
rect 5422 198 5424 200
rect 5428 198 5430 200
rect 5452 198 5454 200
rect 5458 198 5460 200
rect 5482 198 5484 200
rect 5488 198 5490 200
rect 5512 198 5514 200
rect 5518 198 5520 200
rect 5542 198 5544 200
rect 5548 198 5550 200
rect 6260 199 6262 201
rect 6266 199 6268 201
rect 6290 199 6292 201
rect 6296 199 6298 201
rect 6320 199 6322 201
rect 6326 199 6328 201
rect 6350 199 6352 201
rect 6356 199 6358 201
rect 6380 199 6382 201
rect 6386 199 6388 201
rect 6410 199 6412 201
rect 6416 199 6418 201
rect 6440 199 6442 201
rect 6446 199 6448 201
rect 6470 199 6472 201
rect 6476 199 6478 201
rect 6500 199 6502 201
rect 6506 199 6508 201
rect 6530 199 6532 201
rect 6536 199 6538 201
rect 6560 199 6562 201
rect 6566 199 6568 201
rect 6590 199 6592 201
rect 6596 199 6598 201
rect 6620 199 6622 201
rect 6626 199 6628 201
rect 6650 199 6652 201
rect 6656 199 6658 201
rect 6680 199 6682 201
rect 6686 199 6688 201
rect 6710 199 6712 201
rect 6716 199 6718 201
rect 6740 199 6742 201
rect 6746 199 6748 201
rect 4470 196 4472 198
rect 4500 196 4502 198
rect 4530 196 4532 198
rect 4560 196 4562 198
rect 4590 196 4592 198
rect 4620 196 4622 198
rect 4650 196 4652 198
rect 4680 196 4682 198
rect 4710 196 4712 198
rect 4740 196 4742 198
rect 4770 196 4772 198
rect 4800 196 4802 198
rect 4830 196 4832 198
rect 4860 196 4862 198
rect 4890 196 4892 198
rect 4920 196 4922 198
rect 4950 196 4952 198
rect 5070 196 5072 198
rect 5100 196 5102 198
rect 5130 196 5132 198
rect 5160 196 5162 198
rect 5190 196 5192 198
rect 5220 196 5222 198
rect 5250 196 5252 198
rect 5280 196 5282 198
rect 5310 196 5312 198
rect 5340 196 5342 198
rect 5370 196 5372 198
rect 5400 196 5402 198
rect 5430 196 5432 198
rect 5460 196 5462 198
rect 5490 196 5492 198
rect 5520 196 5522 198
rect 5550 196 5552 198
rect 6268 197 6270 199
rect 6298 197 6300 199
rect 6328 197 6330 199
rect 6358 197 6360 199
rect 6388 197 6390 199
rect 6418 197 6420 199
rect 6448 197 6450 199
rect 6478 197 6480 199
rect 6508 197 6510 199
rect 6538 197 6540 199
rect 6568 197 6570 199
rect 6598 197 6600 199
rect 6628 197 6630 199
rect 6658 197 6660 199
rect 6688 197 6690 199
rect 6718 197 6720 199
rect 6748 197 6750 199
rect 1630 192 1632 194
rect 1628 190 1630 192
rect 4470 190 4472 192
rect 4500 190 4502 192
rect 4530 190 4532 192
rect 4560 190 4562 192
rect 4590 190 4592 192
rect 4620 190 4622 192
rect 4650 190 4652 192
rect 4680 190 4682 192
rect 4710 190 4712 192
rect 4740 190 4742 192
rect 4770 190 4772 192
rect 4800 190 4802 192
rect 4830 190 4832 192
rect 4860 190 4862 192
rect 4890 190 4892 192
rect 4920 190 4922 192
rect 4950 190 4952 192
rect 5070 190 5072 192
rect 5100 190 5102 192
rect 5130 190 5132 192
rect 5160 190 5162 192
rect 5190 190 5192 192
rect 5220 190 5222 192
rect 5250 190 5252 192
rect 5280 190 5282 192
rect 5310 190 5312 192
rect 5340 190 5342 192
rect 5370 190 5372 192
rect 5400 190 5402 192
rect 5430 190 5432 192
rect 5460 190 5462 192
rect 5490 190 5492 192
rect 5520 190 5522 192
rect 5550 190 5552 192
rect 6268 191 6270 193
rect 6298 191 6300 193
rect 6328 191 6330 193
rect 6358 191 6360 193
rect 6388 191 6390 193
rect 6418 191 6420 193
rect 6448 191 6450 193
rect 6478 191 6480 193
rect 6508 191 6510 193
rect 6538 191 6540 193
rect 6568 191 6570 193
rect 6598 191 6600 193
rect 6628 191 6630 193
rect 6658 191 6660 193
rect 6688 191 6690 193
rect 6718 191 6720 193
rect 6748 191 6750 193
rect 4462 188 4464 190
rect 4468 188 4470 190
rect 4492 188 4494 190
rect 4498 188 4500 190
rect 4522 188 4524 190
rect 4528 188 4530 190
rect 4552 188 4554 190
rect 4558 188 4560 190
rect 4582 188 4584 190
rect 4588 188 4590 190
rect 4612 188 4614 190
rect 4618 188 4620 190
rect 4642 188 4644 190
rect 4648 188 4650 190
rect 4672 188 4674 190
rect 4678 188 4680 190
rect 4702 188 4704 190
rect 4708 188 4710 190
rect 4732 188 4734 190
rect 4738 188 4740 190
rect 4762 188 4764 190
rect 4768 188 4770 190
rect 4792 188 4794 190
rect 4798 188 4800 190
rect 4822 188 4824 190
rect 4828 188 4830 190
rect 4852 188 4854 190
rect 4858 188 4860 190
rect 4882 188 4884 190
rect 4888 188 4890 190
rect 4912 188 4914 190
rect 4918 188 4920 190
rect 4942 188 4944 190
rect 4948 188 4950 190
rect 5062 188 5064 190
rect 5068 188 5070 190
rect 5092 188 5094 190
rect 5098 188 5100 190
rect 5122 188 5124 190
rect 5128 188 5130 190
rect 5152 188 5154 190
rect 5158 188 5160 190
rect 5182 188 5184 190
rect 5188 188 5190 190
rect 5212 188 5214 190
rect 5218 188 5220 190
rect 5242 188 5244 190
rect 5248 188 5250 190
rect 5272 188 5274 190
rect 5278 188 5280 190
rect 5302 188 5304 190
rect 5308 188 5310 190
rect 5332 188 5334 190
rect 5338 188 5340 190
rect 5362 188 5364 190
rect 5368 188 5370 190
rect 5392 188 5394 190
rect 5398 188 5400 190
rect 5422 188 5424 190
rect 5428 188 5430 190
rect 5452 188 5454 190
rect 5458 188 5460 190
rect 5482 188 5484 190
rect 5488 188 5490 190
rect 5512 188 5514 190
rect 5518 188 5520 190
rect 5542 188 5544 190
rect 5548 188 5550 190
rect 6260 189 6262 191
rect 6266 189 6268 191
rect 6290 189 6292 191
rect 6296 189 6298 191
rect 6320 189 6322 191
rect 6326 189 6328 191
rect 6350 189 6352 191
rect 6356 189 6358 191
rect 6380 189 6382 191
rect 6386 189 6388 191
rect 6410 189 6412 191
rect 6416 189 6418 191
rect 6440 189 6442 191
rect 6446 189 6448 191
rect 6470 189 6472 191
rect 6476 189 6478 191
rect 6500 189 6502 191
rect 6506 189 6508 191
rect 6530 189 6532 191
rect 6536 189 6538 191
rect 6560 189 6562 191
rect 6566 189 6568 191
rect 6590 189 6592 191
rect 6596 189 6598 191
rect 6620 189 6622 191
rect 6626 189 6628 191
rect 6650 189 6652 191
rect 6656 189 6658 191
rect 6680 189 6682 191
rect 6686 189 6688 191
rect 6710 189 6712 191
rect 6716 189 6718 191
rect 6740 189 6742 191
rect 6746 189 6748 191
rect 4460 186 4462 188
rect 4490 186 4492 188
rect 4520 186 4522 188
rect 4550 186 4552 188
rect 4580 186 4582 188
rect 4610 186 4612 188
rect 4640 186 4642 188
rect 4670 186 4672 188
rect 4700 186 4702 188
rect 4730 186 4732 188
rect 4760 186 4762 188
rect 4790 186 4792 188
rect 4820 186 4822 188
rect 4850 186 4852 188
rect 4880 186 4882 188
rect 4910 186 4912 188
rect 4940 186 4942 188
rect 5060 186 5062 188
rect 5090 186 5092 188
rect 5120 186 5122 188
rect 5150 186 5152 188
rect 5180 186 5182 188
rect 5210 186 5212 188
rect 5240 186 5242 188
rect 5270 186 5272 188
rect 5300 186 5302 188
rect 5330 186 5332 188
rect 5360 186 5362 188
rect 5390 186 5392 188
rect 5420 186 5422 188
rect 5450 186 5452 188
rect 5480 186 5482 188
rect 5510 186 5512 188
rect 5540 186 5542 188
rect 6258 187 6260 189
rect 6288 187 6290 189
rect 6318 187 6320 189
rect 6348 187 6350 189
rect 6378 187 6380 189
rect 6408 187 6410 189
rect 6438 187 6440 189
rect 6468 187 6470 189
rect 6498 187 6500 189
rect 6528 187 6530 189
rect 6558 187 6560 189
rect 6588 187 6590 189
rect 6618 187 6620 189
rect 6648 187 6650 189
rect 6678 187 6680 189
rect 6708 187 6710 189
rect 6738 187 6740 189
rect 1620 182 1622 184
rect 1618 180 1620 182
rect 4460 180 4462 182
rect 4490 180 4492 182
rect 4520 180 4522 182
rect 4550 180 4552 182
rect 4580 180 4582 182
rect 4610 180 4612 182
rect 4640 180 4642 182
rect 4670 180 4672 182
rect 4700 180 4702 182
rect 4730 180 4732 182
rect 4760 180 4762 182
rect 4790 180 4792 182
rect 4820 180 4822 182
rect 4850 180 4852 182
rect 4880 180 4882 182
rect 4910 180 4912 182
rect 4940 180 4942 182
rect 5060 180 5062 182
rect 5090 180 5092 182
rect 5120 180 5122 182
rect 5150 180 5152 182
rect 5180 180 5182 182
rect 5210 180 5212 182
rect 5240 180 5242 182
rect 5270 180 5272 182
rect 5300 180 5302 182
rect 5330 180 5332 182
rect 5360 180 5362 182
rect 5390 180 5392 182
rect 5420 180 5422 182
rect 5450 180 5452 182
rect 5480 180 5482 182
rect 5510 180 5512 182
rect 5540 180 5542 182
rect 6258 181 6260 183
rect 6288 181 6290 183
rect 6318 181 6320 183
rect 6348 181 6350 183
rect 6378 181 6380 183
rect 6408 181 6410 183
rect 6438 181 6440 183
rect 6468 181 6470 183
rect 6498 181 6500 183
rect 6528 181 6530 183
rect 6558 181 6560 183
rect 6588 181 6590 183
rect 6618 181 6620 183
rect 6648 181 6650 183
rect 6678 181 6680 183
rect 6708 181 6710 183
rect 6738 181 6740 183
rect 4462 178 4464 180
rect 4468 178 4470 180
rect 4492 178 4494 180
rect 4498 178 4500 180
rect 4522 178 4524 180
rect 4528 178 4530 180
rect 4552 178 4554 180
rect 4558 178 4560 180
rect 4582 178 4584 180
rect 4588 178 4590 180
rect 4612 178 4614 180
rect 4618 178 4620 180
rect 4642 178 4644 180
rect 4648 178 4650 180
rect 4672 178 4674 180
rect 4678 178 4680 180
rect 4702 178 4704 180
rect 4708 178 4710 180
rect 4732 178 4734 180
rect 4738 178 4740 180
rect 4762 178 4764 180
rect 4768 178 4770 180
rect 4792 178 4794 180
rect 4798 178 4800 180
rect 4822 178 4824 180
rect 4828 178 4830 180
rect 4852 178 4854 180
rect 4858 178 4860 180
rect 4882 178 4884 180
rect 4888 178 4890 180
rect 4912 178 4914 180
rect 4918 178 4920 180
rect 4942 178 4944 180
rect 4948 178 4950 180
rect 5062 178 5064 180
rect 5068 178 5070 180
rect 5092 178 5094 180
rect 5098 178 5100 180
rect 5122 178 5124 180
rect 5128 178 5130 180
rect 5152 178 5154 180
rect 5158 178 5160 180
rect 5182 178 5184 180
rect 5188 178 5190 180
rect 5212 178 5214 180
rect 5218 178 5220 180
rect 5242 178 5244 180
rect 5248 178 5250 180
rect 5272 178 5274 180
rect 5278 178 5280 180
rect 5302 178 5304 180
rect 5308 178 5310 180
rect 5332 178 5334 180
rect 5338 178 5340 180
rect 5362 178 5364 180
rect 5368 178 5370 180
rect 5392 178 5394 180
rect 5398 178 5400 180
rect 5422 178 5424 180
rect 5428 178 5430 180
rect 5452 178 5454 180
rect 5458 178 5460 180
rect 5482 178 5484 180
rect 5488 178 5490 180
rect 5512 178 5514 180
rect 5518 178 5520 180
rect 5542 178 5544 180
rect 5548 178 5550 180
rect 6260 179 6262 181
rect 6266 179 6268 181
rect 6290 179 6292 181
rect 6296 179 6298 181
rect 6320 179 6322 181
rect 6326 179 6328 181
rect 6350 179 6352 181
rect 6356 179 6358 181
rect 6380 179 6382 181
rect 6386 179 6388 181
rect 6410 179 6412 181
rect 6416 179 6418 181
rect 6440 179 6442 181
rect 6446 179 6448 181
rect 6470 179 6472 181
rect 6476 179 6478 181
rect 6500 179 6502 181
rect 6506 179 6508 181
rect 6530 179 6532 181
rect 6536 179 6538 181
rect 6560 179 6562 181
rect 6566 179 6568 181
rect 6590 179 6592 181
rect 6596 179 6598 181
rect 6620 179 6622 181
rect 6626 179 6628 181
rect 6650 179 6652 181
rect 6656 179 6658 181
rect 6680 179 6682 181
rect 6686 179 6688 181
rect 6710 179 6712 181
rect 6716 179 6718 181
rect 6740 179 6742 181
rect 6746 179 6748 181
rect 4470 176 4472 178
rect 4500 176 4502 178
rect 4530 176 4532 178
rect 4560 176 4562 178
rect 4590 176 4592 178
rect 4620 176 4622 178
rect 4650 176 4652 178
rect 4680 176 4682 178
rect 4710 176 4712 178
rect 4740 176 4742 178
rect 4770 176 4772 178
rect 4800 176 4802 178
rect 4830 176 4832 178
rect 4860 176 4862 178
rect 4890 176 4892 178
rect 4920 176 4922 178
rect 4950 176 4952 178
rect 5070 176 5072 178
rect 5100 176 5102 178
rect 5130 176 5132 178
rect 5160 176 5162 178
rect 5190 176 5192 178
rect 5220 176 5222 178
rect 5250 176 5252 178
rect 5280 176 5282 178
rect 5310 176 5312 178
rect 5340 176 5342 178
rect 5370 176 5372 178
rect 5400 176 5402 178
rect 5430 176 5432 178
rect 5460 176 5462 178
rect 5490 176 5492 178
rect 5520 176 5522 178
rect 5550 176 5552 178
rect 6268 177 6270 179
rect 6298 177 6300 179
rect 6328 177 6330 179
rect 6358 177 6360 179
rect 6388 177 6390 179
rect 6418 177 6420 179
rect 6448 177 6450 179
rect 6478 177 6480 179
rect 6508 177 6510 179
rect 6538 177 6540 179
rect 6568 177 6570 179
rect 6598 177 6600 179
rect 6628 177 6630 179
rect 6658 177 6660 179
rect 6688 177 6690 179
rect 6718 177 6720 179
rect 6748 177 6750 179
rect 1610 172 1612 174
rect 1608 170 1610 172
rect 4470 170 4472 172
rect 4500 170 4502 172
rect 4530 170 4532 172
rect 4560 170 4562 172
rect 4590 170 4592 172
rect 4620 170 4622 172
rect 4650 170 4652 172
rect 4680 170 4682 172
rect 4710 170 4712 172
rect 4740 170 4742 172
rect 4770 170 4772 172
rect 4800 170 4802 172
rect 4830 170 4832 172
rect 4860 170 4862 172
rect 4890 170 4892 172
rect 4920 170 4922 172
rect 4950 170 4952 172
rect 5070 170 5072 172
rect 5100 170 5102 172
rect 5130 170 5132 172
rect 5160 170 5162 172
rect 5190 170 5192 172
rect 5220 170 5222 172
rect 5250 170 5252 172
rect 5280 170 5282 172
rect 5310 170 5312 172
rect 5340 170 5342 172
rect 5370 170 5372 172
rect 5400 170 5402 172
rect 5430 170 5432 172
rect 5460 170 5462 172
rect 5490 170 5492 172
rect 5520 170 5522 172
rect 5550 170 5552 172
rect 6268 171 6270 173
rect 6298 171 6300 173
rect 6328 171 6330 173
rect 6358 171 6360 173
rect 6388 171 6390 173
rect 6418 171 6420 173
rect 6448 171 6450 173
rect 6478 171 6480 173
rect 6508 171 6510 173
rect 6538 171 6540 173
rect 6568 171 6570 173
rect 6598 171 6600 173
rect 6628 171 6630 173
rect 6658 171 6660 173
rect 6688 171 6690 173
rect 6718 171 6720 173
rect 6748 171 6750 173
rect 4462 168 4464 170
rect 4468 168 4470 170
rect 4492 168 4494 170
rect 4498 168 4500 170
rect 4522 168 4524 170
rect 4528 168 4530 170
rect 4552 168 4554 170
rect 4558 168 4560 170
rect 4582 168 4584 170
rect 4588 168 4590 170
rect 4612 168 4614 170
rect 4618 168 4620 170
rect 4642 168 4644 170
rect 4648 168 4650 170
rect 4672 168 4674 170
rect 4678 168 4680 170
rect 4702 168 4704 170
rect 4708 168 4710 170
rect 4732 168 4734 170
rect 4738 168 4740 170
rect 4762 168 4764 170
rect 4768 168 4770 170
rect 4792 168 4794 170
rect 4798 168 4800 170
rect 4822 168 4824 170
rect 4828 168 4830 170
rect 4852 168 4854 170
rect 4858 168 4860 170
rect 4882 168 4884 170
rect 4888 168 4890 170
rect 4912 168 4914 170
rect 4918 168 4920 170
rect 4942 168 4944 170
rect 4948 168 4950 170
rect 5062 168 5064 170
rect 5068 168 5070 170
rect 5092 168 5094 170
rect 5098 168 5100 170
rect 5122 168 5124 170
rect 5128 168 5130 170
rect 5152 168 5154 170
rect 5158 168 5160 170
rect 5182 168 5184 170
rect 5188 168 5190 170
rect 5212 168 5214 170
rect 5218 168 5220 170
rect 5242 168 5244 170
rect 5248 168 5250 170
rect 5272 168 5274 170
rect 5278 168 5280 170
rect 5302 168 5304 170
rect 5308 168 5310 170
rect 5332 168 5334 170
rect 5338 168 5340 170
rect 5362 168 5364 170
rect 5368 168 5370 170
rect 5392 168 5394 170
rect 5398 168 5400 170
rect 5422 168 5424 170
rect 5428 168 5430 170
rect 5452 168 5454 170
rect 5458 168 5460 170
rect 5482 168 5484 170
rect 5488 168 5490 170
rect 5512 168 5514 170
rect 5518 168 5520 170
rect 5542 168 5544 170
rect 5548 168 5550 170
rect 6260 169 6262 171
rect 6266 169 6268 171
rect 6290 169 6292 171
rect 6296 169 6298 171
rect 6320 169 6322 171
rect 6326 169 6328 171
rect 6350 169 6352 171
rect 6356 169 6358 171
rect 6380 169 6382 171
rect 6386 169 6388 171
rect 6410 169 6412 171
rect 6416 169 6418 171
rect 6440 169 6442 171
rect 6446 169 6448 171
rect 6470 169 6472 171
rect 6476 169 6478 171
rect 6500 169 6502 171
rect 6506 169 6508 171
rect 6530 169 6532 171
rect 6536 169 6538 171
rect 6560 169 6562 171
rect 6566 169 6568 171
rect 6590 169 6592 171
rect 6596 169 6598 171
rect 6620 169 6622 171
rect 6626 169 6628 171
rect 6650 169 6652 171
rect 6656 169 6658 171
rect 6680 169 6682 171
rect 6686 169 6688 171
rect 6710 169 6712 171
rect 6716 169 6718 171
rect 6740 169 6742 171
rect 6746 169 6748 171
rect 4460 166 4462 168
rect 4490 166 4492 168
rect 4520 166 4522 168
rect 4550 166 4552 168
rect 4580 166 4582 168
rect 4610 166 4612 168
rect 4640 166 4642 168
rect 4670 166 4672 168
rect 4700 166 4702 168
rect 4730 166 4732 168
rect 4760 166 4762 168
rect 4790 166 4792 168
rect 4820 166 4822 168
rect 4850 166 4852 168
rect 4880 166 4882 168
rect 4910 166 4912 168
rect 4940 166 4942 168
rect 5060 166 5062 168
rect 5090 166 5092 168
rect 5120 166 5122 168
rect 5150 166 5152 168
rect 5180 166 5182 168
rect 5210 166 5212 168
rect 5240 166 5242 168
rect 5270 166 5272 168
rect 5300 166 5302 168
rect 5330 166 5332 168
rect 5360 166 5362 168
rect 5390 166 5392 168
rect 5420 166 5422 168
rect 5450 166 5452 168
rect 5480 166 5482 168
rect 5510 166 5512 168
rect 5540 166 5542 168
rect 6258 167 6260 169
rect 6288 167 6290 169
rect 6318 167 6320 169
rect 6348 167 6350 169
rect 6378 167 6380 169
rect 6408 167 6410 169
rect 6438 167 6440 169
rect 6468 167 6470 169
rect 6498 167 6500 169
rect 6528 167 6530 169
rect 6558 167 6560 169
rect 6588 167 6590 169
rect 6618 167 6620 169
rect 6648 167 6650 169
rect 6678 167 6680 169
rect 6708 167 6710 169
rect 6738 167 6740 169
rect 1600 162 1602 164
rect 3306 160 3308 162
rect 3692 160 3694 162
rect 3906 160 3908 162
rect 4292 160 4294 162
rect 4460 160 4462 162
rect 4490 160 4492 162
rect 4910 160 4912 162
rect 4940 160 4942 162
rect 5060 160 5062 162
rect 5090 160 5092 162
rect 5510 160 5512 162
rect 5540 160 5542 162
rect 6258 161 6260 163
rect 6288 161 6290 163
rect 6708 161 6710 163
rect 6738 161 6740 163
rect 3304 158 3306 160
rect 3694 158 3696 160
rect 3904 158 3906 160
rect 4294 158 4296 160
rect 4462 158 4464 160
rect 4468 158 4470 160
rect 4492 158 4494 160
rect 4908 158 4910 160
rect 4942 158 4944 160
rect 4948 158 4950 160
rect 5062 158 5064 160
rect 5068 158 5070 160
rect 5092 158 5094 160
rect 5508 158 5510 160
rect 5542 158 5544 160
rect 5548 158 5550 160
rect 5706 158 5708 160
rect 6092 158 6094 160
rect 6260 159 6262 161
rect 6266 159 6268 161
rect 6290 159 6292 161
rect 6706 159 6708 161
rect 6740 159 6742 161
rect 6746 159 6748 161
rect 4470 156 4472 158
rect 4950 156 4952 158
rect 5070 156 5072 158
rect 5550 156 5552 158
rect 5704 156 5706 158
rect 6094 156 6096 158
rect 6268 157 6270 159
rect 6748 157 6750 159
rect 4470 150 4472 152
rect 4950 150 4952 152
rect 5070 150 5072 152
rect 5550 150 5552 152
rect 6268 151 6270 153
rect 6748 151 6750 153
rect 4462 148 4464 150
rect 4468 148 4470 150
rect 4492 148 4494 150
rect 4908 148 4910 150
rect 4942 148 4944 150
rect 4948 148 4950 150
rect 5062 148 5064 150
rect 5068 148 5070 150
rect 5092 148 5094 150
rect 5508 148 5510 150
rect 5542 148 5544 150
rect 5548 148 5550 150
rect 6260 149 6262 151
rect 6266 149 6268 151
rect 6290 149 6292 151
rect 6706 149 6708 151
rect 6740 149 6742 151
rect 6746 149 6748 151
rect 4460 146 4462 148
rect 4490 146 4492 148
rect 4910 146 4912 148
rect 4940 146 4942 148
rect 5060 146 5062 148
rect 5090 146 5092 148
rect 5510 146 5512 148
rect 5540 146 5542 148
rect 6258 147 6260 149
rect 6288 147 6290 149
rect 6708 147 6710 149
rect 6738 147 6740 149
rect 4460 140 4462 142
rect 4490 140 4492 142
rect 4520 140 4522 142
rect 4550 140 4552 142
rect 4580 140 4582 142
rect 4610 140 4612 142
rect 4640 140 4642 142
rect 4670 140 4672 142
rect 4700 140 4702 142
rect 4730 140 4732 142
rect 4760 140 4762 142
rect 4790 140 4792 142
rect 4820 140 4822 142
rect 4850 140 4852 142
rect 4880 140 4882 142
rect 4910 140 4912 142
rect 4940 140 4942 142
rect 5060 140 5062 142
rect 5090 140 5092 142
rect 5120 140 5122 142
rect 5150 140 5152 142
rect 5180 140 5182 142
rect 5210 140 5212 142
rect 5240 140 5242 142
rect 5270 140 5272 142
rect 5300 140 5302 142
rect 5330 140 5332 142
rect 5360 140 5362 142
rect 5390 140 5392 142
rect 5420 140 5422 142
rect 5450 140 5452 142
rect 5480 140 5482 142
rect 5510 140 5512 142
rect 5540 140 5542 142
rect 6258 141 6260 143
rect 6288 141 6290 143
rect 6318 141 6320 143
rect 6348 141 6350 143
rect 6378 141 6380 143
rect 6408 141 6410 143
rect 6438 141 6440 143
rect 6468 141 6470 143
rect 6498 141 6500 143
rect 6528 141 6530 143
rect 6558 141 6560 143
rect 6588 141 6590 143
rect 6618 141 6620 143
rect 6648 141 6650 143
rect 6678 141 6680 143
rect 6708 141 6710 143
rect 6738 141 6740 143
rect 4462 138 4464 140
rect 4468 138 4470 140
rect 4492 138 4494 140
rect 4498 138 4500 140
rect 4522 138 4524 140
rect 4528 138 4530 140
rect 4552 138 4554 140
rect 4558 138 4560 140
rect 4582 138 4584 140
rect 4588 138 4590 140
rect 4612 138 4614 140
rect 4618 138 4620 140
rect 4642 138 4644 140
rect 4648 138 4650 140
rect 4672 138 4674 140
rect 4678 138 4680 140
rect 4702 138 4704 140
rect 4708 138 4710 140
rect 4732 138 4734 140
rect 4738 138 4740 140
rect 4762 138 4764 140
rect 4768 138 4770 140
rect 4792 138 4794 140
rect 4798 138 4800 140
rect 4822 138 4824 140
rect 4828 138 4830 140
rect 4852 138 4854 140
rect 4858 138 4860 140
rect 4882 138 4884 140
rect 4888 138 4890 140
rect 4912 138 4914 140
rect 4918 138 4920 140
rect 4942 138 4944 140
rect 4948 138 4950 140
rect 5062 138 5064 140
rect 5068 138 5070 140
rect 5092 138 5094 140
rect 5098 138 5100 140
rect 5122 138 5124 140
rect 5128 138 5130 140
rect 5152 138 5154 140
rect 5158 138 5160 140
rect 5182 138 5184 140
rect 5188 138 5190 140
rect 5212 138 5214 140
rect 5218 138 5220 140
rect 5242 138 5244 140
rect 5248 138 5250 140
rect 5272 138 5274 140
rect 5278 138 5280 140
rect 5302 138 5304 140
rect 5308 138 5310 140
rect 5332 138 5334 140
rect 5338 138 5340 140
rect 5362 138 5364 140
rect 5368 138 5370 140
rect 5392 138 5394 140
rect 5398 138 5400 140
rect 5422 138 5424 140
rect 5428 138 5430 140
rect 5452 138 5454 140
rect 5458 138 5460 140
rect 5482 138 5484 140
rect 5488 138 5490 140
rect 5512 138 5514 140
rect 5518 138 5520 140
rect 5542 138 5544 140
rect 5548 138 5550 140
rect 6260 139 6262 141
rect 6266 139 6268 141
rect 6290 139 6292 141
rect 6296 139 6298 141
rect 6320 139 6322 141
rect 6326 139 6328 141
rect 6350 139 6352 141
rect 6356 139 6358 141
rect 6380 139 6382 141
rect 6386 139 6388 141
rect 6410 139 6412 141
rect 6416 139 6418 141
rect 6440 139 6442 141
rect 6446 139 6448 141
rect 6470 139 6472 141
rect 6476 139 6478 141
rect 6500 139 6502 141
rect 6506 139 6508 141
rect 6530 139 6532 141
rect 6536 139 6538 141
rect 6560 139 6562 141
rect 6566 139 6568 141
rect 6590 139 6592 141
rect 6596 139 6598 141
rect 6620 139 6622 141
rect 6626 139 6628 141
rect 6650 139 6652 141
rect 6656 139 6658 141
rect 6680 139 6682 141
rect 6686 139 6688 141
rect 6710 139 6712 141
rect 6716 139 6718 141
rect 6740 139 6742 141
rect 6746 139 6748 141
rect 4470 136 4472 138
rect 4500 136 4502 138
rect 4530 136 4532 138
rect 4560 136 4562 138
rect 4590 136 4592 138
rect 4620 136 4622 138
rect 4650 136 4652 138
rect 4680 136 4682 138
rect 4710 136 4712 138
rect 4740 136 4742 138
rect 4770 136 4772 138
rect 4800 136 4802 138
rect 4830 136 4832 138
rect 4860 136 4862 138
rect 4890 136 4892 138
rect 4920 136 4922 138
rect 4950 136 4952 138
rect 5070 136 5072 138
rect 5100 136 5102 138
rect 5130 136 5132 138
rect 5160 136 5162 138
rect 5190 136 5192 138
rect 5220 136 5222 138
rect 5250 136 5252 138
rect 5280 136 5282 138
rect 5310 136 5312 138
rect 5340 136 5342 138
rect 5370 136 5372 138
rect 5400 136 5402 138
rect 5430 136 5432 138
rect 5460 136 5462 138
rect 5490 136 5492 138
rect 5520 136 5522 138
rect 5550 136 5552 138
rect 6268 137 6270 139
rect 6298 137 6300 139
rect 6328 137 6330 139
rect 6358 137 6360 139
rect 6388 137 6390 139
rect 6418 137 6420 139
rect 6448 137 6450 139
rect 6478 137 6480 139
rect 6508 137 6510 139
rect 6538 137 6540 139
rect 6568 137 6570 139
rect 6598 137 6600 139
rect 6628 137 6630 139
rect 6658 137 6660 139
rect 6688 137 6690 139
rect 6718 137 6720 139
rect 6748 137 6750 139
rect 4470 130 4472 132
rect 4500 130 4502 132
rect 4530 130 4532 132
rect 4560 130 4562 132
rect 4590 130 4592 132
rect 4620 130 4622 132
rect 4650 130 4652 132
rect 4680 130 4682 132
rect 4710 130 4712 132
rect 4740 130 4742 132
rect 4770 130 4772 132
rect 4800 130 4802 132
rect 4830 130 4832 132
rect 4860 130 4862 132
rect 4890 130 4892 132
rect 4920 130 4922 132
rect 4950 130 4952 132
rect 5070 130 5072 132
rect 5100 130 5102 132
rect 5130 130 5132 132
rect 5160 130 5162 132
rect 5190 130 5192 132
rect 5220 130 5222 132
rect 5250 130 5252 132
rect 5280 130 5282 132
rect 5310 130 5312 132
rect 5340 130 5342 132
rect 5370 130 5372 132
rect 5400 130 5402 132
rect 5430 130 5432 132
rect 5460 130 5462 132
rect 5490 130 5492 132
rect 5520 130 5522 132
rect 5550 130 5552 132
rect 6268 131 6270 133
rect 6298 131 6300 133
rect 6328 131 6330 133
rect 6358 131 6360 133
rect 6388 131 6390 133
rect 6418 131 6420 133
rect 6448 131 6450 133
rect 6478 131 6480 133
rect 6508 131 6510 133
rect 6538 131 6540 133
rect 6568 131 6570 133
rect 6598 131 6600 133
rect 6628 131 6630 133
rect 6658 131 6660 133
rect 6688 131 6690 133
rect 6718 131 6720 133
rect 6748 131 6750 133
rect 4462 128 4464 130
rect 4468 128 4470 130
rect 4492 128 4494 130
rect 4498 128 4500 130
rect 4522 128 4524 130
rect 4528 128 4530 130
rect 4552 128 4554 130
rect 4558 128 4560 130
rect 4582 128 4584 130
rect 4588 128 4590 130
rect 4612 128 4614 130
rect 4618 128 4620 130
rect 4642 128 4644 130
rect 4648 128 4650 130
rect 4672 128 4674 130
rect 4678 128 4680 130
rect 4702 128 4704 130
rect 4708 128 4710 130
rect 4732 128 4734 130
rect 4738 128 4740 130
rect 4762 128 4764 130
rect 4768 128 4770 130
rect 4792 128 4794 130
rect 4798 128 4800 130
rect 4822 128 4824 130
rect 4828 128 4830 130
rect 4852 128 4854 130
rect 4858 128 4860 130
rect 4882 128 4884 130
rect 4888 128 4890 130
rect 4912 128 4914 130
rect 4918 128 4920 130
rect 4942 128 4944 130
rect 4948 128 4950 130
rect 5062 128 5064 130
rect 5068 128 5070 130
rect 5092 128 5094 130
rect 5098 128 5100 130
rect 5122 128 5124 130
rect 5128 128 5130 130
rect 5152 128 5154 130
rect 5158 128 5160 130
rect 5182 128 5184 130
rect 5188 128 5190 130
rect 5212 128 5214 130
rect 5218 128 5220 130
rect 5242 128 5244 130
rect 5248 128 5250 130
rect 5272 128 5274 130
rect 5278 128 5280 130
rect 5302 128 5304 130
rect 5308 128 5310 130
rect 5332 128 5334 130
rect 5338 128 5340 130
rect 5362 128 5364 130
rect 5368 128 5370 130
rect 5392 128 5394 130
rect 5398 128 5400 130
rect 5422 128 5424 130
rect 5428 128 5430 130
rect 5452 128 5454 130
rect 5458 128 5460 130
rect 5482 128 5484 130
rect 5488 128 5490 130
rect 5512 128 5514 130
rect 5518 128 5520 130
rect 5542 128 5544 130
rect 5548 128 5550 130
rect 6260 129 6262 131
rect 6266 129 6268 131
rect 6290 129 6292 131
rect 6296 129 6298 131
rect 6320 129 6322 131
rect 6326 129 6328 131
rect 6350 129 6352 131
rect 6356 129 6358 131
rect 6380 129 6382 131
rect 6386 129 6388 131
rect 6410 129 6412 131
rect 6416 129 6418 131
rect 6440 129 6442 131
rect 6446 129 6448 131
rect 6470 129 6472 131
rect 6476 129 6478 131
rect 6500 129 6502 131
rect 6506 129 6508 131
rect 6530 129 6532 131
rect 6536 129 6538 131
rect 6560 129 6562 131
rect 6566 129 6568 131
rect 6590 129 6592 131
rect 6596 129 6598 131
rect 6620 129 6622 131
rect 6626 129 6628 131
rect 6650 129 6652 131
rect 6656 129 6658 131
rect 6680 129 6682 131
rect 6686 129 6688 131
rect 6710 129 6712 131
rect 6716 129 6718 131
rect 6740 129 6742 131
rect 6746 129 6748 131
rect 4460 126 4462 128
rect 4490 126 4492 128
rect 4520 126 4522 128
rect 4550 126 4552 128
rect 4580 126 4582 128
rect 4610 126 4612 128
rect 4640 126 4642 128
rect 4670 126 4672 128
rect 4700 126 4702 128
rect 4730 126 4732 128
rect 4760 126 4762 128
rect 4790 126 4792 128
rect 4820 126 4822 128
rect 4850 126 4852 128
rect 4880 126 4882 128
rect 4910 126 4912 128
rect 4940 126 4942 128
rect 5060 126 5062 128
rect 5090 126 5092 128
rect 5120 126 5122 128
rect 5150 126 5152 128
rect 5180 126 5182 128
rect 5210 126 5212 128
rect 5240 126 5242 128
rect 5270 126 5272 128
rect 5300 126 5302 128
rect 5330 126 5332 128
rect 5360 126 5362 128
rect 5390 126 5392 128
rect 5420 126 5422 128
rect 5450 126 5452 128
rect 5480 126 5482 128
rect 5510 126 5512 128
rect 5540 126 5542 128
rect 6258 127 6260 129
rect 6288 127 6290 129
rect 6318 127 6320 129
rect 6348 127 6350 129
rect 6378 127 6380 129
rect 6408 127 6410 129
rect 6438 127 6440 129
rect 6468 127 6470 129
rect 6498 127 6500 129
rect 6528 127 6530 129
rect 6558 127 6560 129
rect 6588 127 6590 129
rect 6618 127 6620 129
rect 6648 127 6650 129
rect 6678 127 6680 129
rect 6708 127 6710 129
rect 6738 127 6740 129
rect 4460 120 4462 122
rect 4490 120 4492 122
rect 4520 120 4522 122
rect 4550 120 4552 122
rect 4580 120 4582 122
rect 4610 120 4612 122
rect 4640 120 4642 122
rect 4670 120 4672 122
rect 4700 120 4702 122
rect 4730 120 4732 122
rect 4760 120 4762 122
rect 4790 120 4792 122
rect 4820 120 4822 122
rect 4850 120 4852 122
rect 4880 120 4882 122
rect 4910 120 4912 122
rect 4940 120 4942 122
rect 5060 120 5062 122
rect 5090 120 5092 122
rect 5120 120 5122 122
rect 5150 120 5152 122
rect 5180 120 5182 122
rect 5210 120 5212 122
rect 5240 120 5242 122
rect 5270 120 5272 122
rect 5300 120 5302 122
rect 5330 120 5332 122
rect 5360 120 5362 122
rect 5390 120 5392 122
rect 5420 120 5422 122
rect 5450 120 5452 122
rect 5480 120 5482 122
rect 5510 120 5512 122
rect 5540 120 5542 122
rect 6258 121 6260 123
rect 6288 121 6290 123
rect 6318 121 6320 123
rect 6348 121 6350 123
rect 6378 121 6380 123
rect 6408 121 6410 123
rect 6438 121 6440 123
rect 6468 121 6470 123
rect 6498 121 6500 123
rect 6528 121 6530 123
rect 6558 121 6560 123
rect 6588 121 6590 123
rect 6618 121 6620 123
rect 6648 121 6650 123
rect 6678 121 6680 123
rect 6708 121 6710 123
rect 6738 121 6740 123
rect 4462 118 4464 120
rect 4468 118 4470 120
rect 4492 118 4494 120
rect 4498 118 4500 120
rect 4522 118 4524 120
rect 4528 118 4530 120
rect 4552 118 4554 120
rect 4558 118 4560 120
rect 4582 118 4584 120
rect 4588 118 4590 120
rect 4612 118 4614 120
rect 4618 118 4620 120
rect 4642 118 4644 120
rect 4648 118 4650 120
rect 4672 118 4674 120
rect 4678 118 4680 120
rect 4702 118 4704 120
rect 4708 118 4710 120
rect 4732 118 4734 120
rect 4738 118 4740 120
rect 4762 118 4764 120
rect 4768 118 4770 120
rect 4792 118 4794 120
rect 4798 118 4800 120
rect 4822 118 4824 120
rect 4828 118 4830 120
rect 4852 118 4854 120
rect 4858 118 4860 120
rect 4882 118 4884 120
rect 4888 118 4890 120
rect 4912 118 4914 120
rect 4918 118 4920 120
rect 4942 118 4944 120
rect 4948 118 4950 120
rect 5062 118 5064 120
rect 5068 118 5070 120
rect 5092 118 5094 120
rect 5098 118 5100 120
rect 5122 118 5124 120
rect 5128 118 5130 120
rect 5152 118 5154 120
rect 5158 118 5160 120
rect 5182 118 5184 120
rect 5188 118 5190 120
rect 5212 118 5214 120
rect 5218 118 5220 120
rect 5242 118 5244 120
rect 5248 118 5250 120
rect 5272 118 5274 120
rect 5278 118 5280 120
rect 5302 118 5304 120
rect 5308 118 5310 120
rect 5332 118 5334 120
rect 5338 118 5340 120
rect 5362 118 5364 120
rect 5368 118 5370 120
rect 5392 118 5394 120
rect 5398 118 5400 120
rect 5422 118 5424 120
rect 5428 118 5430 120
rect 5452 118 5454 120
rect 5458 118 5460 120
rect 5482 118 5484 120
rect 5488 118 5490 120
rect 5512 118 5514 120
rect 5518 118 5520 120
rect 5542 118 5544 120
rect 5548 118 5550 120
rect 6260 119 6262 121
rect 6266 119 6268 121
rect 6290 119 6292 121
rect 6296 119 6298 121
rect 6320 119 6322 121
rect 6326 119 6328 121
rect 6350 119 6352 121
rect 6356 119 6358 121
rect 6380 119 6382 121
rect 6386 119 6388 121
rect 6410 119 6412 121
rect 6416 119 6418 121
rect 6440 119 6442 121
rect 6446 119 6448 121
rect 6470 119 6472 121
rect 6476 119 6478 121
rect 6500 119 6502 121
rect 6506 119 6508 121
rect 6530 119 6532 121
rect 6536 119 6538 121
rect 6560 119 6562 121
rect 6566 119 6568 121
rect 6590 119 6592 121
rect 6596 119 6598 121
rect 6620 119 6622 121
rect 6626 119 6628 121
rect 6650 119 6652 121
rect 6656 119 6658 121
rect 6680 119 6682 121
rect 6686 119 6688 121
rect 6710 119 6712 121
rect 6716 119 6718 121
rect 6740 119 6742 121
rect 6746 119 6748 121
rect 4470 116 4472 118
rect 4500 116 4502 118
rect 4530 116 4532 118
rect 4560 116 4562 118
rect 4590 116 4592 118
rect 4620 116 4622 118
rect 4650 116 4652 118
rect 4680 116 4682 118
rect 4710 116 4712 118
rect 4740 116 4742 118
rect 4770 116 4772 118
rect 4800 116 4802 118
rect 4830 116 4832 118
rect 4860 116 4862 118
rect 4890 116 4892 118
rect 4920 116 4922 118
rect 4950 116 4952 118
rect 5070 116 5072 118
rect 5100 116 5102 118
rect 5130 116 5132 118
rect 5160 116 5162 118
rect 5190 116 5192 118
rect 5220 116 5222 118
rect 5250 116 5252 118
rect 5280 116 5282 118
rect 5310 116 5312 118
rect 5340 116 5342 118
rect 5370 116 5372 118
rect 5400 116 5402 118
rect 5430 116 5432 118
rect 5460 116 5462 118
rect 5490 116 5492 118
rect 5520 116 5522 118
rect 5550 116 5552 118
rect 6268 117 6270 119
rect 6298 117 6300 119
rect 6328 117 6330 119
rect 6358 117 6360 119
rect 6388 117 6390 119
rect 6418 117 6420 119
rect 6448 117 6450 119
rect 6478 117 6480 119
rect 6508 117 6510 119
rect 6538 117 6540 119
rect 6568 117 6570 119
rect 6598 117 6600 119
rect 6628 117 6630 119
rect 6658 117 6660 119
rect 6688 117 6690 119
rect 6718 117 6720 119
rect 6748 117 6750 119
rect 4470 110 4472 112
rect 4500 110 4502 112
rect 4530 110 4532 112
rect 4560 110 4562 112
rect 4590 110 4592 112
rect 4620 110 4622 112
rect 4650 110 4652 112
rect 4680 110 4682 112
rect 4710 110 4712 112
rect 4740 110 4742 112
rect 4770 110 4772 112
rect 4800 110 4802 112
rect 4830 110 4832 112
rect 4860 110 4862 112
rect 4890 110 4892 112
rect 4920 110 4922 112
rect 4950 110 4952 112
rect 5070 110 5072 112
rect 5100 110 5102 112
rect 5130 110 5132 112
rect 5160 110 5162 112
rect 5190 110 5192 112
rect 5220 110 5222 112
rect 5250 110 5252 112
rect 5280 110 5282 112
rect 5310 110 5312 112
rect 5340 110 5342 112
rect 5370 110 5372 112
rect 5400 110 5402 112
rect 5430 110 5432 112
rect 5460 110 5462 112
rect 5490 110 5492 112
rect 5520 110 5522 112
rect 5550 110 5552 112
rect 6268 111 6270 113
rect 6298 111 6300 113
rect 6328 111 6330 113
rect 6358 111 6360 113
rect 6388 111 6390 113
rect 6418 111 6420 113
rect 6448 111 6450 113
rect 6478 111 6480 113
rect 6508 111 6510 113
rect 6538 111 6540 113
rect 6568 111 6570 113
rect 6598 111 6600 113
rect 6628 111 6630 113
rect 6658 111 6660 113
rect 6688 111 6690 113
rect 6718 111 6720 113
rect 6748 111 6750 113
rect 4462 108 4464 110
rect 4468 108 4470 110
rect 4492 108 4494 110
rect 4498 108 4500 110
rect 4522 108 4524 110
rect 4528 108 4530 110
rect 4552 108 4554 110
rect 4558 108 4560 110
rect 4582 108 4584 110
rect 4588 108 4590 110
rect 4612 108 4614 110
rect 4618 108 4620 110
rect 4642 108 4644 110
rect 4648 108 4650 110
rect 4672 108 4674 110
rect 4678 108 4680 110
rect 4702 108 4704 110
rect 4708 108 4710 110
rect 4732 108 4734 110
rect 4738 108 4740 110
rect 4762 108 4764 110
rect 4768 108 4770 110
rect 4792 108 4794 110
rect 4798 108 4800 110
rect 4822 108 4824 110
rect 4828 108 4830 110
rect 4852 108 4854 110
rect 4858 108 4860 110
rect 4882 108 4884 110
rect 4888 108 4890 110
rect 4912 108 4914 110
rect 4918 108 4920 110
rect 4942 108 4944 110
rect 4948 108 4950 110
rect 5062 108 5064 110
rect 5068 108 5070 110
rect 5092 108 5094 110
rect 5098 108 5100 110
rect 5122 108 5124 110
rect 5128 108 5130 110
rect 5152 108 5154 110
rect 5158 108 5160 110
rect 5182 108 5184 110
rect 5188 108 5190 110
rect 5212 108 5214 110
rect 5218 108 5220 110
rect 5242 108 5244 110
rect 5248 108 5250 110
rect 5272 108 5274 110
rect 5278 108 5280 110
rect 5302 108 5304 110
rect 5308 108 5310 110
rect 5332 108 5334 110
rect 5338 108 5340 110
rect 5362 108 5364 110
rect 5368 108 5370 110
rect 5392 108 5394 110
rect 5398 108 5400 110
rect 5422 108 5424 110
rect 5428 108 5430 110
rect 5452 108 5454 110
rect 5458 108 5460 110
rect 5482 108 5484 110
rect 5488 108 5490 110
rect 5512 108 5514 110
rect 5518 108 5520 110
rect 5542 108 5544 110
rect 5548 108 5550 110
rect 6260 109 6262 111
rect 6266 109 6268 111
rect 6290 109 6292 111
rect 6296 109 6298 111
rect 6320 109 6322 111
rect 6326 109 6328 111
rect 6350 109 6352 111
rect 6356 109 6358 111
rect 6380 109 6382 111
rect 6386 109 6388 111
rect 6410 109 6412 111
rect 6416 109 6418 111
rect 6440 109 6442 111
rect 6446 109 6448 111
rect 6470 109 6472 111
rect 6476 109 6478 111
rect 6500 109 6502 111
rect 6506 109 6508 111
rect 6530 109 6532 111
rect 6536 109 6538 111
rect 6560 109 6562 111
rect 6566 109 6568 111
rect 6590 109 6592 111
rect 6596 109 6598 111
rect 6620 109 6622 111
rect 6626 109 6628 111
rect 6650 109 6652 111
rect 6656 109 6658 111
rect 6680 109 6682 111
rect 6686 109 6688 111
rect 6710 109 6712 111
rect 6716 109 6718 111
rect 6740 109 6742 111
rect 6746 109 6748 111
rect 4460 106 4462 108
rect 4490 106 4492 108
rect 4520 106 4522 108
rect 4550 106 4552 108
rect 4580 106 4582 108
rect 4610 106 4612 108
rect 4640 106 4642 108
rect 4670 106 4672 108
rect 4700 106 4702 108
rect 4730 106 4732 108
rect 4760 106 4762 108
rect 4790 106 4792 108
rect 4820 106 4822 108
rect 4850 106 4852 108
rect 4880 106 4882 108
rect 4910 106 4912 108
rect 4940 106 4942 108
rect 5060 106 5062 108
rect 5090 106 5092 108
rect 5120 106 5122 108
rect 5150 106 5152 108
rect 5180 106 5182 108
rect 5210 106 5212 108
rect 5240 106 5242 108
rect 5270 106 5272 108
rect 5300 106 5302 108
rect 5330 106 5332 108
rect 5360 106 5362 108
rect 5390 106 5392 108
rect 5420 106 5422 108
rect 5450 106 5452 108
rect 5480 106 5482 108
rect 5510 106 5512 108
rect 5540 106 5542 108
rect 6258 107 6260 109
rect 6288 107 6290 109
rect 6318 107 6320 109
rect 6348 107 6350 109
rect 6378 107 6380 109
rect 6408 107 6410 109
rect 6438 107 6440 109
rect 6468 107 6470 109
rect 6498 107 6500 109
rect 6528 107 6530 109
rect 6558 107 6560 109
rect 6588 107 6590 109
rect 6618 107 6620 109
rect 6648 107 6650 109
rect 6678 107 6680 109
rect 6708 107 6710 109
rect 6738 107 6740 109
rect 4460 100 4462 102
rect 4490 100 4492 102
rect 4520 100 4522 102
rect 4550 100 4552 102
rect 4580 100 4582 102
rect 4610 100 4612 102
rect 4640 100 4642 102
rect 4670 100 4672 102
rect 4700 100 4702 102
rect 4730 100 4732 102
rect 4760 100 4762 102
rect 4790 100 4792 102
rect 4820 100 4822 102
rect 4850 100 4852 102
rect 4880 100 4882 102
rect 4910 100 4912 102
rect 4940 100 4942 102
rect 5060 100 5062 102
rect 5090 100 5092 102
rect 5120 100 5122 102
rect 5150 100 5152 102
rect 5180 100 5182 102
rect 5210 100 5212 102
rect 5240 100 5242 102
rect 5270 100 5272 102
rect 5300 100 5302 102
rect 5330 100 5332 102
rect 5360 100 5362 102
rect 5390 100 5392 102
rect 5420 100 5422 102
rect 5450 100 5452 102
rect 5480 100 5482 102
rect 5510 100 5512 102
rect 5540 100 5542 102
rect 6258 101 6260 103
rect 6288 101 6290 103
rect 6318 101 6320 103
rect 6348 101 6350 103
rect 6378 101 6380 103
rect 6408 101 6410 103
rect 6438 101 6440 103
rect 6468 101 6470 103
rect 6498 101 6500 103
rect 6528 101 6530 103
rect 6558 101 6560 103
rect 6588 101 6590 103
rect 6618 101 6620 103
rect 6648 101 6650 103
rect 6678 101 6680 103
rect 6708 101 6710 103
rect 6738 101 6740 103
rect 3304 98 3306 100
rect 3694 98 3696 100
rect 3904 98 3906 100
rect 4294 98 4296 100
rect 4462 98 4464 100
rect 4468 98 4470 100
rect 4492 98 4494 100
rect 4498 98 4500 100
rect 4522 98 4524 100
rect 4528 98 4530 100
rect 4552 98 4554 100
rect 4558 98 4560 100
rect 4582 98 4584 100
rect 4588 98 4590 100
rect 4612 98 4614 100
rect 4618 98 4620 100
rect 4642 98 4644 100
rect 4648 98 4650 100
rect 4672 98 4674 100
rect 4678 98 4680 100
rect 4702 98 4704 100
rect 4708 98 4710 100
rect 4732 98 4734 100
rect 4738 98 4740 100
rect 4762 98 4764 100
rect 4768 98 4770 100
rect 4792 98 4794 100
rect 4798 98 4800 100
rect 4822 98 4824 100
rect 4828 98 4830 100
rect 4852 98 4854 100
rect 4858 98 4860 100
rect 4882 98 4884 100
rect 4888 98 4890 100
rect 4912 98 4914 100
rect 4918 98 4920 100
rect 4942 98 4944 100
rect 4948 98 4950 100
rect 5062 98 5064 100
rect 5068 98 5070 100
rect 5092 98 5094 100
rect 5098 98 5100 100
rect 5122 98 5124 100
rect 5128 98 5130 100
rect 5152 98 5154 100
rect 5158 98 5160 100
rect 5182 98 5184 100
rect 5188 98 5190 100
rect 5212 98 5214 100
rect 5218 98 5220 100
rect 5242 98 5244 100
rect 5248 98 5250 100
rect 5272 98 5274 100
rect 5278 98 5280 100
rect 5302 98 5304 100
rect 5308 98 5310 100
rect 5332 98 5334 100
rect 5338 98 5340 100
rect 5362 98 5364 100
rect 5368 98 5370 100
rect 5392 98 5394 100
rect 5398 98 5400 100
rect 5422 98 5424 100
rect 5428 98 5430 100
rect 5452 98 5454 100
rect 5458 98 5460 100
rect 5482 98 5484 100
rect 5488 98 5490 100
rect 5512 98 5514 100
rect 5518 98 5520 100
rect 5542 98 5544 100
rect 5548 98 5550 100
rect 6260 99 6262 101
rect 6266 99 6268 101
rect 6290 99 6292 101
rect 6296 99 6298 101
rect 6320 99 6322 101
rect 6326 99 6328 101
rect 6350 99 6352 101
rect 6356 99 6358 101
rect 6380 99 6382 101
rect 6386 99 6388 101
rect 6410 99 6412 101
rect 6416 99 6418 101
rect 6440 99 6442 101
rect 6446 99 6448 101
rect 6470 99 6472 101
rect 6476 99 6478 101
rect 6500 99 6502 101
rect 6506 99 6508 101
rect 6530 99 6532 101
rect 6536 99 6538 101
rect 6560 99 6562 101
rect 6566 99 6568 101
rect 6590 99 6592 101
rect 6596 99 6598 101
rect 6620 99 6622 101
rect 6626 99 6628 101
rect 6650 99 6652 101
rect 6656 99 6658 101
rect 6680 99 6682 101
rect 6686 99 6688 101
rect 6710 99 6712 101
rect 6716 99 6718 101
rect 6740 99 6742 101
rect 6746 99 6748 101
rect 3306 96 3308 98
rect 3692 96 3694 98
rect 3906 96 3908 98
rect 4292 96 4294 98
rect 4470 96 4472 98
rect 4500 96 4502 98
rect 4530 96 4532 98
rect 4560 96 4562 98
rect 4590 96 4592 98
rect 4620 96 4622 98
rect 4650 96 4652 98
rect 4680 96 4682 98
rect 4710 96 4712 98
rect 4740 96 4742 98
rect 4770 96 4772 98
rect 4800 96 4802 98
rect 4830 96 4832 98
rect 4860 96 4862 98
rect 4890 96 4892 98
rect 4920 96 4922 98
rect 4950 96 4952 98
rect 5070 96 5072 98
rect 5100 96 5102 98
rect 5130 96 5132 98
rect 5160 96 5162 98
rect 5190 96 5192 98
rect 5220 96 5222 98
rect 5250 96 5252 98
rect 5280 96 5282 98
rect 5310 96 5312 98
rect 5340 96 5342 98
rect 5370 96 5372 98
rect 5400 96 5402 98
rect 5430 96 5432 98
rect 5460 96 5462 98
rect 5490 96 5492 98
rect 5520 96 5522 98
rect 5550 96 5552 98
rect 5704 96 5706 98
rect 6094 96 6096 98
rect 6268 97 6270 99
rect 6298 97 6300 99
rect 6328 97 6330 99
rect 6358 97 6360 99
rect 6388 97 6390 99
rect 6418 97 6420 99
rect 6448 97 6450 99
rect 6478 97 6480 99
rect 6508 97 6510 99
rect 6538 97 6540 99
rect 6568 97 6570 99
rect 6598 97 6600 99
rect 6628 97 6630 99
rect 6658 97 6660 99
rect 6688 97 6690 99
rect 6718 97 6720 99
rect 6748 97 6750 99
rect 5706 94 5708 96
rect 6092 94 6094 96
rect 4470 90 4472 92
rect 4500 90 4502 92
rect 4530 90 4532 92
rect 4560 90 4562 92
rect 4590 90 4592 92
rect 4620 90 4622 92
rect 4650 90 4652 92
rect 4680 90 4682 92
rect 4710 90 4712 92
rect 4740 90 4742 92
rect 4770 90 4772 92
rect 4800 90 4802 92
rect 4830 90 4832 92
rect 4860 90 4862 92
rect 4890 90 4892 92
rect 4920 90 4922 92
rect 4950 90 4952 92
rect 5070 90 5072 92
rect 5100 90 5102 92
rect 5130 90 5132 92
rect 5160 90 5162 92
rect 5190 90 5192 92
rect 5220 90 5222 92
rect 5250 90 5252 92
rect 5280 90 5282 92
rect 5310 90 5312 92
rect 5340 90 5342 92
rect 5370 90 5372 92
rect 5400 90 5402 92
rect 5430 90 5432 92
rect 5460 90 5462 92
rect 5490 90 5492 92
rect 5520 90 5522 92
rect 5550 90 5552 92
rect 6268 91 6270 93
rect 6298 91 6300 93
rect 6328 91 6330 93
rect 6358 91 6360 93
rect 6388 91 6390 93
rect 6418 91 6420 93
rect 6448 91 6450 93
rect 6478 91 6480 93
rect 6508 91 6510 93
rect 6538 91 6540 93
rect 6568 91 6570 93
rect 6598 91 6600 93
rect 6628 91 6630 93
rect 6658 91 6660 93
rect 6688 91 6690 93
rect 6718 91 6720 93
rect 6748 91 6750 93
rect 4462 88 4464 90
rect 4468 88 4470 90
rect 4492 88 4494 90
rect 4498 88 4500 90
rect 4522 88 4524 90
rect 4528 88 4530 90
rect 4552 88 4554 90
rect 4558 88 4560 90
rect 4582 88 4584 90
rect 4588 88 4590 90
rect 4612 88 4614 90
rect 4618 88 4620 90
rect 4642 88 4644 90
rect 4648 88 4650 90
rect 4672 88 4674 90
rect 4678 88 4680 90
rect 4702 88 4704 90
rect 4708 88 4710 90
rect 4732 88 4734 90
rect 4738 88 4740 90
rect 4762 88 4764 90
rect 4768 88 4770 90
rect 4792 88 4794 90
rect 4798 88 4800 90
rect 4822 88 4824 90
rect 4828 88 4830 90
rect 4852 88 4854 90
rect 4858 88 4860 90
rect 4882 88 4884 90
rect 4888 88 4890 90
rect 4912 88 4914 90
rect 4918 88 4920 90
rect 4942 88 4944 90
rect 4948 88 4950 90
rect 5062 88 5064 90
rect 5068 88 5070 90
rect 5092 88 5094 90
rect 5098 88 5100 90
rect 5122 88 5124 90
rect 5128 88 5130 90
rect 5152 88 5154 90
rect 5158 88 5160 90
rect 5182 88 5184 90
rect 5188 88 5190 90
rect 5212 88 5214 90
rect 5218 88 5220 90
rect 5242 88 5244 90
rect 5248 88 5250 90
rect 5272 88 5274 90
rect 5278 88 5280 90
rect 5302 88 5304 90
rect 5308 88 5310 90
rect 5332 88 5334 90
rect 5338 88 5340 90
rect 5362 88 5364 90
rect 5368 88 5370 90
rect 5392 88 5394 90
rect 5398 88 5400 90
rect 5422 88 5424 90
rect 5428 88 5430 90
rect 5452 88 5454 90
rect 5458 88 5460 90
rect 5482 88 5484 90
rect 5488 88 5490 90
rect 5512 88 5514 90
rect 5518 88 5520 90
rect 5542 88 5544 90
rect 5548 88 5550 90
rect 6260 89 6262 91
rect 6266 89 6268 91
rect 6290 89 6292 91
rect 6296 89 6298 91
rect 6320 89 6322 91
rect 6326 89 6328 91
rect 6350 89 6352 91
rect 6356 89 6358 91
rect 6380 89 6382 91
rect 6386 89 6388 91
rect 6410 89 6412 91
rect 6416 89 6418 91
rect 6440 89 6442 91
rect 6446 89 6448 91
rect 6470 89 6472 91
rect 6476 89 6478 91
rect 6500 89 6502 91
rect 6506 89 6508 91
rect 6530 89 6532 91
rect 6536 89 6538 91
rect 6560 89 6562 91
rect 6566 89 6568 91
rect 6590 89 6592 91
rect 6596 89 6598 91
rect 6620 89 6622 91
rect 6626 89 6628 91
rect 6650 89 6652 91
rect 6656 89 6658 91
rect 6680 89 6682 91
rect 6686 89 6688 91
rect 6710 89 6712 91
rect 6716 89 6718 91
rect 6740 89 6742 91
rect 6746 89 6748 91
rect 4460 86 4462 88
rect 4490 86 4492 88
rect 4520 86 4522 88
rect 4550 86 4552 88
rect 4580 86 4582 88
rect 4610 86 4612 88
rect 4640 86 4642 88
rect 4670 86 4672 88
rect 4700 86 4702 88
rect 4730 86 4732 88
rect 4760 86 4762 88
rect 4790 86 4792 88
rect 4820 86 4822 88
rect 4850 86 4852 88
rect 4880 86 4882 88
rect 4910 86 4912 88
rect 4940 86 4942 88
rect 5060 86 5062 88
rect 5090 86 5092 88
rect 5120 86 5122 88
rect 5150 86 5152 88
rect 5180 86 5182 88
rect 5210 86 5212 88
rect 5240 86 5242 88
rect 5270 86 5272 88
rect 5300 86 5302 88
rect 5330 86 5332 88
rect 5360 86 5362 88
rect 5390 86 5392 88
rect 5420 86 5422 88
rect 5450 86 5452 88
rect 5480 86 5482 88
rect 5510 86 5512 88
rect 5540 86 5542 88
rect 6258 87 6260 89
rect 6288 87 6290 89
rect 6318 87 6320 89
rect 6348 87 6350 89
rect 6378 87 6380 89
rect 6408 87 6410 89
rect 6438 87 6440 89
rect 6468 87 6470 89
rect 6498 87 6500 89
rect 6528 87 6530 89
rect 6558 87 6560 89
rect 6588 87 6590 89
rect 6618 87 6620 89
rect 6648 87 6650 89
rect 6678 87 6680 89
rect 6708 87 6710 89
rect 6738 87 6740 89
rect 4460 80 4462 82
rect 4490 80 4492 82
rect 4520 80 4522 82
rect 4550 80 4552 82
rect 4580 80 4582 82
rect 4610 80 4612 82
rect 4640 80 4642 82
rect 4670 80 4672 82
rect 4700 80 4702 82
rect 4730 80 4732 82
rect 4760 80 4762 82
rect 4790 80 4792 82
rect 4820 80 4822 82
rect 4850 80 4852 82
rect 4880 80 4882 82
rect 4910 80 4912 82
rect 4940 80 4942 82
rect 5060 80 5062 82
rect 5090 80 5092 82
rect 5120 80 5122 82
rect 5150 80 5152 82
rect 5180 80 5182 82
rect 5210 80 5212 82
rect 5240 80 5242 82
rect 5270 80 5272 82
rect 5300 80 5302 82
rect 5330 80 5332 82
rect 5360 80 5362 82
rect 5390 80 5392 82
rect 5420 80 5422 82
rect 5450 80 5452 82
rect 5480 80 5482 82
rect 5510 80 5512 82
rect 5540 80 5542 82
rect 6258 81 6260 83
rect 6288 81 6290 83
rect 6318 81 6320 83
rect 6348 81 6350 83
rect 6378 81 6380 83
rect 6408 81 6410 83
rect 6438 81 6440 83
rect 6468 81 6470 83
rect 6498 81 6500 83
rect 6528 81 6530 83
rect 6558 81 6560 83
rect 6588 81 6590 83
rect 6618 81 6620 83
rect 6648 81 6650 83
rect 6678 81 6680 83
rect 6708 81 6710 83
rect 6738 81 6740 83
rect 4462 78 4464 80
rect 4468 78 4470 80
rect 4492 78 4494 80
rect 4498 78 4500 80
rect 4522 78 4524 80
rect 4528 78 4530 80
rect 4552 78 4554 80
rect 4558 78 4560 80
rect 4582 78 4584 80
rect 4588 78 4590 80
rect 4612 78 4614 80
rect 4618 78 4620 80
rect 4642 78 4644 80
rect 4648 78 4650 80
rect 4672 78 4674 80
rect 4678 78 4680 80
rect 4702 78 4704 80
rect 4708 78 4710 80
rect 4732 78 4734 80
rect 4738 78 4740 80
rect 4762 78 4764 80
rect 4768 78 4770 80
rect 4792 78 4794 80
rect 4798 78 4800 80
rect 4822 78 4824 80
rect 4828 78 4830 80
rect 4852 78 4854 80
rect 4858 78 4860 80
rect 4882 78 4884 80
rect 4888 78 4890 80
rect 4912 78 4914 80
rect 4918 78 4920 80
rect 4942 78 4944 80
rect 4948 78 4950 80
rect 5062 78 5064 80
rect 5068 78 5070 80
rect 5092 78 5094 80
rect 5098 78 5100 80
rect 5122 78 5124 80
rect 5128 78 5130 80
rect 5152 78 5154 80
rect 5158 78 5160 80
rect 5182 78 5184 80
rect 5188 78 5190 80
rect 5212 78 5214 80
rect 5218 78 5220 80
rect 5242 78 5244 80
rect 5248 78 5250 80
rect 5272 78 5274 80
rect 5278 78 5280 80
rect 5302 78 5304 80
rect 5308 78 5310 80
rect 5332 78 5334 80
rect 5338 78 5340 80
rect 5362 78 5364 80
rect 5368 78 5370 80
rect 5392 78 5394 80
rect 5398 78 5400 80
rect 5422 78 5424 80
rect 5428 78 5430 80
rect 5452 78 5454 80
rect 5458 78 5460 80
rect 5482 78 5484 80
rect 5488 78 5490 80
rect 5512 78 5514 80
rect 5518 78 5520 80
rect 5542 78 5544 80
rect 5548 78 5550 80
rect 6260 79 6262 81
rect 6266 79 6268 81
rect 6290 79 6292 81
rect 6296 79 6298 81
rect 6320 79 6322 81
rect 6326 79 6328 81
rect 6350 79 6352 81
rect 6356 79 6358 81
rect 6380 79 6382 81
rect 6386 79 6388 81
rect 6410 79 6412 81
rect 6416 79 6418 81
rect 6440 79 6442 81
rect 6446 79 6448 81
rect 6470 79 6472 81
rect 6476 79 6478 81
rect 6500 79 6502 81
rect 6506 79 6508 81
rect 6530 79 6532 81
rect 6536 79 6538 81
rect 6560 79 6562 81
rect 6566 79 6568 81
rect 6590 79 6592 81
rect 6596 79 6598 81
rect 6620 79 6622 81
rect 6626 79 6628 81
rect 6650 79 6652 81
rect 6656 79 6658 81
rect 6680 79 6682 81
rect 6686 79 6688 81
rect 6710 79 6712 81
rect 6716 79 6718 81
rect 6740 79 6742 81
rect 6746 79 6748 81
rect 4470 76 4472 78
rect 4500 76 4502 78
rect 4530 76 4532 78
rect 4560 76 4562 78
rect 4590 76 4592 78
rect 4620 76 4622 78
rect 4650 76 4652 78
rect 4680 76 4682 78
rect 4710 76 4712 78
rect 4740 76 4742 78
rect 4770 76 4772 78
rect 4800 76 4802 78
rect 4830 76 4832 78
rect 4860 76 4862 78
rect 4890 76 4892 78
rect 4920 76 4922 78
rect 4950 76 4952 78
rect 5070 76 5072 78
rect 5100 76 5102 78
rect 5130 76 5132 78
rect 5160 76 5162 78
rect 5190 76 5192 78
rect 5220 76 5222 78
rect 5250 76 5252 78
rect 5280 76 5282 78
rect 5310 76 5312 78
rect 5340 76 5342 78
rect 5370 76 5372 78
rect 5400 76 5402 78
rect 5430 76 5432 78
rect 5460 76 5462 78
rect 5490 76 5492 78
rect 5520 76 5522 78
rect 5550 76 5552 78
rect 6268 77 6270 79
rect 6298 77 6300 79
rect 6328 77 6330 79
rect 6358 77 6360 79
rect 6388 77 6390 79
rect 6418 77 6420 79
rect 6448 77 6450 79
rect 6478 77 6480 79
rect 6508 77 6510 79
rect 6538 77 6540 79
rect 6568 77 6570 79
rect 6598 77 6600 79
rect 6628 77 6630 79
rect 6658 77 6660 79
rect 6688 77 6690 79
rect 6718 77 6720 79
rect 6748 77 6750 79
rect 4470 70 4472 72
rect 4500 70 4502 72
rect 4530 70 4532 72
rect 4560 70 4562 72
rect 4590 70 4592 72
rect 4620 70 4622 72
rect 4650 70 4652 72
rect 4680 70 4682 72
rect 4710 70 4712 72
rect 4740 70 4742 72
rect 4770 70 4772 72
rect 4800 70 4802 72
rect 4830 70 4832 72
rect 4860 70 4862 72
rect 4890 70 4892 72
rect 4920 70 4922 72
rect 4950 70 4952 72
rect 5070 70 5072 72
rect 5100 70 5102 72
rect 5130 70 5132 72
rect 5160 70 5162 72
rect 5190 70 5192 72
rect 5220 70 5222 72
rect 5250 70 5252 72
rect 5280 70 5282 72
rect 5310 70 5312 72
rect 5340 70 5342 72
rect 5370 70 5372 72
rect 5400 70 5402 72
rect 5430 70 5432 72
rect 5460 70 5462 72
rect 5490 70 5492 72
rect 5520 70 5522 72
rect 5550 70 5552 72
rect 6268 71 6270 73
rect 6298 71 6300 73
rect 6328 71 6330 73
rect 6358 71 6360 73
rect 6388 71 6390 73
rect 6418 71 6420 73
rect 6448 71 6450 73
rect 6478 71 6480 73
rect 6508 71 6510 73
rect 6538 71 6540 73
rect 6568 71 6570 73
rect 6598 71 6600 73
rect 6628 71 6630 73
rect 6658 71 6660 73
rect 6688 71 6690 73
rect 6718 71 6720 73
rect 6748 71 6750 73
rect 4462 68 4464 70
rect 4468 68 4470 70
rect 4492 68 4494 70
rect 4498 68 4500 70
rect 4522 68 4524 70
rect 4528 68 4530 70
rect 4552 68 4554 70
rect 4558 68 4560 70
rect 4582 68 4584 70
rect 4588 68 4590 70
rect 4612 68 4614 70
rect 4618 68 4620 70
rect 4642 68 4644 70
rect 4648 68 4650 70
rect 4672 68 4674 70
rect 4678 68 4680 70
rect 4702 68 4704 70
rect 4708 68 4710 70
rect 4732 68 4734 70
rect 4738 68 4740 70
rect 4762 68 4764 70
rect 4768 68 4770 70
rect 4792 68 4794 70
rect 4798 68 4800 70
rect 4822 68 4824 70
rect 4828 68 4830 70
rect 4852 68 4854 70
rect 4858 68 4860 70
rect 4882 68 4884 70
rect 4888 68 4890 70
rect 4912 68 4914 70
rect 4918 68 4920 70
rect 4942 68 4944 70
rect 4948 68 4950 70
rect 5062 68 5064 70
rect 5068 68 5070 70
rect 5092 68 5094 70
rect 5098 68 5100 70
rect 5122 68 5124 70
rect 5128 68 5130 70
rect 5152 68 5154 70
rect 5158 68 5160 70
rect 5182 68 5184 70
rect 5188 68 5190 70
rect 5212 68 5214 70
rect 5218 68 5220 70
rect 5242 68 5244 70
rect 5248 68 5250 70
rect 5272 68 5274 70
rect 5278 68 5280 70
rect 5302 68 5304 70
rect 5308 68 5310 70
rect 5332 68 5334 70
rect 5338 68 5340 70
rect 5362 68 5364 70
rect 5368 68 5370 70
rect 5392 68 5394 70
rect 5398 68 5400 70
rect 5422 68 5424 70
rect 5428 68 5430 70
rect 5452 68 5454 70
rect 5458 68 5460 70
rect 5482 68 5484 70
rect 5488 68 5490 70
rect 5512 68 5514 70
rect 5518 68 5520 70
rect 5542 68 5544 70
rect 5548 68 5550 70
rect 6260 69 6262 71
rect 6266 69 6268 71
rect 6290 69 6292 71
rect 6296 69 6298 71
rect 6320 69 6322 71
rect 6326 69 6328 71
rect 6350 69 6352 71
rect 6356 69 6358 71
rect 6380 69 6382 71
rect 6386 69 6388 71
rect 6410 69 6412 71
rect 6416 69 6418 71
rect 6440 69 6442 71
rect 6446 69 6448 71
rect 6470 69 6472 71
rect 6476 69 6478 71
rect 6500 69 6502 71
rect 6506 69 6508 71
rect 6530 69 6532 71
rect 6536 69 6538 71
rect 6560 69 6562 71
rect 6566 69 6568 71
rect 6590 69 6592 71
rect 6596 69 6598 71
rect 6620 69 6622 71
rect 6626 69 6628 71
rect 6650 69 6652 71
rect 6656 69 6658 71
rect 6680 69 6682 71
rect 6686 69 6688 71
rect 6710 69 6712 71
rect 6716 69 6718 71
rect 6740 69 6742 71
rect 6746 69 6748 71
rect 4460 66 4462 68
rect 4490 66 4492 68
rect 4520 66 4522 68
rect 4550 66 4552 68
rect 4580 66 4582 68
rect 4610 66 4612 68
rect 4640 66 4642 68
rect 4670 66 4672 68
rect 4700 66 4702 68
rect 4730 66 4732 68
rect 4760 66 4762 68
rect 4790 66 4792 68
rect 4820 66 4822 68
rect 4850 66 4852 68
rect 4880 66 4882 68
rect 4910 66 4912 68
rect 4940 66 4942 68
rect 5060 66 5062 68
rect 5090 66 5092 68
rect 5120 66 5122 68
rect 5150 66 5152 68
rect 5180 66 5182 68
rect 5210 66 5212 68
rect 5240 66 5242 68
rect 5270 66 5272 68
rect 5300 66 5302 68
rect 5330 66 5332 68
rect 5360 66 5362 68
rect 5390 66 5392 68
rect 5420 66 5422 68
rect 5450 66 5452 68
rect 5480 66 5482 68
rect 5510 66 5512 68
rect 5540 66 5542 68
rect 6258 67 6260 69
rect 6288 67 6290 69
rect 6318 67 6320 69
rect 6348 67 6350 69
rect 6378 67 6380 69
rect 6408 67 6410 69
rect 6438 67 6440 69
rect 6468 67 6470 69
rect 6498 67 6500 69
rect 6528 67 6530 69
rect 6558 67 6560 69
rect 6588 67 6590 69
rect 6618 67 6620 69
rect 6648 67 6650 69
rect 6678 67 6680 69
rect 6708 67 6710 69
rect 6738 67 6740 69
rect 2068 60 2078 64
rect 2668 60 2678 64
rect 4460 60 4462 62
rect 4490 60 4492 62
rect 4520 60 4522 62
rect 4550 60 4552 62
rect 4580 60 4582 62
rect 4610 60 4612 62
rect 4640 60 4642 62
rect 4670 60 4672 62
rect 4700 60 4702 62
rect 4730 60 4732 62
rect 4760 60 4762 62
rect 4790 60 4792 62
rect 4820 60 4822 62
rect 4850 60 4852 62
rect 4880 60 4882 62
rect 4910 60 4912 62
rect 4940 60 4942 62
rect 5060 60 5062 62
rect 5090 60 5092 62
rect 5120 60 5122 62
rect 5150 60 5152 62
rect 5180 60 5182 62
rect 5210 60 5212 62
rect 5240 60 5242 62
rect 5270 60 5272 62
rect 5300 60 5302 62
rect 5330 60 5332 62
rect 5360 60 5362 62
rect 5390 60 5392 62
rect 5420 60 5422 62
rect 5450 60 5452 62
rect 5480 60 5482 62
rect 5510 60 5512 62
rect 5540 60 5542 62
rect 6258 61 6260 63
rect 6288 61 6290 63
rect 6318 61 6320 63
rect 6348 61 6350 63
rect 6378 61 6380 63
rect 6408 61 6410 63
rect 6438 61 6440 63
rect 6468 61 6470 63
rect 6498 61 6500 63
rect 6528 61 6530 63
rect 6558 61 6560 63
rect 6588 61 6590 63
rect 6618 61 6620 63
rect 6648 61 6650 63
rect 6678 61 6680 63
rect 6708 61 6710 63
rect 6738 61 6740 63
rect 2068 58 2080 60
rect 2668 58 2680 60
rect 4462 58 4464 60
rect 4468 58 4470 60
rect 4492 58 4494 60
rect 4498 58 4500 60
rect 4522 58 4524 60
rect 4528 58 4530 60
rect 4552 58 4554 60
rect 4558 58 4560 60
rect 4582 58 4584 60
rect 4588 58 4590 60
rect 4612 58 4614 60
rect 4618 58 4620 60
rect 4642 58 4644 60
rect 4648 58 4650 60
rect 4672 58 4674 60
rect 4678 58 4680 60
rect 4702 58 4704 60
rect 4708 58 4710 60
rect 4732 58 4734 60
rect 4738 58 4740 60
rect 4762 58 4764 60
rect 4768 58 4770 60
rect 4792 58 4794 60
rect 4798 58 4800 60
rect 4822 58 4824 60
rect 4828 58 4830 60
rect 4852 58 4854 60
rect 4858 58 4860 60
rect 4882 58 4884 60
rect 4888 58 4890 60
rect 4912 58 4914 60
rect 4918 58 4920 60
rect 4942 58 4944 60
rect 4948 58 4950 60
rect 5062 58 5064 60
rect 5068 58 5070 60
rect 5092 58 5094 60
rect 5098 58 5100 60
rect 5122 58 5124 60
rect 5128 58 5130 60
rect 5152 58 5154 60
rect 5158 58 5160 60
rect 5182 58 5184 60
rect 5188 58 5190 60
rect 5212 58 5214 60
rect 5218 58 5220 60
rect 5242 58 5244 60
rect 5248 58 5250 60
rect 5272 58 5274 60
rect 5278 58 5280 60
rect 5302 58 5304 60
rect 5308 58 5310 60
rect 5332 58 5334 60
rect 5338 58 5340 60
rect 5362 58 5364 60
rect 5368 58 5370 60
rect 5392 58 5394 60
rect 5398 58 5400 60
rect 5422 58 5424 60
rect 5428 58 5430 60
rect 5452 58 5454 60
rect 5458 58 5460 60
rect 5482 58 5484 60
rect 5488 58 5490 60
rect 5512 58 5514 60
rect 5518 58 5520 60
rect 5542 58 5544 60
rect 5548 58 5550 60
rect 6260 59 6262 61
rect 6266 59 6268 61
rect 6290 59 6292 61
rect 6296 59 6298 61
rect 6320 59 6322 61
rect 6326 59 6328 61
rect 6350 59 6352 61
rect 6356 59 6358 61
rect 6380 59 6382 61
rect 6386 59 6388 61
rect 6410 59 6412 61
rect 6416 59 6418 61
rect 6440 59 6442 61
rect 6446 59 6448 61
rect 6470 59 6472 61
rect 6476 59 6478 61
rect 6500 59 6502 61
rect 6506 59 6508 61
rect 6530 59 6532 61
rect 6536 59 6538 61
rect 6560 59 6562 61
rect 6566 59 6568 61
rect 6590 59 6592 61
rect 6596 59 6598 61
rect 6620 59 6622 61
rect 6626 59 6628 61
rect 6650 59 6652 61
rect 6656 59 6658 61
rect 6680 59 6682 61
rect 6686 59 6688 61
rect 6710 59 6712 61
rect 6716 59 6718 61
rect 6740 59 6742 61
rect 6746 59 6748 61
rect 6868 60 6878 64
rect 2076 56 2078 58
rect 2676 56 2678 58
rect 4470 56 4472 58
rect 4500 56 4502 58
rect 4530 56 4532 58
rect 4560 56 4562 58
rect 4590 56 4592 58
rect 4620 56 4622 58
rect 4650 56 4652 58
rect 4680 56 4682 58
rect 4710 56 4712 58
rect 4740 56 4742 58
rect 4770 56 4772 58
rect 4800 56 4802 58
rect 4830 56 4832 58
rect 4860 56 4862 58
rect 4890 56 4892 58
rect 4920 56 4922 58
rect 4950 56 4952 58
rect 5070 56 5072 58
rect 5100 56 5102 58
rect 5130 56 5132 58
rect 5160 56 5162 58
rect 5190 56 5192 58
rect 5220 56 5222 58
rect 5250 56 5252 58
rect 5280 56 5282 58
rect 5310 56 5312 58
rect 5340 56 5342 58
rect 5370 56 5372 58
rect 5400 56 5402 58
rect 5430 56 5432 58
rect 5460 56 5462 58
rect 5490 56 5492 58
rect 5520 56 5522 58
rect 5550 56 5552 58
rect 5686 56 5688 58
rect 5696 56 5698 58
rect 5706 56 5708 58
rect 5716 56 5718 58
rect 5726 56 5728 58
rect 5736 56 5738 58
rect 5746 56 5748 58
rect 5756 56 5758 58
rect 5766 56 5768 58
rect 5776 56 5778 58
rect 5786 56 5788 58
rect 6012 56 6014 58
rect 6022 56 6024 58
rect 6032 56 6034 58
rect 6042 56 6044 58
rect 6052 56 6054 58
rect 6062 56 6064 58
rect 6072 56 6074 58
rect 6082 56 6084 58
rect 6092 56 6094 58
rect 6102 56 6104 58
rect 6112 56 6114 58
rect 6268 57 6270 59
rect 6298 57 6300 59
rect 6328 57 6330 59
rect 6358 57 6360 59
rect 6388 57 6390 59
rect 6418 57 6420 59
rect 6448 57 6450 59
rect 6478 57 6480 59
rect 6508 57 6510 59
rect 6538 57 6540 59
rect 6568 57 6570 59
rect 6598 57 6600 59
rect 6628 57 6630 59
rect 6658 57 6660 59
rect 6688 57 6690 59
rect 6718 57 6720 59
rect 6748 57 6750 59
rect 6868 58 6880 60
rect 6876 56 6878 58
rect 2074 54 2076 56
rect 2674 54 2676 56
rect 5684 54 5686 56
rect 5698 54 5700 56
rect 5704 54 5706 56
rect 5718 54 5720 56
rect 5724 54 5726 56
rect 5738 54 5740 56
rect 5744 54 5746 56
rect 5758 54 5760 56
rect 5764 54 5766 56
rect 5778 54 5780 56
rect 5784 54 5786 56
rect 6014 54 6016 56
rect 6020 54 6022 56
rect 6034 54 6036 56
rect 6040 54 6042 56
rect 6054 54 6056 56
rect 6060 54 6062 56
rect 6074 54 6076 56
rect 6080 54 6082 56
rect 6094 54 6096 56
rect 6100 54 6102 56
rect 6114 54 6116 56
rect 6874 54 6876 56
rect 2068 50 2078 54
rect 2668 50 2678 54
rect 4470 50 4472 52
rect 4500 50 4502 52
rect 4530 50 4532 52
rect 4560 50 4562 52
rect 4590 50 4592 52
rect 4620 50 4622 52
rect 4650 50 4652 52
rect 4680 50 4682 52
rect 4710 50 4712 52
rect 4740 50 4742 52
rect 4770 50 4772 52
rect 4800 50 4802 52
rect 4830 50 4832 52
rect 4860 50 4862 52
rect 4890 50 4892 52
rect 4920 50 4922 52
rect 4950 50 4952 52
rect 5070 50 5072 52
rect 5100 50 5102 52
rect 5130 50 5132 52
rect 5160 50 5162 52
rect 5190 50 5192 52
rect 5220 50 5222 52
rect 5250 50 5252 52
rect 5280 50 5282 52
rect 5310 50 5312 52
rect 5340 50 5342 52
rect 5370 50 5372 52
rect 5400 50 5402 52
rect 5430 50 5432 52
rect 5460 50 5462 52
rect 5490 50 5492 52
rect 5520 50 5522 52
rect 5550 50 5552 52
rect 6268 51 6270 53
rect 6298 51 6300 53
rect 6328 51 6330 53
rect 6358 51 6360 53
rect 6388 51 6390 53
rect 6418 51 6420 53
rect 6448 51 6450 53
rect 6478 51 6480 53
rect 6508 51 6510 53
rect 6538 51 6540 53
rect 6568 51 6570 53
rect 6598 51 6600 53
rect 6628 51 6630 53
rect 6658 51 6660 53
rect 6688 51 6690 53
rect 6718 51 6720 53
rect 6748 51 6750 53
rect 2068 48 2080 50
rect 2668 48 2680 50
rect 4462 48 4464 50
rect 4468 48 4470 50
rect 4492 48 4494 50
rect 4498 48 4500 50
rect 4522 48 4524 50
rect 4528 48 4530 50
rect 4552 48 4554 50
rect 4558 48 4560 50
rect 4582 48 4584 50
rect 4588 48 4590 50
rect 4612 48 4614 50
rect 4618 48 4620 50
rect 4642 48 4644 50
rect 4648 48 4650 50
rect 4672 48 4674 50
rect 4678 48 4680 50
rect 4702 48 4704 50
rect 4708 48 4710 50
rect 4732 48 4734 50
rect 4738 48 4740 50
rect 4762 48 4764 50
rect 4768 48 4770 50
rect 4792 48 4794 50
rect 4798 48 4800 50
rect 4822 48 4824 50
rect 4828 48 4830 50
rect 4852 48 4854 50
rect 4858 48 4860 50
rect 4882 48 4884 50
rect 4888 48 4890 50
rect 4912 48 4914 50
rect 4918 48 4920 50
rect 4942 48 4944 50
rect 4948 48 4950 50
rect 5062 48 5064 50
rect 5068 48 5070 50
rect 5092 48 5094 50
rect 5098 48 5100 50
rect 5122 48 5124 50
rect 5128 48 5130 50
rect 5152 48 5154 50
rect 5158 48 5160 50
rect 5182 48 5184 50
rect 5188 48 5190 50
rect 5212 48 5214 50
rect 5218 48 5220 50
rect 5242 48 5244 50
rect 5248 48 5250 50
rect 5272 48 5274 50
rect 5278 48 5280 50
rect 5302 48 5304 50
rect 5308 48 5310 50
rect 5332 48 5334 50
rect 5338 48 5340 50
rect 5362 48 5364 50
rect 5368 48 5370 50
rect 5392 48 5394 50
rect 5398 48 5400 50
rect 5422 48 5424 50
rect 5428 48 5430 50
rect 5452 48 5454 50
rect 5458 48 5460 50
rect 5482 48 5484 50
rect 5488 48 5490 50
rect 5512 48 5514 50
rect 5518 48 5520 50
rect 5542 48 5544 50
rect 5548 48 5550 50
rect 6260 49 6262 51
rect 6266 49 6268 51
rect 6290 49 6292 51
rect 6296 49 6298 51
rect 6320 49 6322 51
rect 6326 49 6328 51
rect 6350 49 6352 51
rect 6356 49 6358 51
rect 6380 49 6382 51
rect 6386 49 6388 51
rect 6410 49 6412 51
rect 6416 49 6418 51
rect 6440 49 6442 51
rect 6446 49 6448 51
rect 6470 49 6472 51
rect 6476 49 6478 51
rect 6500 49 6502 51
rect 6506 49 6508 51
rect 6530 49 6532 51
rect 6536 49 6538 51
rect 6560 49 6562 51
rect 6566 49 6568 51
rect 6590 49 6592 51
rect 6596 49 6598 51
rect 6620 49 6622 51
rect 6626 49 6628 51
rect 6650 49 6652 51
rect 6656 49 6658 51
rect 6680 49 6682 51
rect 6686 49 6688 51
rect 6710 49 6712 51
rect 6716 49 6718 51
rect 6740 49 6742 51
rect 6746 49 6748 51
rect 6868 50 6878 54
rect 2076 46 2078 48
rect 2676 46 2678 48
rect 4460 46 4462 48
rect 4490 46 4492 48
rect 4520 46 4522 48
rect 4550 46 4552 48
rect 4580 46 4582 48
rect 4610 46 4612 48
rect 4640 46 4642 48
rect 4670 46 4672 48
rect 4700 46 4702 48
rect 4730 46 4732 48
rect 4760 46 4762 48
rect 4790 46 4792 48
rect 4820 46 4822 48
rect 4850 46 4852 48
rect 4880 46 4882 48
rect 4910 46 4912 48
rect 4940 46 4942 48
rect 5060 46 5062 48
rect 5090 46 5092 48
rect 5120 46 5122 48
rect 5150 46 5152 48
rect 5180 46 5182 48
rect 5210 46 5212 48
rect 5240 46 5242 48
rect 5270 46 5272 48
rect 5300 46 5302 48
rect 5330 46 5332 48
rect 5360 46 5362 48
rect 5390 46 5392 48
rect 5420 46 5422 48
rect 5450 46 5452 48
rect 5480 46 5482 48
rect 5510 46 5512 48
rect 5540 46 5542 48
rect 6258 47 6260 49
rect 6288 47 6290 49
rect 6318 47 6320 49
rect 6348 47 6350 49
rect 6378 47 6380 49
rect 6408 47 6410 49
rect 6438 47 6440 49
rect 6468 47 6470 49
rect 6498 47 6500 49
rect 6528 47 6530 49
rect 6558 47 6560 49
rect 6588 47 6590 49
rect 6618 47 6620 49
rect 6648 47 6650 49
rect 6678 47 6680 49
rect 6708 47 6710 49
rect 6738 47 6740 49
rect 6868 48 6880 50
rect 6876 46 6878 48
rect 2074 44 2076 46
rect 2674 44 2676 46
rect 6874 44 6876 46
rect 2068 40 2078 44
rect 2668 40 2678 44
rect 4460 40 4462 42
rect 4490 40 4492 42
rect 4520 40 4522 42
rect 4550 40 4552 42
rect 4580 40 4582 42
rect 4610 40 4612 42
rect 4640 40 4642 42
rect 4670 40 4672 42
rect 4700 40 4702 42
rect 4730 40 4732 42
rect 4760 40 4762 42
rect 4790 40 4792 42
rect 4820 40 4822 42
rect 4850 40 4852 42
rect 4880 40 4882 42
rect 4910 40 4912 42
rect 4940 40 4942 42
rect 5060 40 5062 42
rect 5090 40 5092 42
rect 5120 40 5122 42
rect 5150 40 5152 42
rect 5180 40 5182 42
rect 5210 40 5212 42
rect 5240 40 5242 42
rect 5270 40 5272 42
rect 5300 40 5302 42
rect 5330 40 5332 42
rect 5360 40 5362 42
rect 5390 40 5392 42
rect 5420 40 5422 42
rect 5450 40 5452 42
rect 5480 40 5482 42
rect 5510 40 5512 42
rect 5540 40 5542 42
rect 6258 41 6260 43
rect 6288 41 6290 43
rect 6318 41 6320 43
rect 6348 41 6350 43
rect 6378 41 6380 43
rect 6408 41 6410 43
rect 6438 41 6440 43
rect 6468 41 6470 43
rect 6498 41 6500 43
rect 6528 41 6530 43
rect 6558 41 6560 43
rect 6588 41 6590 43
rect 6618 41 6620 43
rect 6648 41 6650 43
rect 6678 41 6680 43
rect 6708 41 6710 43
rect 6738 41 6740 43
rect 2068 38 2080 40
rect 2668 38 2680 40
rect 4462 38 4464 40
rect 4468 38 4470 40
rect 4492 38 4494 40
rect 4498 38 4500 40
rect 4522 38 4524 40
rect 4528 38 4530 40
rect 4552 38 4554 40
rect 4558 38 4560 40
rect 4582 38 4584 40
rect 4588 38 4590 40
rect 4612 38 4614 40
rect 4618 38 4620 40
rect 4642 38 4644 40
rect 4648 38 4650 40
rect 4672 38 4674 40
rect 4678 38 4680 40
rect 4702 38 4704 40
rect 4708 38 4710 40
rect 4732 38 4734 40
rect 4738 38 4740 40
rect 4762 38 4764 40
rect 4768 38 4770 40
rect 4792 38 4794 40
rect 4798 38 4800 40
rect 4822 38 4824 40
rect 4828 38 4830 40
rect 4852 38 4854 40
rect 4858 38 4860 40
rect 4882 38 4884 40
rect 4888 38 4890 40
rect 4912 38 4914 40
rect 4918 38 4920 40
rect 4942 38 4944 40
rect 4948 38 4950 40
rect 5062 38 5064 40
rect 5068 38 5070 40
rect 5092 38 5094 40
rect 5098 38 5100 40
rect 5122 38 5124 40
rect 5128 38 5130 40
rect 5152 38 5154 40
rect 5158 38 5160 40
rect 5182 38 5184 40
rect 5188 38 5190 40
rect 5212 38 5214 40
rect 5218 38 5220 40
rect 5242 38 5244 40
rect 5248 38 5250 40
rect 5272 38 5274 40
rect 5278 38 5280 40
rect 5302 38 5304 40
rect 5308 38 5310 40
rect 5332 38 5334 40
rect 5338 38 5340 40
rect 5362 38 5364 40
rect 5368 38 5370 40
rect 5392 38 5394 40
rect 5398 38 5400 40
rect 5422 38 5424 40
rect 5428 38 5430 40
rect 5452 38 5454 40
rect 5458 38 5460 40
rect 5482 38 5484 40
rect 5488 38 5490 40
rect 5512 38 5514 40
rect 5518 38 5520 40
rect 5542 38 5544 40
rect 5548 38 5550 40
rect 6260 39 6262 41
rect 6266 39 6268 41
rect 6290 39 6292 41
rect 6296 39 6298 41
rect 6320 39 6322 41
rect 6326 39 6328 41
rect 6350 39 6352 41
rect 6356 39 6358 41
rect 6380 39 6382 41
rect 6386 39 6388 41
rect 6410 39 6412 41
rect 6416 39 6418 41
rect 6440 39 6442 41
rect 6446 39 6448 41
rect 6470 39 6472 41
rect 6476 39 6478 41
rect 6500 39 6502 41
rect 6506 39 6508 41
rect 6530 39 6532 41
rect 6536 39 6538 41
rect 6560 39 6562 41
rect 6566 39 6568 41
rect 6590 39 6592 41
rect 6596 39 6598 41
rect 6620 39 6622 41
rect 6626 39 6628 41
rect 6650 39 6652 41
rect 6656 39 6658 41
rect 6680 39 6682 41
rect 6686 39 6688 41
rect 6710 39 6712 41
rect 6716 39 6718 41
rect 6740 39 6742 41
rect 6746 39 6748 41
rect 6868 40 6878 44
rect 2076 36 2078 38
rect 2676 36 2678 38
rect 4470 36 4472 38
rect 4500 36 4502 38
rect 4530 36 4532 38
rect 4560 36 4562 38
rect 4590 36 4592 38
rect 4620 36 4622 38
rect 4650 36 4652 38
rect 4680 36 4682 38
rect 4710 36 4712 38
rect 4740 36 4742 38
rect 4770 36 4772 38
rect 4800 36 4802 38
rect 4830 36 4832 38
rect 4860 36 4862 38
rect 4890 36 4892 38
rect 4920 36 4922 38
rect 4950 36 4952 38
rect 5070 36 5072 38
rect 5100 36 5102 38
rect 5130 36 5132 38
rect 5160 36 5162 38
rect 5190 36 5192 38
rect 5220 36 5222 38
rect 5250 36 5252 38
rect 5280 36 5282 38
rect 5310 36 5312 38
rect 5340 36 5342 38
rect 5370 36 5372 38
rect 5400 36 5402 38
rect 5430 36 5432 38
rect 5460 36 5462 38
rect 5490 36 5492 38
rect 5520 36 5522 38
rect 5550 36 5552 38
rect 6268 37 6270 39
rect 6298 37 6300 39
rect 6328 37 6330 39
rect 6358 37 6360 39
rect 6388 37 6390 39
rect 6418 37 6420 39
rect 6448 37 6450 39
rect 6478 37 6480 39
rect 6508 37 6510 39
rect 6538 37 6540 39
rect 6568 37 6570 39
rect 6598 37 6600 39
rect 6628 37 6630 39
rect 6658 37 6660 39
rect 6688 37 6690 39
rect 6718 37 6720 39
rect 6748 37 6750 39
rect 6868 38 6880 40
rect 6876 36 6878 38
rect 2074 34 2076 36
rect 2674 34 2676 36
rect 6874 34 6876 36
rect 2578 14 2580 22
rect 2586 14 2590 16
rect 3178 14 3180 22
rect 3186 14 3190 16
rect 5612 14 5622 16
rect 2580 12 2582 14
rect 2584 12 2588 14
rect 2590 12 2592 14
rect 3180 12 3182 14
rect 3184 12 3188 14
rect 3190 12 3192 14
rect 3210 12 3212 14
rect 3788 12 3790 14
rect 3810 12 3812 14
rect 4388 12 4390 14
rect 5610 12 5622 14
rect 6178 14 6188 16
rect 6178 12 6190 14
rect 6210 12 6212 14
rect 6788 12 6790 14
rect 2010 10 2022 12
rect 2046 10 2058 12
rect 2072 10 2084 12
rect 2106 10 2118 12
rect 2474 10 2486 12
rect 2528 10 2540 12
rect 2578 10 2580 12
rect 2610 10 2622 12
rect 2646 10 2658 12
rect 2672 10 2684 12
rect 2706 10 2718 12
rect 3074 10 3086 12
rect 3128 10 3140 12
rect 3178 10 3180 12
rect 3212 10 3214 12
rect 3786 10 3788 12
rect 3812 10 3814 12
rect 4386 10 4388 12
rect 2012 8 2014 10
rect 2054 8 2056 10
rect 2074 8 2076 10
rect 2114 8 2116 10
rect 2476 8 2478 10
rect 2536 8 2538 10
rect 2612 8 2614 10
rect 2654 8 2656 10
rect 2674 8 2676 10
rect 2714 8 2716 10
rect 3076 8 3078 10
rect 3136 8 3138 10
rect 5612 8 5614 12
rect 6186 8 6188 12
rect 6212 10 6214 12
rect 6786 10 6788 12
rect 6810 10 6822 12
rect 6846 10 6858 12
rect 6872 10 6884 12
rect 6906 10 6918 12
rect 6812 8 6814 10
rect 6854 8 6856 10
rect 6874 8 6876 10
rect 6914 8 6916 10
rect 5614 6 5616 8
rect 6184 6 6186 8
rect 2012 4 2014 6
rect 2054 4 2056 6
rect 2074 4 2076 6
rect 2114 4 2116 6
rect 2476 4 2478 6
rect 2536 4 2538 6
rect 2612 4 2614 6
rect 2654 4 2656 6
rect 2674 4 2676 6
rect 2714 4 2716 6
rect 3076 4 3078 6
rect 3136 4 3138 6
rect 6812 4 6814 6
rect 6854 4 6856 6
rect 6874 4 6876 6
rect 6914 4 6916 6
rect 2014 2 2016 4
rect 2052 2 2054 4
rect 2076 2 2078 4
rect 2112 2 2114 4
rect 2478 2 2480 4
rect 2534 2 2536 4
rect 2614 2 2616 4
rect 2652 2 2654 4
rect 2676 2 2678 4
rect 2712 2 2714 4
rect 3078 2 3080 4
rect 3134 2 3136 4
rect 6814 2 6816 4
rect 6852 2 6854 4
rect 6876 2 6878 4
rect 6912 2 6914 4
use PadFC  PadFC_0
timestamp 1570494029
transform 1 0 0 0 1 0
box 660 -6 2006 1340
use PadInC  PadInC_0
timestamp 1570494029
transform 1 0 2000 0 1 0
box -12 -6 606 2000
use PadOut  PadOut_0
timestamp 1570494029
transform 1 0 2600 0 1 0
box -12 -6 606 2000
use PadIO  PadIO_0
timestamp 1570494029
transform 1 0 3200 0 1 0
box -6 -6 606 2000
use PadARef  PadARef_0
timestamp 1570494029
transform 1 0 3800 0 1 0
box -6 -6 606 2000
use PadNC  PadNC_0
timestamp 1570494029
transform 1 0 4400 0 1 0
box -6 -6 606 2000
use PadSpace  PadSpace_0
timestamp 1570494029
transform 1 0 5000 0 1 0
box -6 -6 606 1340
use PadGnd  PadGnd_0
timestamp 1570494029
transform 1 0 6200 0 1 0
box -6 -6 606 2000
use Pad_BidirHE  Pad_BidirHE_0
timestamp 1570494029
transform 1 0 6800 0 1 0
box -12 -6 606 2000
use PadVdd  PadVdd_0
timestamp 1570494029
transform 1 0 5600 0 1 0
box -6 -8 606 2000
<< end >>
