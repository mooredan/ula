magic
tech scmos
timestamp 1550344365
<< metal1 >>
rect 110 40 121 45
use dlyrc_7ns  dlyrc_7ns_0
timestamp 1545342674
transform 1 0 -31 0 1 0
box 31 0 148 79
use dlyrc_7ns  dlyrc_7ns_1
timestamp 1545342674
transform 1 0 86 0 1 0
box 31 0 148 79
<< labels >>
rlabel metal1 s 0 79 0 79 4 vdd
port 3 se
rlabel metal1 s 0 0 0 0 2 vss
port 4 ne
rlabel metal1 s 113 41 113 41 2 n1
rlabel metal1 s 0 43 0 43 2 a
port 2 ne
rlabel metal1 s 227 43 227 43 8 b
port 1 nw
<< end >>
