magic
tech scmos
timestamp 1606713361
<< error_p >>
rect -3800 1000 -3780 1040
rect -3930 980 -3780 1000
rect -3740 940 -3720 1000
<< nwell >>
rect 570 760 1290 2320
<< ntransistor >>
rect -3950 1090 -3890 1200
rect -3950 730 -3890 890
rect 900 10 960 580
<< ptransistor >>
rect -3950 1540 -3890 1800
rect 900 940 960 2140
<< nselect >>
rect -4100 1060 -3350 1280
rect -4100 650 -3730 920
rect 690 -50 1170 640
<< pselect >>
rect -4100 1510 -3740 1830
rect 690 880 1170 2200
<< ndiffusion >>
rect -4070 1170 -3950 1200
rect -4070 1120 -4040 1170
rect -3990 1120 -3950 1170
rect -4070 1090 -3950 1120
rect -3890 1170 -3770 1200
rect -3890 1120 -3850 1170
rect -3800 1120 -3770 1170
rect -3890 1090 -3770 1120
rect -3670 1170 -3510 1220
rect -3670 1120 -3640 1170
rect -3590 1120 -3510 1170
rect -3670 1090 -3510 1120
rect -4070 860 -3950 890
rect -4070 810 -4040 860
rect -3990 810 -3950 860
rect -4070 730 -3950 810
rect -3890 860 -3770 890
rect -3890 810 -3850 860
rect -3800 810 -3770 860
rect -3890 730 -3770 810
rect 750 545 900 580
rect 750 495 785 545
rect 835 495 900 545
rect 750 395 900 495
rect 750 345 785 395
rect 835 345 900 395
rect 750 245 900 345
rect 750 195 785 245
rect 835 195 900 245
rect 750 95 900 195
rect 750 45 785 95
rect 835 45 900 95
rect 750 10 900 45
rect 960 545 1110 580
rect 960 495 1025 545
rect 1075 495 1110 545
rect 960 335 1110 495
rect 960 285 1025 335
rect 1075 285 1110 335
rect 960 155 1110 285
rect 960 105 1025 155
rect 1075 105 1110 155
rect 960 10 1110 105
<< pdiffusion >>
rect 750 2105 900 2140
rect 750 2055 785 2105
rect 835 2055 900 2105
rect 750 1925 900 2055
rect 750 1875 785 1925
rect 835 1875 900 1925
rect -4070 1770 -3950 1800
rect -4070 1720 -4040 1770
rect -3990 1720 -3950 1770
rect -4070 1540 -3950 1720
rect -3890 1770 -3770 1800
rect -3890 1720 -3850 1770
rect -3800 1720 -3770 1770
rect -3890 1540 -3770 1720
rect 750 1775 900 1875
rect 750 1725 785 1775
rect 835 1725 900 1775
rect 750 1625 900 1725
rect 750 1575 785 1625
rect 835 1575 900 1625
rect 750 1475 900 1575
rect 750 1425 785 1475
rect 835 1425 900 1475
rect 750 1325 900 1425
rect 750 1275 785 1325
rect 835 1275 900 1325
rect 750 1175 900 1275
rect 750 1125 785 1175
rect 835 1125 900 1175
rect 750 1025 900 1125
rect 750 975 785 1025
rect 835 975 900 1025
rect 750 940 900 975
rect 960 2045 1110 2140
rect 960 1995 1025 2045
rect 1075 1995 1110 2045
rect 960 1895 1110 1995
rect 960 1845 1025 1895
rect 1075 1845 1110 1895
rect 960 1715 1110 1845
rect 960 1665 1025 1715
rect 1075 1665 1110 1715
rect 960 1535 1110 1665
rect 960 1485 1025 1535
rect 1075 1485 1110 1535
rect 960 1355 1110 1485
rect 960 1305 1025 1355
rect 1075 1305 1110 1355
rect 960 1175 1110 1305
rect 960 1125 1025 1175
rect 1075 1125 1110 1175
rect 960 1025 1110 1125
rect 960 975 1025 1025
rect 1075 975 1110 1025
rect 960 940 1110 975
<< ndcontact >>
rect -4040 1120 -3990 1170
rect -3850 1120 -3800 1170
rect -3640 1120 -3590 1170
rect -4040 810 -3990 860
rect -3850 810 -3800 860
rect 785 495 835 545
rect 785 345 835 395
rect 785 195 835 245
rect 785 45 835 95
rect 1025 495 1075 545
rect 1025 285 1075 335
rect 1025 105 1075 155
<< pdcontact >>
rect 785 2055 835 2105
rect 785 1875 835 1925
rect -4040 1720 -3990 1770
rect -3850 1720 -3800 1770
rect 785 1725 835 1775
rect 785 1575 835 1625
rect 785 1425 835 1475
rect 785 1275 835 1325
rect 785 1125 835 1175
rect 785 975 835 1025
rect 1025 1995 1075 2045
rect 1025 1845 1075 1895
rect 1025 1665 1075 1715
rect 1025 1485 1075 1535
rect 1025 1305 1075 1355
rect 1025 1125 1075 1175
rect 1025 975 1075 1025
<< polysilicon >>
rect 900 2140 960 2205
rect -3950 1800 -3890 1870
rect -3950 1200 -3890 1540
rect -3950 1020 -3890 1090
rect -3950 890 -3890 960
rect 900 850 960 940
rect 750 785 960 850
rect 750 735 815 785
rect 865 735 960 785
rect -3950 660 -3890 730
rect 750 670 960 735
rect 900 580 960 670
rect 900 -55 960 10
<< polycontact >>
rect 815 735 865 785
<< metal1 >>
rect 690 2170 1170 2260
rect 750 2105 870 2170
rect 750 2055 785 2105
rect 835 2055 870 2105
rect 750 1925 870 2055
rect -4060 1850 -3780 1910
rect 750 1875 785 1925
rect 835 1875 870 1925
rect -4060 1770 -3970 1850
rect -4060 1720 -4040 1770
rect -3990 1720 -3970 1770
rect -4060 1700 -3970 1720
rect -3870 1770 -3780 1790
rect -3870 1720 -3850 1770
rect -3800 1720 -3780 1770
rect -4060 1410 -3970 1500
rect -4060 1170 -3970 1190
rect -4060 1120 -4040 1170
rect -3990 1120 -3970 1170
rect -4060 1040 -3970 1120
rect -3870 1170 -3780 1720
rect 750 1775 870 1875
rect 750 1725 785 1775
rect 835 1725 870 1775
rect 750 1625 870 1725
rect 750 1575 785 1625
rect 835 1575 870 1625
rect 750 1475 870 1575
rect 750 1425 785 1475
rect 835 1425 870 1475
rect 750 1325 870 1425
rect 750 1275 785 1325
rect 835 1275 870 1325
rect -3870 1120 -3850 1170
rect -3800 1120 -3780 1170
rect -3870 1100 -3780 1120
rect -3660 1170 -3570 1190
rect -3660 1120 -3640 1170
rect -3590 1120 -3570 1170
rect -3660 1100 -3570 1120
rect 750 1175 870 1275
rect 750 1125 785 1175
rect 835 1125 870 1175
rect -4060 980 -3780 1040
rect 750 1025 870 1125
rect -3740 940 -3590 1000
rect 750 975 785 1025
rect 835 975 870 1025
rect 750 940 870 975
rect 990 2045 1110 2080
rect 990 1995 1025 2045
rect 1075 1995 1110 2045
rect 990 1895 1110 1995
rect 990 1845 1025 1895
rect 1075 1845 1110 1895
rect 990 1715 1110 1845
rect 990 1665 1025 1715
rect 1075 1665 1110 1715
rect 990 1535 1110 1665
rect 990 1485 1025 1535
rect 1075 1485 1110 1535
rect 990 1355 1110 1485
rect 990 1305 1025 1355
rect 1075 1305 1110 1355
rect 990 1175 1110 1305
rect 990 1125 1025 1175
rect 1075 1125 1110 1175
rect 990 1025 1110 1125
rect 990 975 1025 1025
rect 1075 975 1110 1025
rect -4060 860 -3970 880
rect -4060 810 -4040 860
rect -3990 810 -3970 860
rect -4060 790 -3970 810
rect -3870 860 -3780 940
rect -3870 810 -3850 860
rect -3800 810 -3780 860
rect -3870 790 -3780 810
rect 780 785 900 820
rect 780 735 815 785
rect 865 735 900 785
rect 780 700 900 735
rect 750 545 870 580
rect 750 495 785 545
rect 835 495 870 545
rect 750 395 870 495
rect 750 345 785 395
rect 835 345 870 395
rect 750 245 870 345
rect 750 195 785 245
rect 835 195 870 245
rect 750 95 870 195
rect 750 45 785 95
rect 835 45 870 95
rect 990 545 1110 975
rect 990 495 1025 545
rect 1075 495 1110 545
rect 990 335 1110 495
rect 990 285 1025 335
rect 1075 285 1110 335
rect 990 155 1110 285
rect 990 105 1025 155
rect 1075 105 1110 155
rect 990 70 1110 105
rect 750 -20 870 45
rect 690 -110 1170 -20
rect -2320 -740 -2230 -600
rect -2320 -790 -2300 -740
rect -2250 -790 -2230 -740
rect -2320 -900 -2230 -790
rect -2320 -950 -2300 -900
rect -2250 -950 -2230 -900
rect -2320 -1030 -2230 -950
rect -2170 -740 -2080 -610
rect -2170 -790 -2150 -740
rect -2100 -790 -2080 -740
rect -2170 -900 -2080 -790
rect -2170 -950 -2150 -900
rect -2100 -950 -2080 -900
rect -2170 -1010 -2080 -950
<< via1 >>
rect -2300 -790 -2250 -740
rect -2300 -950 -2250 -900
rect -2150 -790 -2100 -740
rect -2150 -950 -2100 -900
<< metal2 >>
rect -2960 2680 330 2770
rect -2960 2520 330 2610
rect -2960 2360 330 2450
rect -2960 2200 330 2290
rect -2960 2040 330 2130
rect -2960 1880 330 1970
rect -2960 1720 330 1810
rect -2960 1560 330 1650
rect -2960 1400 330 1490
rect -2960 1240 330 1330
rect -2960 1080 330 1170
rect -4200 945 -4080 1035
rect -2960 920 330 1010
rect -2960 760 330 850
rect -2960 600 330 690
rect -2960 440 330 530
rect -2960 280 330 370
rect -2960 120 330 210
rect -2960 -40 330 50
rect -2960 -200 330 -110
rect -2960 -360 330 -270
rect -2960 -520 330 -430
rect -2910 -740 -1830 -720
rect -2910 -790 -2815 -740
rect -2765 -790 -2655 -740
rect -2605 -790 -2300 -740
rect -2250 -790 -2150 -740
rect -2100 -790 -1830 -740
rect -2910 -810 -1830 -790
rect -2910 -900 -1830 -880
rect -2910 -950 -2815 -900
rect -2765 -950 -2655 -900
rect -2605 -950 -2300 -900
rect -2250 -950 -2150 -900
rect -2100 -950 -1830 -900
rect -2910 -970 -1830 -950
<< via2 >>
rect -2815 -790 -2765 -740
rect -2655 -790 -2605 -740
rect -2815 -950 -2765 -900
rect -2655 -950 -2605 -900
<< metal3 >>
rect -2830 -720 -2750 -650
rect -2670 -720 -2590 -650
rect -2835 -740 -2745 -720
rect -2835 -790 -2815 -740
rect -2765 -790 -2745 -740
rect -2835 -810 -2745 -790
rect -2675 -740 -2585 -720
rect -2675 -790 -2655 -740
rect -2605 -790 -2585 -740
rect -2675 -810 -2585 -790
rect -2830 -880 -2750 -810
rect -2670 -880 -2590 -810
rect -2835 -900 -2745 -880
rect -2835 -950 -2815 -900
rect -2765 -950 -2745 -900
rect -2835 -970 -2745 -950
rect -2675 -900 -2585 -880
rect -2675 -950 -2655 -900
rect -2605 -950 -2585 -900
rect -2675 -970 -2585 -950
rect -2830 -1030 -2750 -970
rect -2670 -1030 -2590 -970
<< labels >>
flabel nwell 690 820 690 820 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 720 -80 720 -80 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 720 2200 720 2200 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 1050 700 1050 700 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 840 760 840 760 2 FreeSans 400 0 0 0 a
port 2 ne
<< end >>
