`celldefine
module decap4 ();
endmodule
`endcelldefine
