`celldefine
module and2_c (z, a, b);
  output z;
  input  a;
  input  b;

  and G1 (z, a, b);
endmodule
`endcelldefine
