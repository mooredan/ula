magic
tech amic5n
timestamp 1608317707
<< nwell >>
rect -90 870 1320 2430
<< nselect >>
rect 0 60 1200 750
<< pselect >>
rect 30 990 1200 2310
<< ntransistor >>
rect 210 120 270 690
rect 450 120 510 690
rect 930 120 990 690
<< ptransistor >>
rect 240 1050 300 2250
rect 450 1050 510 2250
rect 930 1050 990 2250
<< ndiffusion >>
rect 60 120 210 690
rect 270 120 450 690
rect 510 120 930 690
rect 990 120 1140 690
<< pdiffusion >>
rect 90 1050 240 2250
rect 300 1050 450 2250
rect 510 1050 660 2250
rect 780 1050 930 2250
rect 990 1050 1140 2250
<< polysilicon >>
rect 240 2250 300 2310
rect 450 2250 510 2310
rect 930 2250 990 2310
rect 240 960 300 1050
rect 60 780 300 960
rect 450 960 510 1050
rect 930 960 990 1050
rect 450 780 660 960
rect 780 780 990 960
rect 210 690 270 780
rect 450 690 510 780
rect 930 690 990 780
rect 210 60 270 120
rect 450 60 510 120
rect 930 60 990 120
<< pdcontact >>
rect 125 2165 175 2215
<< pdcontact >>
rect 815 2165 865 2215
<< pdcontact >>
rect 575 2105 625 2155
<< pdcontact >>
rect 1055 2105 1105 2155
<< pdcontact >>
rect 125 1985 175 2035
<< pdcontact >>
rect 815 2015 865 2065
<< pdcontact >>
rect 575 1955 625 2005
<< pdcontact >>
rect 1055 1955 1105 2005
<< pdcontact >>
rect 125 1835 175 1885
<< pdcontact >>
rect 815 1865 865 1915
<< pdcontact >>
rect 575 1775 625 1825
<< pdcontact >>
rect 1055 1775 1105 1825
<< pdcontact >>
rect 125 1685 175 1735
<< pdcontact >>
rect 815 1715 865 1765
<< pdcontact >>
rect 575 1595 625 1645
<< pdcontact >>
rect 125 1535 175 1585
<< pdcontact >>
rect 815 1565 865 1615
<< pdcontact >>
rect 1055 1595 1105 1645
<< pdcontact >>
rect 125 1385 175 1435
<< pdcontact >>
rect 575 1415 625 1465
<< pdcontact >>
rect 815 1415 865 1465
<< pdcontact >>
rect 1055 1415 1105 1465
<< pdcontact >>
rect 125 1235 175 1285
<< pdcontact >>
rect 575 1235 625 1285
<< pdcontact >>
rect 815 1265 865 1315
<< pdcontact >>
rect 1055 1235 1105 1285
<< pdcontact >>
rect 125 1085 175 1135
<< pdcontact >>
rect 575 1085 625 1135
<< pdcontact >>
rect 1055 1085 1105 1135
<< polycontact >>
rect 125 845 175 895
<< polycontact >>
rect 545 845 595 895
<< polycontact >>
rect 845 845 895 895
<< ndcontact >>
rect 95 605 145 655
<< ndcontact >>
rect 335 605 385 655
<< ndcontact >>
rect 575 605 625 655
<< ndcontact >>
rect 815 605 865 655
<< ndcontact >>
rect 1055 605 1105 655
<< ndcontact >>
rect 95 455 145 505
<< ndcontact >>
rect 575 455 625 505
<< ndcontact >>
rect 815 455 865 505
<< ndcontact >>
rect 335 395 385 445
<< ndcontact >>
rect 1055 395 1105 445
<< ndcontact >>
rect 95 305 145 355
<< ndcontact >>
rect 575 305 625 355
<< ndcontact >>
rect 815 305 865 355
<< ndcontact >>
rect 335 215 385 265
<< ndcontact >>
rect 1055 215 1105 265
<< ndcontact >>
rect 95 155 145 205
<< ndcontact >>
rect 575 155 625 205
<< ndcontact >>
rect 815 155 865 205
<< metal1 >>
rect 0 2280 1200 2370
rect 90 1050 210 2280
rect 540 1140 660 2190
rect 780 1230 900 2280
rect 300 1020 930 1140
rect 90 810 210 930
rect 60 90 180 690
rect 300 180 420 1020
rect 510 810 630 930
rect 810 810 930 1020
rect 540 90 900 690
rect 1020 180 1140 2190
rect 0 0 1200 90
<< labels >>
flabel nwell  0 930 0 930 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 30 30 30 30 2 FreeSans 400 0 0 0 vss
port 5 ne
flabel metal1 s 30 2310 30 2310 2 FreeSans 400 0 0 0 vdd
port 4 ne
flabel metal1 s 570 870 570 870 2 FreeSans 400 0 0 0 b
port 3 ne
flabel metal1 s 150 870 150 870 2 FreeSans 400 0 0 0 a
port 2 ne
flabel metal1 s 1080 810 1080 810 2 FreeSans 400 0 0 0 z
port 1 ne
flabel pdiffusion s 360 1620 360 1620 2 FreeSans 400 0 0 0 x1
flabel metal1 s 690 1050 690 1050 2 FreeSans 400 0 0 0 n1
<< checkpaint >>
rect -100 -10 1330 2440
<< end >>
