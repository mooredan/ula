magic
tech amic5n
timestamp 1625072543
<< nwell >>
rect -130 550 880 1495
<< ntransistor >>
rect 225 95 285 400
rect 465 95 525 400
<< ptransistor >>
rect 225 705 285 1345
rect 465 705 525 1345
<< nselect >>
rect -10 0 760 430
<< pselect >>
rect -10 670 760 1440
<< ndiffusion >>
rect 105 370 225 400
rect 105 320 135 370
rect 185 320 225 370
rect 105 175 225 320
rect 105 125 135 175
rect 185 125 225 175
rect 105 95 225 125
rect 285 95 465 400
rect 525 345 645 400
rect 525 295 565 345
rect 615 295 645 345
rect 525 185 645 295
rect 525 135 565 185
rect 615 135 645 185
rect 525 95 645 135
<< pdiffusion >>
rect 105 1315 225 1345
rect 105 1265 135 1315
rect 185 1265 225 1315
rect 105 1215 225 1265
rect 105 1165 135 1215
rect 185 1165 225 1215
rect 105 1085 225 1165
rect 105 1035 135 1085
rect 185 1035 225 1085
rect 105 950 225 1035
rect 105 900 135 950
rect 185 900 225 950
rect 105 830 225 900
rect 105 780 135 830
rect 185 780 225 830
rect 105 705 225 780
rect 285 1315 465 1345
rect 285 1265 350 1315
rect 400 1265 465 1315
rect 285 1185 465 1265
rect 285 1135 350 1185
rect 400 1135 465 1185
rect 285 1085 465 1135
rect 285 1035 350 1085
rect 400 1035 465 1085
rect 285 985 465 1035
rect 285 935 350 985
rect 400 935 465 985
rect 285 885 465 935
rect 285 835 350 885
rect 400 835 465 885
rect 285 785 465 835
rect 285 735 350 785
rect 400 735 465 785
rect 285 705 465 735
rect 525 1315 645 1345
rect 525 1265 565 1315
rect 615 1265 645 1315
rect 525 1215 645 1265
rect 525 1165 565 1215
rect 615 1165 645 1215
rect 525 1115 645 1165
rect 525 1065 565 1115
rect 615 1065 645 1115
rect 525 1015 645 1065
rect 525 965 565 1015
rect 615 965 645 1015
rect 525 915 645 965
rect 525 865 565 915
rect 615 865 645 915
rect 525 815 645 865
rect 525 765 565 815
rect 615 765 645 815
rect 525 705 645 765
<< ndcontact >>
rect 135 320 185 370
rect 135 125 185 175
rect 565 295 615 345
rect 565 135 615 185
<< pdcontact >>
rect 135 1265 185 1315
rect 135 1165 185 1215
rect 135 1035 185 1085
rect 135 900 185 950
rect 135 780 185 830
rect 350 1265 400 1315
rect 350 1135 400 1185
rect 350 1035 400 1085
rect 350 935 400 985
rect 350 835 400 885
rect 350 735 400 785
rect 565 1265 615 1315
rect 565 1165 615 1215
rect 565 1065 615 1115
rect 565 965 615 1015
rect 565 865 615 915
rect 565 765 615 815
<< polysilicon >>
rect 225 1345 285 1410
rect 465 1345 525 1410
rect 225 685 285 705
rect 115 665 285 685
rect 115 615 135 665
rect 185 615 285 665
rect 115 595 285 615
rect 225 400 285 595
rect 465 525 525 705
rect 465 505 635 525
rect 465 455 565 505
rect 615 455 635 505
rect 465 435 635 455
rect 465 400 525 435
rect 225 30 285 95
rect 465 30 525 95
<< polycontact >>
rect 135 615 185 665
rect 565 455 615 505
<< metal1 >>
rect 0 1395 750 1485
rect 115 1315 205 1395
rect 115 1265 135 1315
rect 185 1265 205 1315
rect 115 1215 205 1265
rect 115 1165 135 1215
rect 185 1165 205 1215
rect 115 1085 205 1165
rect 115 1035 135 1085
rect 185 1035 205 1085
rect 115 950 205 1035
rect 115 900 135 950
rect 185 900 205 950
rect 115 830 205 900
rect 115 780 135 830
rect 185 780 205 830
rect 115 760 205 780
rect 330 1315 420 1335
rect 330 1265 350 1315
rect 400 1265 420 1315
rect 330 1185 420 1265
rect 330 1135 350 1185
rect 400 1135 420 1185
rect 330 1085 420 1135
rect 330 1035 350 1085
rect 400 1035 420 1085
rect 330 985 420 1035
rect 330 935 350 985
rect 400 935 420 985
rect 330 885 420 935
rect 330 835 350 885
rect 400 835 420 885
rect 330 785 420 835
rect 330 735 350 785
rect 400 735 420 785
rect 545 1315 635 1395
rect 545 1265 565 1315
rect 615 1265 635 1315
rect 545 1215 635 1265
rect 545 1165 565 1215
rect 615 1165 635 1215
rect 545 1115 635 1165
rect 545 1065 565 1115
rect 615 1065 635 1115
rect 545 1015 635 1065
rect 545 965 565 1015
rect 615 965 635 1015
rect 545 915 635 965
rect 545 865 565 915
rect 615 865 635 915
rect 545 815 635 865
rect 545 765 565 815
rect 615 765 635 815
rect 545 745 635 765
rect 30 665 205 685
rect 30 615 135 665
rect 185 615 205 665
rect 30 595 205 615
rect 115 370 205 390
rect 115 320 135 370
rect 185 320 205 370
rect 115 175 205 320
rect 330 365 420 735
rect 545 505 720 525
rect 545 455 565 505
rect 615 455 720 505
rect 545 435 720 455
rect 330 345 635 365
rect 330 295 565 345
rect 615 295 635 345
rect 330 275 635 295
rect 115 125 135 175
rect 185 125 205 175
rect 115 45 205 125
rect 545 185 635 275
rect 545 135 565 185
rect 615 135 635 185
rect 545 105 635 135
rect 0 -45 750 45
<< labels >>
flabel metal1 s 360 470 360 470 2 FreeSans 400 0 0 0 z
port 0 ne
flabel metal1 s 616 445 616 445 2 FreeSans 400 0 0 0 b
port 2 ne
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel nwell 5 585 5 585 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 135 605 135 605 2 FreeSans 400 0 0 0 a
port 1 ne
<< properties >>
string LEFclass CORE
string LEFsite core
string FIXED_BBOX 0 0 750 1440
string LEFsymmetry X Y
<< end >>
