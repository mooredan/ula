magic
tech amic5n
timestamp 1624378881
<< nwell >>
rect -130 550 1330 1495
<< ntransistor >>
rect 205 95 265 400
rect 595 125 655 400
rect 785 125 845 400
rect 975 125 1035 400
<< ptransistor >>
rect 205 705 265 1345
rect 595 705 655 1290
rect 785 705 845 1290
rect 975 705 1035 1290
<< nselect >>
rect -10 0 1210 430
<< pselect >>
rect -10 670 1210 1440
<< ndiffusion >>
rect 85 370 205 400
rect 85 320 115 370
rect 165 320 205 370
rect 85 175 205 320
rect 85 125 115 175
rect 165 125 205 175
rect 85 95 205 125
rect 265 370 385 400
rect 265 320 305 370
rect 355 320 385 370
rect 265 175 385 320
rect 265 125 305 175
rect 355 125 385 175
rect 475 370 595 400
rect 475 320 505 370
rect 555 320 595 370
rect 475 205 595 320
rect 475 155 505 205
rect 555 155 595 205
rect 475 125 595 155
rect 655 370 785 400
rect 655 320 695 370
rect 745 320 785 370
rect 655 205 785 320
rect 655 155 695 205
rect 745 155 785 205
rect 655 125 785 155
rect 845 345 975 400
rect 845 295 885 345
rect 935 295 975 345
rect 845 205 975 295
rect 845 155 885 205
rect 935 155 975 205
rect 845 125 975 155
rect 1035 370 1155 400
rect 1035 320 1075 370
rect 1125 320 1155 370
rect 1035 205 1155 320
rect 1035 155 1075 205
rect 1125 155 1155 205
rect 1035 125 1155 155
rect 265 95 385 125
<< pdiffusion >>
rect 85 1315 205 1345
rect 85 1265 115 1315
rect 165 1265 205 1315
rect 85 1215 205 1265
rect 85 1165 115 1215
rect 165 1165 205 1215
rect 85 1115 205 1165
rect 85 1065 115 1115
rect 165 1065 205 1115
rect 85 1015 205 1065
rect 85 965 115 1015
rect 165 965 205 1015
rect 85 915 205 965
rect 85 865 115 915
rect 165 865 205 915
rect 85 815 205 865
rect 85 765 115 815
rect 165 765 205 815
rect 85 705 205 765
rect 265 1315 385 1345
rect 265 1265 305 1315
rect 355 1265 385 1315
rect 265 1185 385 1265
rect 265 1135 305 1185
rect 355 1135 385 1185
rect 265 1085 385 1135
rect 265 1035 305 1085
rect 355 1035 385 1085
rect 265 985 385 1035
rect 265 935 305 985
rect 355 935 385 985
rect 265 885 385 935
rect 265 835 305 885
rect 355 835 385 885
rect 265 785 385 835
rect 265 735 305 785
rect 355 735 385 785
rect 265 705 385 735
rect 475 1260 595 1290
rect 475 1210 505 1260
rect 555 1210 595 1260
rect 475 1115 595 1210
rect 475 1065 505 1115
rect 555 1065 595 1115
rect 475 1015 595 1065
rect 475 965 505 1015
rect 555 965 595 1015
rect 475 915 595 965
rect 475 865 505 915
rect 555 865 595 915
rect 475 815 595 865
rect 475 765 505 815
rect 555 765 595 815
rect 475 705 595 765
rect 655 1260 785 1290
rect 655 1210 695 1260
rect 745 1210 785 1260
rect 655 1080 785 1210
rect 655 1030 695 1080
rect 745 1030 785 1080
rect 655 980 785 1030
rect 655 930 695 980
rect 745 930 785 980
rect 655 825 785 930
rect 655 775 695 825
rect 745 775 785 825
rect 655 705 785 775
rect 845 1260 975 1290
rect 845 1210 885 1260
rect 935 1210 975 1260
rect 845 1115 975 1210
rect 845 1065 885 1115
rect 935 1065 975 1115
rect 845 975 975 1065
rect 845 925 885 975
rect 935 925 975 975
rect 845 705 975 925
rect 1035 1260 1155 1290
rect 1035 1210 1075 1260
rect 1125 1210 1155 1260
rect 1035 1085 1155 1210
rect 1035 1035 1075 1085
rect 1125 1035 1155 1085
rect 1035 985 1155 1035
rect 1035 935 1075 985
rect 1125 935 1155 985
rect 1035 885 1155 935
rect 1035 835 1075 885
rect 1125 835 1155 885
rect 1035 785 1155 835
rect 1035 735 1075 785
rect 1125 735 1155 785
rect 1035 705 1155 735
<< ndcontact >>
rect 115 320 165 370
rect 115 125 165 175
rect 305 320 355 370
rect 305 125 355 175
rect 505 320 555 370
rect 505 155 555 205
rect 695 320 745 370
rect 695 155 745 205
rect 885 295 935 345
rect 885 155 935 205
rect 1075 320 1125 370
rect 1075 155 1125 205
<< pdcontact >>
rect 115 1265 165 1315
rect 115 1165 165 1215
rect 115 1065 165 1115
rect 115 965 165 1015
rect 115 865 165 915
rect 115 765 165 815
rect 305 1265 355 1315
rect 305 1135 355 1185
rect 305 1035 355 1085
rect 305 935 355 985
rect 305 835 355 885
rect 305 735 355 785
rect 505 1210 555 1260
rect 505 1065 555 1115
rect 505 965 555 1015
rect 505 865 555 915
rect 505 765 555 815
rect 695 1210 745 1260
rect 695 1030 745 1080
rect 695 930 745 980
rect 695 775 745 825
rect 885 1210 935 1260
rect 885 1065 935 1115
rect 885 925 935 975
rect 1075 1210 1125 1260
rect 1075 1035 1125 1085
rect 1075 935 1125 985
rect 1075 835 1125 885
rect 1075 735 1125 785
<< polysilicon >>
rect 205 1345 265 1410
rect 595 1290 655 1355
rect 785 1290 845 1355
rect 975 1290 1035 1355
rect 205 685 265 705
rect 595 685 655 705
rect 785 685 845 705
rect 975 685 1035 705
rect 95 665 265 685
rect 95 615 115 665
rect 165 615 265 665
rect 95 595 265 615
rect 485 665 1035 685
rect 485 615 505 665
rect 555 615 605 665
rect 655 615 705 665
rect 755 615 805 665
rect 855 615 905 665
rect 955 615 1035 665
rect 485 595 1035 615
rect 205 400 265 595
rect 595 400 655 595
rect 785 400 845 595
rect 975 400 1035 595
rect 205 30 265 95
rect 595 60 655 125
rect 785 60 845 125
rect 975 60 1035 125
<< polycontact >>
rect 115 615 165 665
rect 505 615 555 665
rect 605 615 655 665
rect 705 615 755 665
rect 805 615 855 665
rect 905 615 955 665
<< metal1 >>
rect 0 1395 1200 1485
rect 95 1315 185 1395
rect 95 1265 115 1315
rect 165 1265 185 1315
rect 95 1215 185 1265
rect 95 1165 115 1215
rect 165 1165 185 1215
rect 95 1115 185 1165
rect 95 1065 115 1115
rect 165 1065 185 1115
rect 95 1015 185 1065
rect 95 965 115 1015
rect 165 965 185 1015
rect 95 915 185 965
rect 95 865 115 915
rect 165 865 185 915
rect 95 815 185 865
rect 95 765 115 815
rect 165 765 185 815
rect 95 745 185 765
rect 285 1315 375 1335
rect 285 1265 305 1315
rect 355 1265 375 1315
rect 285 1185 375 1265
rect 285 1135 305 1185
rect 355 1135 375 1185
rect 285 1085 375 1135
rect 285 1035 305 1085
rect 355 1035 375 1085
rect 285 985 375 1035
rect 285 935 305 985
rect 355 935 375 985
rect 285 885 375 935
rect 285 835 305 885
rect 355 835 375 885
rect 285 785 375 835
rect 285 735 305 785
rect 355 735 375 785
rect 485 1260 575 1395
rect 485 1210 505 1260
rect 555 1210 575 1260
rect 485 1115 575 1210
rect 485 1065 505 1115
rect 555 1065 575 1115
rect 485 1015 575 1065
rect 485 965 505 1015
rect 555 965 575 1015
rect 485 915 575 965
rect 485 865 505 915
rect 555 865 575 915
rect 485 815 575 865
rect 485 765 505 815
rect 555 765 575 815
rect 485 745 575 765
rect 675 1260 765 1280
rect 675 1210 695 1260
rect 745 1210 765 1260
rect 675 1080 765 1210
rect 675 1030 695 1080
rect 745 1030 765 1080
rect 675 980 765 1030
rect 675 930 695 980
rect 745 930 765 980
rect 675 845 765 930
rect 865 1260 955 1395
rect 865 1210 885 1260
rect 935 1210 955 1260
rect 865 1115 955 1210
rect 865 1065 885 1115
rect 935 1065 955 1115
rect 865 975 955 1065
rect 865 925 885 975
rect 935 925 955 975
rect 865 905 955 925
rect 1055 1260 1145 1280
rect 1055 1210 1075 1260
rect 1125 1210 1145 1260
rect 1055 1085 1145 1210
rect 1055 1035 1075 1085
rect 1125 1035 1145 1085
rect 1055 985 1145 1035
rect 1055 935 1075 985
rect 1125 935 1145 985
rect 1055 885 1145 935
rect 1055 845 1075 885
rect 675 835 1075 845
rect 1125 835 1145 885
rect 675 825 1145 835
rect 675 775 695 825
rect 745 785 1145 825
rect 745 775 1075 785
rect 675 755 1075 775
rect 285 685 375 735
rect 1055 735 1075 755
rect 1125 735 1145 785
rect 95 665 185 685
rect 95 615 115 665
rect 165 615 185 665
rect 95 595 185 615
rect 285 665 975 685
rect 285 615 505 665
rect 555 615 605 665
rect 655 615 705 665
rect 755 615 805 665
rect 855 615 905 665
rect 955 615 975 665
rect 285 595 975 615
rect 95 370 185 390
rect 95 320 115 370
rect 165 320 185 370
rect 95 175 185 320
rect 95 125 115 175
rect 165 125 185 175
rect 95 45 185 125
rect 285 370 375 595
rect 1055 525 1145 735
rect 675 435 1145 525
rect 285 320 305 370
rect 355 320 375 370
rect 285 175 375 320
rect 285 125 305 175
rect 355 125 375 175
rect 285 105 375 125
rect 485 370 575 390
rect 485 320 505 370
rect 555 320 575 370
rect 485 205 575 320
rect 485 155 505 205
rect 555 155 575 205
rect 485 45 575 155
rect 675 370 765 435
rect 675 320 695 370
rect 745 320 765 370
rect 1055 370 1145 435
rect 675 205 765 320
rect 675 155 695 205
rect 745 155 765 205
rect 675 135 765 155
rect 865 345 955 365
rect 865 295 885 345
rect 935 295 955 345
rect 865 205 955 295
rect 865 155 885 205
rect 935 155 955 205
rect 865 45 955 155
rect 1055 320 1075 370
rect 1125 320 1145 370
rect 1055 205 1145 320
rect 1055 155 1075 205
rect 1125 155 1145 205
rect 1055 135 1145 155
rect 0 -45 1200 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 200 0 0 0 vss
port 3 ne
flabel metal1 s 75 1415 75 1415 2 FreeSans 400 0 0 0 vdd
port 2 ne
flabel metal1 s 1095 485 1095 485 2 FreeSans 400 0 0 0 z
port 0 ne
flabel nwell 385 560 385 560 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 115 605 115 605 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 310 470 310 470 2 FreeSans 200 0 0 0 x1
<< properties >>
string FIXED_BBOX 0 0 1200 1440
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
