magic
tech amic5n
timestamp 1624387535
<< nwell >>
rect -130 550 1030 1495
<< ntransistor >>
rect 295 125 355 400
rect 485 125 545 400
rect 675 125 735 400
<< ptransistor >>
rect 295 705 355 1290
rect 485 705 545 1290
rect 675 705 735 1290
<< nselect >>
rect 10 765 175 1290
rect -10 350 910 430
rect 175 125 910 350
rect -10 0 910 125
<< pselect >>
rect -10 1290 910 1440
rect 175 765 910 1290
rect -10 670 910 765
rect 10 125 175 350
<< ndiffusion >>
rect 175 370 295 400
rect 175 320 205 370
rect 255 320 295 370
rect 175 205 295 320
rect 175 155 205 205
rect 255 155 295 205
rect 175 125 295 155
rect 355 370 485 400
rect 355 320 395 370
rect 445 320 485 370
rect 355 205 485 320
rect 355 155 395 205
rect 445 155 485 205
rect 355 125 485 155
rect 545 345 675 400
rect 545 295 585 345
rect 635 295 675 345
rect 545 205 675 295
rect 545 155 585 205
rect 635 155 675 205
rect 545 125 675 155
rect 735 370 855 400
rect 735 320 775 370
rect 825 320 855 370
rect 735 205 855 320
rect 735 155 775 205
rect 825 155 855 205
rect 735 125 855 155
<< pdiffusion >>
rect 175 1260 295 1290
rect 175 1210 205 1260
rect 255 1210 295 1260
rect 175 1115 295 1210
rect 175 1065 205 1115
rect 255 1065 295 1115
rect 175 1015 295 1065
rect 175 965 205 1015
rect 255 965 295 1015
rect 175 915 295 965
rect 175 865 205 915
rect 255 865 295 915
rect 175 815 295 865
rect 175 765 205 815
rect 255 765 295 815
rect 175 705 295 765
rect 355 1260 485 1290
rect 355 1210 395 1260
rect 445 1210 485 1260
rect 355 1080 485 1210
rect 355 1030 395 1080
rect 445 1030 485 1080
rect 355 980 485 1030
rect 355 930 395 980
rect 445 930 485 980
rect 355 825 485 930
rect 355 775 395 825
rect 445 775 485 825
rect 355 705 485 775
rect 545 1260 675 1290
rect 545 1210 585 1260
rect 635 1210 675 1260
rect 545 1115 675 1210
rect 545 1065 585 1115
rect 635 1065 675 1115
rect 545 975 675 1065
rect 545 925 585 975
rect 635 925 675 975
rect 545 705 675 925
rect 735 1260 855 1290
rect 735 1210 775 1260
rect 825 1210 855 1260
rect 735 1085 855 1210
rect 735 1035 775 1085
rect 825 1035 855 1085
rect 735 985 855 1035
rect 735 935 775 985
rect 825 935 855 985
rect 735 885 855 935
rect 735 835 775 885
rect 825 835 855 885
rect 735 785 855 835
rect 735 735 775 785
rect 825 735 855 785
rect 735 705 855 735
<< psubstratepdiff >>
rect 60 320 175 350
rect 60 270 90 320
rect 140 270 175 320
rect 60 205 175 270
rect 60 155 90 205
rect 140 155 175 205
rect 60 125 175 155
<< nsubstratendiff >>
rect 60 1260 175 1290
rect 60 1210 95 1260
rect 145 1210 175 1260
rect 60 1160 175 1210
rect 60 1110 90 1160
rect 140 1110 175 1160
rect 60 1060 175 1110
rect 60 1010 90 1060
rect 140 1010 175 1060
rect 60 960 175 1010
rect 60 910 90 960
rect 140 910 175 960
rect 60 855 175 910
rect 60 805 90 855
rect 140 805 175 855
rect 60 765 175 805
<< nsubstratencontact >>
rect 95 1210 145 1260
rect 90 1110 140 1160
rect 90 1010 140 1060
rect 90 910 140 960
rect 90 805 140 855
<< psubstratepcontact >>
rect 90 270 140 320
rect 90 155 140 205
<< ndcontact >>
rect 205 320 255 370
rect 205 155 255 205
rect 395 320 445 370
rect 395 155 445 205
rect 585 295 635 345
rect 585 155 635 205
rect 775 320 825 370
rect 775 155 825 205
<< pdcontact >>
rect 205 1210 255 1260
rect 205 1065 255 1115
rect 205 965 255 1015
rect 205 865 255 915
rect 205 765 255 815
rect 395 1210 445 1260
rect 395 1030 445 1080
rect 395 930 445 980
rect 395 775 445 825
rect 585 1210 635 1260
rect 585 1065 635 1115
rect 585 925 635 975
rect 775 1210 825 1260
rect 775 1035 825 1085
rect 775 935 825 985
rect 775 835 825 885
rect 775 735 825 785
<< polysilicon >>
rect 295 1290 355 1355
rect 485 1290 545 1355
rect 675 1290 735 1355
rect 295 685 355 705
rect 485 685 545 705
rect 675 685 735 705
rect 185 665 735 685
rect 185 615 205 665
rect 255 615 305 665
rect 355 615 405 665
rect 455 615 505 665
rect 555 615 605 665
rect 655 615 735 665
rect 185 595 735 615
rect 295 400 355 595
rect 485 400 545 595
rect 675 400 735 595
rect 295 60 355 125
rect 485 60 545 125
rect 675 60 735 125
<< polycontact >>
rect 205 615 255 665
rect 305 615 355 665
rect 405 615 455 665
rect 505 615 555 665
rect 605 615 655 665
<< metal1 >>
rect 0 1395 900 1485
rect 70 1260 275 1395
rect 70 1210 95 1260
rect 145 1210 205 1260
rect 255 1210 275 1260
rect 70 1160 275 1210
rect 70 1110 90 1160
rect 140 1115 275 1160
rect 140 1110 205 1115
rect 70 1065 205 1110
rect 255 1065 275 1115
rect 70 1060 275 1065
rect 70 1010 90 1060
rect 140 1015 275 1060
rect 140 1010 205 1015
rect 70 965 205 1010
rect 255 965 275 1015
rect 70 960 275 965
rect 70 910 90 960
rect 140 915 275 960
rect 140 910 205 915
rect 70 865 205 910
rect 255 865 275 915
rect 70 855 275 865
rect 70 805 90 855
rect 140 815 275 855
rect 140 805 205 815
rect 70 765 205 805
rect 255 765 275 815
rect 70 760 275 765
rect 180 745 275 760
rect 375 1260 465 1280
rect 375 1210 395 1260
rect 445 1210 465 1260
rect 375 1080 465 1210
rect 375 1030 395 1080
rect 445 1030 465 1080
rect 375 980 465 1030
rect 375 930 395 980
rect 445 930 465 980
rect 375 845 465 930
rect 565 1260 655 1395
rect 565 1210 585 1260
rect 635 1210 655 1260
rect 565 1115 655 1210
rect 565 1065 585 1115
rect 635 1065 655 1115
rect 565 975 655 1065
rect 565 925 585 975
rect 635 925 655 975
rect 565 905 655 925
rect 755 1260 845 1280
rect 755 1210 775 1260
rect 825 1210 845 1260
rect 755 1085 845 1210
rect 755 1035 775 1085
rect 825 1035 845 1085
rect 755 985 845 1035
rect 755 935 775 985
rect 825 935 845 985
rect 755 885 845 935
rect 755 845 775 885
rect 375 835 775 845
rect 825 835 845 885
rect 375 825 845 835
rect 375 775 395 825
rect 445 785 845 825
rect 445 775 775 785
rect 375 755 775 775
rect 755 735 775 755
rect 825 735 845 785
rect 185 665 675 685
rect 185 615 205 665
rect 255 615 305 665
rect 355 615 405 665
rect 455 615 505 665
rect 555 615 605 665
rect 655 615 675 665
rect 185 595 675 615
rect 755 525 845 735
rect 375 435 845 525
rect 185 370 275 390
rect 185 340 205 370
rect 70 320 205 340
rect 255 320 275 370
rect 70 270 90 320
rect 140 270 275 320
rect 70 205 275 270
rect 70 155 90 205
rect 140 155 205 205
rect 255 155 275 205
rect 70 45 275 155
rect 375 370 465 435
rect 375 320 395 370
rect 445 320 465 370
rect 755 370 845 435
rect 375 205 465 320
rect 375 155 395 205
rect 445 155 465 205
rect 375 135 465 155
rect 565 345 655 365
rect 565 295 585 345
rect 635 295 655 345
rect 565 205 655 295
rect 565 155 585 205
rect 635 155 655 205
rect 565 45 655 155
rect 755 320 775 370
rect 825 320 845 370
rect 755 205 845 320
rect 755 155 775 205
rect 825 155 845 205
rect 755 135 845 155
rect 0 -45 900 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 3 ne
flabel metal1 s 20 1430 20 1430 2 FreeSans 400 0 0 0 vdd
port 2 ne
flabel nwell 170 555 170 555 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 205 605 205 605 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 405 470 405 470 2 FreeSans 400 0 0 0 z
port 0 ne
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
