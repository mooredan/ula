magic
tech amic5n
timestamp 1625182294
<< nwell >>
rect -130 550 880 1495
rect 105 150 645 550
<< polysilicon >>
rect 105 1240 645 1290
rect 105 1220 225 1240
rect 105 1170 125 1220
rect 175 1170 225 1220
rect 525 1220 645 1240
rect 105 1120 225 1170
rect 525 1170 575 1220
rect 625 1170 645 1220
rect 105 1070 125 1120
rect 175 1070 225 1120
rect 525 1120 645 1170
rect 525 1070 575 1120
rect 625 1070 645 1120
rect 105 1020 225 1070
rect 525 1020 645 1070
rect 105 970 125 1020
rect 175 970 225 1020
rect 105 920 225 970
rect 525 970 575 1020
rect 625 970 645 1020
rect 105 870 125 920
rect 175 870 225 920
rect 525 920 645 970
rect 105 820 225 870
rect 525 870 575 920
rect 625 870 645 920
rect 105 770 125 820
rect 175 770 225 820
rect 525 820 645 870
rect 105 720 225 770
rect 525 770 575 820
rect 625 770 645 820
rect 105 670 125 720
rect 175 670 225 720
rect 525 720 645 770
rect 105 620 225 670
rect 525 670 575 720
rect 625 670 645 720
rect 105 570 125 620
rect 175 570 225 620
rect 525 620 645 670
rect 105 520 225 570
rect 525 570 575 620
rect 625 570 645 620
rect 525 520 645 570
rect 105 470 125 520
rect 175 470 225 520
rect 525 470 575 520
rect 625 470 645 520
rect 105 420 225 470
rect 105 370 125 420
rect 175 370 225 420
rect 525 420 645 470
rect 105 320 225 370
rect 525 370 575 420
rect 625 370 645 420
rect 105 270 125 320
rect 175 270 225 320
rect 525 320 645 370
rect 105 220 225 270
rect 525 270 575 320
rect 625 270 645 320
rect 105 170 125 220
rect 175 200 225 220
rect 525 220 645 270
rect 525 200 575 220
rect 175 170 575 200
rect 625 170 645 220
rect 105 150 645 170
<< polycontact >>
rect 125 1170 175 1220
rect 575 1170 625 1220
rect 125 1070 175 1120
rect 575 1070 625 1120
rect 125 970 175 1020
rect 575 970 625 1020
rect 125 870 175 920
rect 575 870 625 920
rect 125 770 175 820
rect 575 770 625 820
rect 125 670 175 720
rect 575 670 625 720
rect 125 570 175 620
rect 575 570 625 620
rect 125 470 175 520
rect 575 470 625 520
rect 125 370 175 420
rect 575 370 625 420
rect 125 270 175 320
rect 575 270 625 320
rect 125 170 175 220
rect 575 170 625 220
<< poly2cap >>
rect 225 1180 525 1240
rect 225 1130 275 1180
rect 325 1130 425 1180
rect 475 1130 525 1180
rect 225 1070 525 1130
rect 225 1020 275 1070
rect 325 1020 425 1070
rect 475 1020 525 1070
rect 225 960 525 1020
rect 225 910 275 960
rect 325 910 425 960
rect 475 910 525 960
rect 225 850 525 910
rect 225 800 275 850
rect 325 800 425 850
rect 475 800 525 850
rect 225 740 525 800
rect 225 690 275 740
rect 325 690 425 740
rect 475 690 525 740
rect 225 630 525 690
rect 225 580 275 630
rect 325 580 425 630
rect 475 580 525 630
rect 225 520 525 580
rect 225 470 275 520
rect 325 470 425 520
rect 475 470 525 520
rect 225 410 525 470
rect 225 360 275 410
rect 325 360 425 410
rect 475 360 525 410
rect 225 300 525 360
rect 225 250 275 300
rect 325 250 425 300
rect 475 250 525 300
rect 225 200 525 250
<< poly2capcontact >>
rect 275 1130 325 1180
rect 425 1130 475 1180
rect 275 1020 325 1070
rect 425 1020 475 1070
rect 275 910 325 960
rect 425 910 475 960
rect 275 800 325 850
rect 425 800 475 850
rect 275 690 325 740
rect 425 690 475 740
rect 275 580 325 630
rect 425 580 475 630
rect 275 470 325 520
rect 425 470 475 520
rect 275 360 325 410
rect 425 360 475 410
rect 275 250 325 300
rect 425 250 475 300
<< metal1 >>
rect 0 1395 750 1485
rect 165 1305 585 1395
rect 105 1220 195 1240
rect 105 1170 125 1220
rect 175 1170 195 1220
rect 105 1120 195 1170
rect 105 1070 125 1120
rect 175 1070 195 1120
rect 105 1020 195 1070
rect 105 970 125 1020
rect 175 970 195 1020
rect 105 920 195 970
rect 105 870 125 920
rect 175 870 195 920
rect 105 820 195 870
rect 105 770 125 820
rect 175 770 195 820
rect 105 720 195 770
rect 105 670 125 720
rect 175 670 195 720
rect 105 620 195 670
rect 105 570 125 620
rect 175 570 195 620
rect 105 520 195 570
rect 105 470 125 520
rect 175 470 195 520
rect 105 420 195 470
rect 105 370 125 420
rect 175 370 195 420
rect 105 320 195 370
rect 105 270 125 320
rect 175 270 195 320
rect 105 220 195 270
rect 255 1180 495 1305
rect 255 1130 275 1180
rect 325 1130 425 1180
rect 475 1130 495 1180
rect 255 1070 495 1130
rect 255 1020 275 1070
rect 325 1020 425 1070
rect 475 1020 495 1070
rect 255 960 495 1020
rect 255 910 275 960
rect 325 910 425 960
rect 475 910 495 960
rect 255 850 495 910
rect 255 800 275 850
rect 325 800 425 850
rect 475 800 495 850
rect 255 740 495 800
rect 255 690 275 740
rect 325 690 425 740
rect 475 690 495 740
rect 255 630 495 690
rect 255 580 275 630
rect 325 580 425 630
rect 475 580 495 630
rect 255 520 495 580
rect 255 470 275 520
rect 325 470 425 520
rect 475 470 495 520
rect 255 410 495 470
rect 255 360 275 410
rect 325 360 425 410
rect 475 360 495 410
rect 255 300 495 360
rect 255 250 275 300
rect 325 250 425 300
rect 475 250 495 300
rect 255 230 495 250
rect 555 1220 645 1240
rect 555 1170 575 1220
rect 625 1170 645 1220
rect 555 1120 645 1170
rect 555 1070 575 1120
rect 625 1070 645 1120
rect 555 1020 645 1070
rect 555 970 575 1020
rect 625 970 645 1020
rect 555 920 645 970
rect 555 870 575 920
rect 625 870 645 920
rect 555 820 645 870
rect 555 770 575 820
rect 625 770 645 820
rect 555 720 645 770
rect 555 670 575 720
rect 625 670 645 720
rect 555 620 645 670
rect 555 570 575 620
rect 625 570 645 620
rect 555 520 645 570
rect 555 470 575 520
rect 625 470 645 520
rect 555 420 645 470
rect 555 370 575 420
rect 625 370 645 420
rect 555 320 645 370
rect 555 270 575 320
rect 625 270 645 320
rect 105 170 125 220
rect 175 170 195 220
rect 105 150 195 170
rect 555 220 645 270
rect 555 170 575 220
rect 625 170 645 220
rect 555 150 645 170
rect 105 45 645 150
rect 0 -45 750 45
<< labels >>
flabel metal1 s 95 1415 95 1415 2 FreeSans 400 0 0 0 vdd
port 0 ne
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 1 ne
flabel nwell 5 580 5 580 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFclass CORE
string LEFsite core
string FIXED_BBOX 0 0 750 1440
string LEFsymmetry X Y
<< end >>
