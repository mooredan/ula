magic
tech amic5n
timestamp 1621830667
use inv_c  inv_c_3
timestamp 1621808710
transform -1 0 -1505 0 1 -40
box -105 -45 495 2455
use inv_c  inv_c_2
timestamp 1621808710
transform 1 0 -1505 0 1 -40
box -105 -45 495 2455
use inv_c  inv_c_1
timestamp 1621808710
transform -1 0 -725 0 1 -40
box -105 -45 495 2455
use inv_c  inv_c_0
timestamp 1621808710
transform -1 0 -335 0 1 -40
box -105 -45 495 2455
use inv_c  inv_c_9
timestamp 1621808710
transform -1 0 -335 0 -1 -40
box -105 -45 495 2455
use inv_c  inv_c_8
timestamp 1621808710
transform -1 0 -725 0 -1 -40
box -105 -45 495 2455
use inv_c  inv_c_7
timestamp 1621808710
transform 1 0 -1505 0 -1 -40
box -105 -45 495 2455
use inv_c  inv_c_6
timestamp 1621808710
transform -1 0 -1505 0 -1 -40
box -105 -45 495 2455
use inv_c  inv_c_11
timestamp 1621808710
transform -1 0 -1505 0 -1 4760
box -105 -45 495 2455
use inv_c  inv_c_10
timestamp 1621808710
transform 1 0 -1505 0 -1 4760
box -105 -45 495 2455
use inv_c  inv_c_5
timestamp 1621808710
transform -1 0 -725 0 -1 4760
box -105 -45 495 2455
use inv_c  inv_c_4
timestamp 1621808710
transform -1 0 -335 0 -1 4760
box -105 -45 495 2455
<< end >>
