magic
tech amic5n
timestamp 1608317708
<< nwell >>
rect -120 870 600 2430
<< nselect >>
rect 0 60 480 750
<< pselect >>
rect 0 990 480 2310
<< ntransistor >>
rect 210 120 270 690
<< ptransistor >>
rect 210 1050 270 2250
<< ndiffusion >>
rect 60 120 210 690
rect 270 120 420 690
<< pdiffusion >>
rect 60 1050 210 2250
rect 270 1050 420 2250
<< polysilicon >>
rect 210 2250 270 2310
rect 210 960 270 1050
rect 60 780 270 960
rect 210 690 270 780
rect 210 60 270 120
<< pdcontact >>
rect 95 2165 145 2215
<< pdcontact >>
rect 335 2105 385 2155
<< pdcontact >>
rect 95 1985 145 2035
<< pdcontact >>
rect 335 1955 385 2005
<< pdcontact >>
rect 95 1835 145 1885
<< pdcontact >>
rect 335 1775 385 1825
<< pdcontact >>
rect 95 1685 145 1735
<< pdcontact >>
rect 335 1595 385 1645
<< pdcontact >>
rect 95 1535 145 1585
<< pdcontact >>
rect 95 1385 145 1435
<< pdcontact >>
rect 335 1415 385 1465
<< pdcontact >>
rect 95 1235 145 1285
<< pdcontact >>
rect 335 1235 385 1285
<< pdcontact >>
rect 95 1085 145 1135
<< pdcontact >>
rect 335 1085 385 1135
<< polycontact >>
rect 125 845 175 895
<< ndcontact >>
rect 95 605 145 655
<< ndcontact >>
rect 335 605 385 655
<< ndcontact >>
rect 95 455 145 505
<< ndcontact >>
rect 335 395 385 445
<< ndcontact >>
rect 95 305 145 355
<< ndcontact >>
rect 335 215 385 265
<< ndcontact >>
rect 95 155 145 205
<< metal1 >>
rect 0 2280 480 2370
rect 60 1050 180 2280
rect 300 1050 420 2190
rect 90 810 420 930
rect 60 90 180 690
rect 300 180 420 810
rect 0 0 480 90
<< labels >>
flabel metal1 s 30 30 30 30 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 30 2310 30 2310 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel nwell  0 930 0 930 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 360 1170 360 1170 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 330 810 330 810 2 FreeSans 400 0 0 0 n1
<< checkpaint >>
rect -130 -10 610 2440
<< end >>
