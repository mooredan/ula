`celldefine
module decap6 ();
endmodule
`endcelldefine
