magic
tech scmos
timestamp 1606579561
<< nwell >>
rect -14 -3 22 24
<< ntransistor >>
rect 7 -29 9 -12
<< ptransistor >>
rect 7 3 9 18
<< ndiffusion >>
rect 3 -29 7 -12
rect 9 -29 13 -12
<< pdiffusion >>
rect 5 12 7 18
rect -1 9 7 12
rect 5 3 7 9
rect 9 3 16 18
<< pdcontact >>
rect -1 12 5 18
rect -1 3 5 9
<< nsubstratendiff >>
rect -8 9 -1 11
rect -2 3 -1 9
<< nsubstratencontact >>
rect -8 3 -2 9
<< polysilicon >>
rect 7 18 9 20
rect 7 -12 9 3
rect 7 -31 9 -29
<< metal1 >>
rect -2 3 -1 9
<< end >>
