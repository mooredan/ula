magic
tech scmos
timestamp 1591495604
<< nwell >>
rect -1 29 57 81
<< nselect >>
rect 15 2 29 25
<< pselect >>
rect 12 33 40 77
<< ntransistor >>
rect 21 4 23 23
<< ptransistor >>
rect 20 35 22 75
rect 29 35 31 75
<< ndiffusion >>
rect 17 4 21 23
rect 23 4 27 23
<< pdiffusion >>
rect 14 35 20 75
rect 22 35 29 75
rect 31 35 38 75
<< polysilicon >>
rect 20 75 22 77
rect 29 75 31 77
rect 20 33 22 35
rect 29 33 31 35
rect 21 23 23 30
rect 21 2 23 4
<< metal1 >>
rect 5 76 51 79
rect 6 69 16 73
rect 40 69 50 73
rect 6 62 17 66
rect 40 62 50 66
rect 6 55 17 59
rect 40 55 50 59
rect 6 48 17 52
rect 40 48 50 52
rect 6 41 17 45
rect 40 41 50 45
rect 6 34 17 38
rect 40 34 50 38
rect 6 27 17 31
rect 40 27 50 31
rect 6 20 15 24
rect 39 20 50 24
rect 6 13 15 17
rect 39 13 50 17
rect 6 6 15 10
rect 39 6 50 10
rect 5 0 51 3
rect -2 -10 2 -3
rect 5 -10 9 -3
rect 12 -10 16 -3
rect 19 -10 23 -3
rect 26 -10 30 -3
rect 33 -10 37 -3
rect 40 -10 44 -3
rect 47 -10 51 -3
rect 54 -10 58 -3
<< bb >>
rect 0 0 56 79
<< labels >>
rlabel metal1 5 0 5 0 2 Gnd
port 3 ne
rlabel nwell 5 30 5 30 2 Vdd
rlabel metal1 5 76 5 76 2 Vdd
port 2 ne
<< end >>
