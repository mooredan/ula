magic
tech amic5n
timestamp 1608397441
<< metal1 >>
rect 900 2100 1470 2190
rect 960 -180 4470 -90
<< metal2 >>
rect 840 630 1950 750
<< via1 >>
rect 875 665 925 715
use inv_e  inv_e_1
transform 1 0 55 0 1 -6
box -120 0 1320 2430
use inv_e  inv_e_0
transform 1 0 -6 0 1 -6
box -120 0 1320 2430
use subc_2  subc_2_0
transform 1 0 38 0 1 -6
box -30 0 450 2430
<< labels >>
flabel metal1 s 1110 -150 1110 -150 2 FreeSans 400 0 0 0 vss
flabel metal1 s 1170 2130 1170 2130 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 2400 -150 2400 -150 2 FreeSans 400 0 0 0 vss
flabel metal1 s 2490 900 2490 900 2 FreeSans 400 0 0 0 z1
flabel metal2 s 2340 660 2340 660 2 FreeSans 400 0 0 0 n1
flabel metal2 s 330 660 330 660 2 FreeSans 400 0 0 0 a2
<< checkpaint >>
rect -10 -190 4480 2200
<< end >>
