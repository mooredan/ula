magic
tech scmos
timestamp 1591575340
use newsub  newsub_0 mag
timestamp 1591575201
transform 1 0 32 0 1 0
box -1 0 15 81
use inv_c  inv_c_0 mag
timestamp 1591570911
transform 1 0 0 0 1 0
box -4 0 20 81
<< end >>
