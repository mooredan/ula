magic
tech scmos
timestamp 1591543887
<< error_s >>
rect 42 76 44 79
rect 42 0 44 6
use newsub  newsub_0
timestamp 1591542839
transform 1 0 37 0 1 0
box -1 0 15 81
use inv_c  inv_c_1 ~/projects/ula/mag
timestamp 1591543887
transform 1 0 18 0 1 0
box -1 0 29 81
use inv_c  inv_c_0
timestamp 1591543887
transform 1 0 0 0 1 0
box -1 0 29 81
<< end >>
