magic
tech scmos
timestamp 1591539261
<< nwell >>
rect -1 29 36 81
<< nselect >>
rect 15 2 29 25
<< pselect >>
rect 12 33 29 77
<< ntransistor >>
rect 21 4 23 23
<< ptransistor >>
rect 20 35 22 75
<< ndiffusion >>
rect 17 4 21 23
rect 23 4 27 23
<< pdiffusion >>
rect 14 35 20 75
rect 22 35 27 75
<< polysilicon >>
rect 20 75 22 77
rect 20 33 22 35
rect 21 23 23 30
rect 21 2 23 4
<< metal1 >>
rect 5 76 30 79
rect 6 69 9 73
rect 26 69 29 73
rect 6 62 9 66
rect 26 62 29 66
rect 6 55 9 59
rect 26 55 29 59
rect 6 48 9 52
rect 26 48 29 52
rect 6 41 9 45
rect 26 41 29 45
rect 6 34 9 38
rect 26 34 29 38
rect 6 27 9 31
rect 26 27 29 31
rect 6 20 9 24
rect 26 20 29 24
rect 6 13 9 17
rect 26 13 29 17
rect 6 6 9 10
rect 26 6 29 10
rect 5 0 30 3
rect -2 -10 2 -3
rect 5 -10 9 -3
rect 12 -10 16 -3
rect 19 -10 23 -3
rect 26 -10 30 -3
rect 33 -10 37 -3
<< bb >>
rect 0 0 35 79
<< labels >>
rlabel metal1 5 0 5 0 2 Gnd
port 3 ne
rlabel nwell 5 30 5 30 2 Vdd
rlabel metal1 5 76 5 76 2 Vdd
port 2 ne
<< end >>
