magic
tech amic5n
timestamp 1624412454
<< nwell >>
rect -130 550 2830 1495
<< ntransistor >>
rect 295 125 355 400
rect 485 125 545 400
rect 675 125 735 400
rect 1075 115 1135 400
rect 1265 115 1325 400
rect 1455 115 1515 400
rect 1645 115 1705 400
rect 1835 115 1895 400
rect 2025 115 2085 400
rect 2215 115 2275 400
rect 2405 115 2465 400
<< ptransistor >>
rect 295 705 355 1290
rect 485 705 545 1290
rect 675 705 735 1290
rect 1075 705 1135 1300
rect 1265 705 1325 1300
rect 1455 705 1515 1300
rect 1645 705 1705 1300
rect 1835 705 1895 1300
rect 2025 705 2085 1300
rect 2215 705 2275 1300
rect 2405 705 2465 1300
<< nselect >>
rect 10 765 175 1290
rect -10 350 2710 430
rect 175 125 2710 350
rect -10 0 2710 125
<< pselect >>
rect -10 1290 2710 1440
rect 175 765 2710 1290
rect -10 670 2710 765
rect 10 125 175 350
<< ndiffusion >>
rect 175 370 295 400
rect 175 320 205 370
rect 255 320 295 370
rect 175 205 295 320
rect 175 155 205 205
rect 255 155 295 205
rect 175 125 295 155
rect 355 370 485 400
rect 355 320 395 370
rect 445 320 485 370
rect 355 205 485 320
rect 355 155 395 205
rect 445 155 485 205
rect 355 125 485 155
rect 545 345 675 400
rect 545 295 585 345
rect 635 295 675 345
rect 545 205 675 295
rect 545 155 585 205
rect 635 155 675 205
rect 545 125 675 155
rect 735 370 855 400
rect 735 320 775 370
rect 825 320 855 370
rect 735 205 855 320
rect 735 155 775 205
rect 825 155 855 205
rect 735 125 855 155
rect 955 355 1075 400
rect 955 305 985 355
rect 1035 305 1075 355
rect 955 205 1075 305
rect 955 155 985 205
rect 1035 155 1075 205
rect 955 115 1075 155
rect 1135 370 1265 400
rect 1135 320 1175 370
rect 1225 320 1265 370
rect 1135 205 1265 320
rect 1135 155 1175 205
rect 1225 155 1265 205
rect 1135 115 1265 155
rect 1325 345 1455 400
rect 1325 295 1365 345
rect 1415 295 1455 345
rect 1325 205 1455 295
rect 1325 155 1365 205
rect 1415 155 1455 205
rect 1325 115 1455 155
rect 1515 370 1645 400
rect 1515 320 1555 370
rect 1605 320 1645 370
rect 1515 205 1645 320
rect 1515 155 1555 205
rect 1605 155 1645 205
rect 1515 115 1645 155
rect 1705 345 1835 400
rect 1705 295 1745 345
rect 1795 295 1835 345
rect 1705 205 1835 295
rect 1705 155 1745 205
rect 1795 155 1835 205
rect 1705 115 1835 155
rect 1895 370 2025 400
rect 1895 320 1935 370
rect 1985 320 2025 370
rect 1895 205 2025 320
rect 1895 155 1935 205
rect 1985 155 2025 205
rect 1895 115 2025 155
rect 2085 355 2215 400
rect 2085 305 2125 355
rect 2175 305 2215 355
rect 2085 205 2215 305
rect 2085 155 2125 205
rect 2175 155 2215 205
rect 2085 115 2215 155
rect 2275 370 2405 400
rect 2275 320 2315 370
rect 2365 320 2405 370
rect 2275 205 2405 320
rect 2275 155 2315 205
rect 2365 155 2405 205
rect 2275 115 2405 155
rect 2465 345 2595 400
rect 2465 295 2505 345
rect 2555 295 2595 345
rect 2465 205 2595 295
rect 2465 155 2505 205
rect 2555 155 2595 205
rect 2465 115 2595 155
<< pdiffusion >>
rect 175 1260 295 1290
rect 175 1210 205 1260
rect 255 1210 295 1260
rect 175 1115 295 1210
rect 175 1065 205 1115
rect 255 1065 295 1115
rect 175 1015 295 1065
rect 175 965 205 1015
rect 255 965 295 1015
rect 175 915 295 965
rect 175 865 205 915
rect 255 865 295 915
rect 175 815 295 865
rect 175 765 205 815
rect 255 765 295 815
rect 175 705 295 765
rect 355 1260 485 1290
rect 355 1210 395 1260
rect 445 1210 485 1260
rect 355 1080 485 1210
rect 355 1030 395 1080
rect 445 1030 485 1080
rect 355 980 485 1030
rect 355 930 395 980
rect 445 930 485 980
rect 355 825 485 930
rect 355 775 395 825
rect 445 775 485 825
rect 355 705 485 775
rect 545 1260 675 1290
rect 545 1210 585 1260
rect 635 1210 675 1260
rect 545 1115 675 1210
rect 545 1065 585 1115
rect 635 1065 675 1115
rect 545 975 675 1065
rect 545 925 585 975
rect 635 925 675 975
rect 545 705 675 925
rect 735 1260 855 1290
rect 735 1210 775 1260
rect 825 1210 855 1260
rect 735 1085 855 1210
rect 735 1035 775 1085
rect 825 1035 855 1085
rect 735 985 855 1035
rect 735 935 775 985
rect 825 935 855 985
rect 735 885 855 935
rect 735 835 775 885
rect 825 835 855 885
rect 735 785 855 835
rect 735 735 775 785
rect 825 735 855 785
rect 735 705 855 735
rect 955 1260 1075 1300
rect 955 1210 985 1260
rect 1035 1210 1075 1260
rect 955 1115 1075 1210
rect 955 1065 985 1115
rect 1035 1065 1075 1115
rect 955 1015 1075 1065
rect 955 965 985 1015
rect 1035 965 1075 1015
rect 955 915 1075 965
rect 955 865 985 915
rect 1035 865 1075 915
rect 955 815 1075 865
rect 955 765 985 815
rect 1035 765 1075 815
rect 955 705 1075 765
rect 1135 1260 1265 1300
rect 1135 1210 1175 1260
rect 1225 1210 1265 1260
rect 1135 1080 1265 1210
rect 1135 1030 1175 1080
rect 1225 1030 1265 1080
rect 1135 980 1265 1030
rect 1135 930 1175 980
rect 1225 930 1265 980
rect 1135 825 1265 930
rect 1135 775 1175 825
rect 1225 775 1265 825
rect 1135 705 1265 775
rect 1325 1260 1455 1300
rect 1325 1210 1365 1260
rect 1415 1210 1455 1260
rect 1325 1115 1455 1210
rect 1325 1065 1365 1115
rect 1415 1065 1455 1115
rect 1325 975 1455 1065
rect 1325 925 1365 975
rect 1415 925 1455 975
rect 1325 705 1455 925
rect 1515 1260 1645 1300
rect 1515 1210 1555 1260
rect 1605 1210 1645 1260
rect 1515 1080 1645 1210
rect 1515 1030 1555 1080
rect 1605 1030 1645 1080
rect 1515 980 1645 1030
rect 1515 930 1555 980
rect 1605 930 1645 980
rect 1515 825 1645 930
rect 1515 775 1555 825
rect 1605 775 1645 825
rect 1515 705 1645 775
rect 1705 1260 1835 1300
rect 1705 1210 1745 1260
rect 1795 1210 1835 1260
rect 1705 1115 1835 1210
rect 1705 1065 1745 1115
rect 1795 1065 1835 1115
rect 1705 975 1835 1065
rect 1705 925 1745 975
rect 1795 925 1835 975
rect 1705 705 1835 925
rect 1895 1260 2025 1300
rect 1895 1210 1935 1260
rect 1985 1210 2025 1260
rect 1895 1080 2025 1210
rect 1895 1030 1935 1080
rect 1985 1030 2025 1080
rect 1895 980 2025 1030
rect 1895 930 1935 980
rect 1985 930 2025 980
rect 1895 825 2025 930
rect 1895 775 1935 825
rect 1985 775 2025 825
rect 1895 705 2025 775
rect 2085 1260 2215 1300
rect 2085 1210 2125 1260
rect 2175 1210 2215 1260
rect 2085 1115 2215 1210
rect 2085 1065 2125 1115
rect 2175 1065 2215 1115
rect 2085 975 2215 1065
rect 2085 925 2125 975
rect 2175 925 2215 975
rect 2085 705 2215 925
rect 2275 1260 2405 1300
rect 2275 1210 2315 1260
rect 2365 1210 2405 1260
rect 2275 1080 2405 1210
rect 2275 1030 2315 1080
rect 2365 1030 2405 1080
rect 2275 980 2405 1030
rect 2275 930 2315 980
rect 2365 930 2405 980
rect 2275 825 2405 930
rect 2275 775 2315 825
rect 2365 775 2405 825
rect 2275 705 2405 775
rect 2465 1260 2595 1300
rect 2465 1210 2505 1260
rect 2555 1210 2595 1260
rect 2465 1115 2595 1210
rect 2465 1065 2505 1115
rect 2555 1065 2595 1115
rect 2465 975 2595 1065
rect 2465 925 2505 975
rect 2555 925 2595 975
rect 2465 705 2595 925
<< psubstratepdiff >>
rect 60 320 175 350
rect 60 270 90 320
rect 140 270 175 320
rect 60 205 175 270
rect 60 155 90 205
rect 140 155 175 205
rect 60 125 175 155
<< nsubstratendiff >>
rect 60 1260 175 1290
rect 60 1210 95 1260
rect 145 1210 175 1260
rect 60 1160 175 1210
rect 60 1110 90 1160
rect 140 1110 175 1160
rect 60 1060 175 1110
rect 60 1010 90 1060
rect 140 1010 175 1060
rect 60 960 175 1010
rect 60 910 90 960
rect 140 910 175 960
rect 60 855 175 910
rect 60 805 90 855
rect 140 805 175 855
rect 60 765 175 805
<< nsubstratencontact >>
rect 95 1210 145 1260
rect 90 1110 140 1160
rect 90 1010 140 1060
rect 90 910 140 960
rect 90 805 140 855
<< psubstratepcontact >>
rect 90 270 140 320
rect 90 155 140 205
<< ndcontact >>
rect 205 320 255 370
rect 205 155 255 205
rect 395 320 445 370
rect 395 155 445 205
rect 585 295 635 345
rect 585 155 635 205
rect 775 320 825 370
rect 775 155 825 205
rect 985 305 1035 355
rect 985 155 1035 205
rect 1175 320 1225 370
rect 1175 155 1225 205
rect 1365 295 1415 345
rect 1365 155 1415 205
rect 1555 320 1605 370
rect 1555 155 1605 205
rect 1745 295 1795 345
rect 1745 155 1795 205
rect 1935 320 1985 370
rect 1935 155 1985 205
rect 2125 305 2175 355
rect 2125 155 2175 205
rect 2315 320 2365 370
rect 2315 155 2365 205
rect 2505 295 2555 345
rect 2505 155 2555 205
<< pdcontact >>
rect 205 1210 255 1260
rect 205 1065 255 1115
rect 205 965 255 1015
rect 205 865 255 915
rect 205 765 255 815
rect 395 1210 445 1260
rect 395 1030 445 1080
rect 395 930 445 980
rect 395 775 445 825
rect 585 1210 635 1260
rect 585 1065 635 1115
rect 585 925 635 975
rect 775 1210 825 1260
rect 775 1035 825 1085
rect 775 935 825 985
rect 775 835 825 885
rect 775 735 825 785
rect 985 1210 1035 1260
rect 985 1065 1035 1115
rect 985 965 1035 1015
rect 985 865 1035 915
rect 985 765 1035 815
rect 1175 1210 1225 1260
rect 1175 1030 1225 1080
rect 1175 930 1225 980
rect 1175 775 1225 825
rect 1365 1210 1415 1260
rect 1365 1065 1415 1115
rect 1365 925 1415 975
rect 1555 1210 1605 1260
rect 1555 1030 1605 1080
rect 1555 930 1605 980
rect 1555 775 1605 825
rect 1745 1210 1795 1260
rect 1745 1065 1795 1115
rect 1745 925 1795 975
rect 1935 1210 1985 1260
rect 1935 1030 1985 1080
rect 1935 930 1985 980
rect 1935 775 1985 825
rect 2125 1210 2175 1260
rect 2125 1065 2175 1115
rect 2125 925 2175 975
rect 2315 1210 2365 1260
rect 2315 1030 2365 1080
rect 2315 930 2365 980
rect 2315 775 2365 825
rect 2505 1210 2555 1260
rect 2505 1065 2555 1115
rect 2505 925 2555 975
<< polysilicon >>
rect 295 1290 355 1355
rect 485 1290 545 1355
rect 675 1290 735 1355
rect 1075 1300 1135 1365
rect 1265 1300 1325 1365
rect 1455 1300 1515 1365
rect 1645 1300 1705 1365
rect 1835 1300 1895 1365
rect 2025 1300 2085 1365
rect 2215 1300 2275 1365
rect 2405 1300 2465 1365
rect 295 685 355 705
rect 485 685 545 705
rect 675 685 735 705
rect 1075 685 1135 705
rect 1265 685 1325 705
rect 1455 685 1515 705
rect 1645 685 1705 705
rect 1835 685 1895 705
rect 2025 685 2085 705
rect 2215 685 2275 705
rect 2405 685 2465 705
rect 185 665 735 685
rect 185 615 205 665
rect 255 615 305 665
rect 355 615 405 665
rect 455 615 505 665
rect 555 615 605 665
rect 655 615 735 665
rect 185 595 735 615
rect 965 665 2465 685
rect 965 615 985 665
rect 1035 615 1085 665
rect 1135 615 1185 665
rect 1235 615 1285 665
rect 1335 615 1385 665
rect 1435 615 1485 665
rect 1535 615 1585 665
rect 1635 615 1725 665
rect 1775 615 1825 665
rect 1875 615 1925 665
rect 1975 615 2025 665
rect 2075 615 2125 665
rect 2175 615 2225 665
rect 2275 615 2325 665
rect 2375 615 2465 665
rect 965 595 2465 615
rect 295 400 355 595
rect 485 400 545 595
rect 675 400 735 595
rect 1075 400 1135 595
rect 1265 400 1325 595
rect 1455 400 1515 595
rect 1645 400 1705 595
rect 1835 400 1895 595
rect 2025 400 2085 595
rect 2215 400 2275 595
rect 2405 400 2465 595
rect 295 60 355 125
rect 485 60 545 125
rect 675 60 735 125
rect 1075 50 1135 115
rect 1265 50 1325 115
rect 1455 50 1515 115
rect 1645 50 1705 115
rect 1835 50 1895 115
rect 2025 50 2085 115
rect 2215 50 2275 115
rect 2405 50 2465 115
<< polycontact >>
rect 205 615 255 665
rect 305 615 355 665
rect 405 615 455 665
rect 505 615 555 665
rect 605 615 655 665
rect 985 615 1035 665
rect 1085 615 1135 665
rect 1185 615 1235 665
rect 1285 615 1335 665
rect 1385 615 1435 665
rect 1485 615 1535 665
rect 1585 615 1635 665
rect 1725 615 1775 665
rect 1825 615 1875 665
rect 1925 615 1975 665
rect 2025 615 2075 665
rect 2125 615 2175 665
rect 2225 615 2275 665
rect 2325 615 2375 665
<< metal1 >>
rect 0 1395 2700 1485
rect 70 1260 275 1395
rect 70 1210 95 1260
rect 145 1210 205 1260
rect 255 1210 275 1260
rect 70 1160 275 1210
rect 70 1110 90 1160
rect 140 1115 275 1160
rect 140 1110 205 1115
rect 70 1065 205 1110
rect 255 1065 275 1115
rect 70 1060 275 1065
rect 70 1010 90 1060
rect 140 1015 275 1060
rect 140 1010 205 1015
rect 70 965 205 1010
rect 255 965 275 1015
rect 70 960 275 965
rect 70 910 90 960
rect 140 915 275 960
rect 140 910 205 915
rect 70 865 205 910
rect 255 865 275 915
rect 70 855 275 865
rect 70 805 90 855
rect 140 815 275 855
rect 140 805 205 815
rect 70 765 205 805
rect 255 765 275 815
rect 70 760 275 765
rect 180 745 275 760
rect 375 1260 465 1280
rect 375 1210 395 1260
rect 445 1210 465 1260
rect 375 1080 465 1210
rect 375 1030 395 1080
rect 445 1030 465 1080
rect 375 980 465 1030
rect 375 930 395 980
rect 445 930 465 980
rect 375 845 465 930
rect 565 1260 655 1395
rect 565 1210 585 1260
rect 635 1210 655 1260
rect 565 1115 655 1210
rect 565 1065 585 1115
rect 635 1065 655 1115
rect 565 975 655 1065
rect 565 925 585 975
rect 635 925 655 975
rect 565 905 655 925
rect 755 1260 845 1280
rect 755 1210 775 1260
rect 825 1210 845 1260
rect 755 1085 845 1210
rect 755 1035 775 1085
rect 825 1035 845 1085
rect 755 985 845 1035
rect 755 935 775 985
rect 825 935 845 985
rect 755 885 845 935
rect 755 845 775 885
rect 375 835 775 845
rect 825 835 845 885
rect 375 825 845 835
rect 375 775 395 825
rect 445 785 845 825
rect 445 775 775 785
rect 375 755 775 775
rect 755 735 775 755
rect 825 735 845 785
rect 965 1260 1055 1395
rect 965 1210 985 1260
rect 1035 1210 1055 1260
rect 965 1115 1055 1210
rect 965 1065 985 1115
rect 1035 1065 1055 1115
rect 965 1015 1055 1065
rect 965 965 985 1015
rect 1035 965 1055 1015
rect 965 915 1055 965
rect 965 865 985 915
rect 1035 865 1055 915
rect 965 815 1055 865
rect 965 765 985 815
rect 1035 765 1055 815
rect 965 745 1055 765
rect 1155 1260 1245 1290
rect 1155 1210 1175 1260
rect 1225 1210 1245 1260
rect 1155 1080 1245 1210
rect 1155 1030 1175 1080
rect 1225 1030 1245 1080
rect 1155 980 1245 1030
rect 1155 930 1175 980
rect 1225 930 1245 980
rect 1155 845 1245 930
rect 1345 1260 1435 1395
rect 1345 1210 1365 1260
rect 1415 1210 1435 1260
rect 1345 1115 1435 1210
rect 1345 1065 1365 1115
rect 1415 1065 1435 1115
rect 1345 975 1435 1065
rect 1345 925 1365 975
rect 1415 925 1435 975
rect 1345 905 1435 925
rect 1535 1260 1625 1290
rect 1535 1210 1555 1260
rect 1605 1210 1625 1260
rect 1535 1080 1625 1210
rect 1535 1030 1555 1080
rect 1605 1030 1625 1080
rect 1535 980 1625 1030
rect 1535 930 1555 980
rect 1605 930 1625 980
rect 1535 845 1625 930
rect 1725 1260 1815 1395
rect 1725 1210 1745 1260
rect 1795 1210 1815 1260
rect 1725 1115 1815 1210
rect 1725 1065 1745 1115
rect 1795 1065 1815 1115
rect 1725 975 1815 1065
rect 1725 925 1745 975
rect 1795 925 1815 975
rect 1725 905 1815 925
rect 1915 1260 2005 1290
rect 1915 1210 1935 1260
rect 1985 1210 2005 1260
rect 1915 1080 2005 1210
rect 1915 1030 1935 1080
rect 1985 1030 2005 1080
rect 1915 980 2005 1030
rect 1915 930 1935 980
rect 1985 930 2005 980
rect 1915 845 2005 930
rect 2105 1260 2195 1395
rect 2105 1210 2125 1260
rect 2175 1210 2195 1260
rect 2105 1115 2195 1210
rect 2105 1065 2125 1115
rect 2175 1065 2195 1115
rect 2105 975 2195 1065
rect 2105 925 2125 975
rect 2175 925 2195 975
rect 2105 905 2195 925
rect 2295 1260 2385 1290
rect 2295 1210 2315 1260
rect 2365 1210 2385 1260
rect 2295 1080 2385 1210
rect 2295 1030 2315 1080
rect 2365 1030 2385 1080
rect 2295 980 2385 1030
rect 2295 930 2315 980
rect 2365 930 2385 980
rect 2295 845 2385 930
rect 2485 1260 2575 1395
rect 2485 1210 2505 1260
rect 2555 1210 2575 1260
rect 2485 1115 2575 1210
rect 2485 1065 2505 1115
rect 2555 1065 2575 1115
rect 2485 975 2575 1065
rect 2485 925 2505 975
rect 2555 925 2575 975
rect 2485 905 2575 925
rect 1155 825 2575 845
rect 1155 775 1175 825
rect 1225 775 1555 825
rect 1605 775 1935 825
rect 1985 775 2315 825
rect 2365 775 2575 825
rect 1155 755 2575 775
rect 755 685 845 735
rect 185 665 675 685
rect 185 615 205 665
rect 255 615 305 665
rect 355 615 405 665
rect 455 615 505 665
rect 555 615 605 665
rect 655 615 675 665
rect 185 595 675 615
rect 755 665 2405 685
rect 755 615 985 665
rect 1035 615 1085 665
rect 1135 615 1185 665
rect 1235 615 1285 665
rect 1335 615 1385 665
rect 1435 615 1485 665
rect 1535 615 1585 665
rect 1635 615 1725 665
rect 1775 615 1825 665
rect 1875 615 1925 665
rect 1975 615 2025 665
rect 2075 615 2125 665
rect 2175 615 2225 665
rect 2275 615 2325 665
rect 2375 615 2405 665
rect 755 595 2405 615
rect 755 525 1055 595
rect 2485 525 2575 755
rect 375 435 1055 525
rect 1155 435 2575 525
rect 185 370 275 390
rect 185 340 205 370
rect 70 320 205 340
rect 255 320 275 370
rect 70 270 90 320
rect 140 270 275 320
rect 70 205 275 270
rect 70 155 90 205
rect 140 155 205 205
rect 255 155 275 205
rect 70 45 275 155
rect 375 370 465 435
rect 375 320 395 370
rect 445 320 465 370
rect 755 370 845 435
rect 375 205 465 320
rect 375 155 395 205
rect 445 155 465 205
rect 375 135 465 155
rect 565 345 655 365
rect 565 295 585 345
rect 635 295 655 345
rect 565 205 655 295
rect 565 155 585 205
rect 635 155 655 205
rect 565 45 655 155
rect 755 320 775 370
rect 825 320 845 370
rect 755 205 845 320
rect 755 155 775 205
rect 825 155 845 205
rect 755 135 845 155
rect 965 355 1055 375
rect 965 305 985 355
rect 1035 305 1055 355
rect 965 205 1055 305
rect 965 155 985 205
rect 1035 155 1055 205
rect 965 45 1055 155
rect 1155 370 1245 435
rect 1155 320 1175 370
rect 1225 320 1245 370
rect 1535 370 1625 435
rect 1155 205 1245 320
rect 1155 155 1175 205
rect 1225 155 1245 205
rect 1155 125 1245 155
rect 1345 345 1435 365
rect 1345 295 1365 345
rect 1415 295 1435 345
rect 1345 205 1435 295
rect 1345 155 1365 205
rect 1415 155 1435 205
rect 1345 45 1435 155
rect 1535 320 1555 370
rect 1605 320 1625 370
rect 1915 370 2005 435
rect 1535 205 1625 320
rect 1535 155 1555 205
rect 1605 155 1625 205
rect 1535 125 1625 155
rect 1725 345 1815 365
rect 1725 295 1745 345
rect 1795 295 1815 345
rect 1725 205 1815 295
rect 1725 155 1745 205
rect 1795 155 1815 205
rect 1725 45 1815 155
rect 1915 320 1935 370
rect 1985 320 2005 370
rect 1915 205 2005 320
rect 1915 155 1935 205
rect 1985 155 2005 205
rect 1915 125 2005 155
rect 2105 355 2195 375
rect 2105 305 2125 355
rect 2175 305 2195 355
rect 2105 205 2195 305
rect 2105 155 2125 205
rect 2175 155 2195 205
rect 2105 45 2195 155
rect 2295 370 2385 435
rect 2295 320 2315 370
rect 2365 320 2385 370
rect 2295 205 2385 320
rect 2295 155 2315 205
rect 2365 155 2385 205
rect 2295 125 2385 155
rect 2485 345 2575 365
rect 2485 295 2505 345
rect 2555 295 2575 345
rect 2485 205 2575 295
rect 2485 155 2505 205
rect 2555 155 2575 205
rect 2485 45 2575 155
rect 0 -45 2700 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 3 ne
flabel metal1 s 20 1430 20 1430 2 FreeSans 400 0 0 0 vdd
port 2 ne
flabel nwell 170 555 170 555 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 205 605 205 605 2 FreeSans 400 0 0 0 a
port 1 ne
flabel metal1 s 1185 470 1185 470 2 FreeSans 400 0 0 0 z
port 0 ne
<< properties >>
string LEFsite core
string LEFclass CORE
string LEFsymmetry X Y
<< end >>
