magic
tech amic5n
timestamp 1607374361
<< nwell >>
rect -120 1470 3180 2430
rect -120 870 600 1470
rect 2460 870 3180 1470
<< ntransistor >>
rect 210 390 270 690
rect 2790 120 2850 690
<< ptransistor >>
rect 210 1050 270 1620
rect 2790 1050 2850 2250
<< nselect >>
rect 120 1710 360 2220
rect 0 300 480 750
rect 0 60 120 300
rect 360 60 480 300
rect 2580 60 3060 750
<< pselect >>
rect 0 2220 480 2310
rect 0 1710 120 2220
rect 360 1710 480 2220
rect 0 990 480 1710
rect 2580 990 3060 2310
rect 120 60 360 300
<< ndiffusion >>
rect 60 655 210 690
rect 60 605 95 655
rect 145 605 210 655
rect 60 505 210 605
rect 60 455 95 505
rect 145 455 210 505
rect 60 390 210 455
rect 270 655 420 690
rect 270 605 335 655
rect 385 605 420 655
rect 270 505 420 605
rect 270 455 335 505
rect 385 455 420 505
rect 270 390 420 455
rect 2640 655 2790 690
rect 2640 605 2675 655
rect 2725 605 2790 655
rect 2640 505 2790 605
rect 2640 455 2675 505
rect 2725 455 2790 505
rect 2640 355 2790 455
rect 2640 305 2675 355
rect 2725 305 2790 355
rect 2640 205 2790 305
rect 2640 155 2675 205
rect 2725 155 2790 205
rect 2640 120 2790 155
rect 2850 655 3000 690
rect 2850 605 2915 655
rect 2965 605 3000 655
rect 2850 445 3000 605
rect 2850 395 2915 445
rect 2965 395 3000 445
rect 2850 265 3000 395
rect 2850 215 2915 265
rect 2965 215 3000 265
rect 2850 120 3000 215
<< pdiffusion >>
rect 60 1525 210 1620
rect 60 1475 95 1525
rect 145 1475 210 1525
rect 60 1315 210 1475
rect 60 1265 95 1315
rect 145 1265 210 1315
rect 60 1135 210 1265
rect 60 1085 95 1135
rect 145 1085 210 1135
rect 60 1050 210 1085
rect 270 1525 420 1620
rect 270 1475 335 1525
rect 385 1475 420 1525
rect 2640 2215 2790 2250
rect 2640 2165 2675 2215
rect 2725 2165 2790 2215
rect 2640 2035 2790 2165
rect 2640 1985 2675 2035
rect 2725 1985 2790 2035
rect 2640 1885 2790 1985
rect 2640 1835 2675 1885
rect 2725 1835 2790 1885
rect 2640 1735 2790 1835
rect 2640 1685 2675 1735
rect 2725 1685 2790 1735
rect 2640 1585 2790 1685
rect 2640 1535 2675 1585
rect 2725 1535 2790 1585
rect 270 1315 420 1475
rect 2640 1435 2790 1535
rect 2640 1385 2675 1435
rect 2725 1385 2790 1435
rect 270 1265 335 1315
rect 385 1265 420 1315
rect 270 1135 420 1265
rect 2640 1285 2790 1385
rect 2640 1235 2675 1285
rect 2725 1235 2790 1285
rect 270 1085 335 1135
rect 385 1085 420 1135
rect 270 1050 420 1085
rect 2640 1050 2790 1235
rect 2850 2155 3000 2250
rect 2850 2105 2915 2155
rect 2965 2105 3000 2155
rect 2850 2005 3000 2105
rect 2850 1955 2915 2005
rect 2965 1955 3000 2005
rect 2850 1825 3000 1955
rect 2850 1775 2915 1825
rect 2965 1775 3000 1825
rect 2850 1645 3000 1775
rect 2850 1595 2915 1645
rect 2965 1595 3000 1645
rect 2850 1465 3000 1595
rect 2850 1415 2915 1465
rect 2965 1415 3000 1465
rect 2850 1285 3000 1415
rect 2850 1235 2915 1285
rect 2965 1235 3000 1285
rect 2850 1135 3000 1235
rect 2850 1085 2915 1135
rect 2965 1085 3000 1135
rect 2850 1050 3000 1085
<< psubstratepdiff >>
rect 180 205 300 240
rect 180 155 215 205
rect 265 155 300 205
rect 180 120 300 155
<< nsubstratendiff >>
rect 180 2125 300 2160
rect 180 2075 215 2125
rect 265 2075 300 2125
rect 180 1855 300 2075
rect 180 1805 215 1855
rect 265 1805 300 1855
rect 180 1770 300 1805
<< nsubstratencontact >>
rect 215 2075 265 2125
rect 215 1805 265 1855
<< psubstratepcontact >>
rect 215 155 265 205
<< ndcontact >>
rect 95 605 145 655
rect 95 455 145 505
rect 335 605 385 655
rect 335 455 385 505
rect 2675 605 2725 655
rect 2675 455 2725 505
rect 2675 305 2725 355
rect 2675 155 2725 205
rect 2915 605 2965 655
rect 2915 395 2965 445
rect 2915 215 2965 265
<< pdcontact >>
rect 95 1475 145 1525
rect 95 1265 145 1315
rect 95 1085 145 1135
rect 335 1475 385 1525
rect 2675 2165 2725 2215
rect 2675 1985 2725 2035
rect 2675 1835 2725 1885
rect 2675 1685 2725 1735
rect 2675 1535 2725 1585
rect 2675 1385 2725 1435
rect 335 1265 385 1315
rect 2675 1235 2725 1285
rect 335 1085 385 1135
rect 2915 2105 2965 2155
rect 2915 1955 2965 2005
rect 2915 1775 2965 1825
rect 2915 1595 2965 1645
rect 2915 1415 2965 1465
rect 2915 1235 2965 1285
rect 2915 1085 2965 1135
<< polysilicon >>
rect 720 2130 2460 2310
rect 2790 2250 2850 2315
rect 720 2125 900 2130
rect 720 2075 755 2125
rect 805 2075 900 2125
rect 720 1975 900 2075
rect 2280 2125 2460 2130
rect 2280 2075 2375 2125
rect 2425 2075 2460 2125
rect 720 1925 755 1975
rect 805 1925 900 1975
rect 720 1825 900 1925
rect 720 1775 755 1825
rect 805 1775 900 1825
rect 2280 1975 2460 2075
rect 2280 1925 2375 1975
rect 2425 1925 2460 1975
rect 2280 1825 2460 1925
rect 210 1620 270 1685
rect 720 1675 900 1775
rect 2280 1775 2375 1825
rect 2425 1775 2460 1825
rect 720 1625 755 1675
rect 805 1650 900 1675
rect 2280 1675 2460 1775
rect 2280 1650 2375 1675
rect 805 1625 2375 1650
rect 2425 1625 2460 1675
rect 720 1500 2460 1625
rect 210 960 270 1050
rect 60 895 270 960
rect 60 845 125 895
rect 175 845 270 895
rect 60 780 270 845
rect 210 690 270 780
rect 660 895 2460 990
rect 2790 960 2850 1050
rect 660 845 695 895
rect 745 860 2460 895
rect 745 845 840 860
rect 660 745 840 845
rect 660 695 695 745
rect 745 695 840 745
rect 2280 745 2460 860
rect 2640 895 2850 960
rect 2640 845 2705 895
rect 2755 845 2850 895
rect 2640 780 2850 845
rect 660 595 840 695
rect 2280 695 2375 745
rect 2425 695 2460 745
rect 2280 595 2460 695
rect 2790 690 2850 780
rect 660 545 695 595
rect 745 545 840 595
rect 2280 545 2375 595
rect 2425 545 2460 595
rect 660 445 840 545
rect 660 395 695 445
rect 745 395 840 445
rect 210 325 270 390
rect 660 295 840 395
rect 2280 445 2460 545
rect 2280 395 2375 445
rect 2425 395 2460 445
rect 660 245 695 295
rect 745 245 840 295
rect 660 160 840 245
rect 2280 295 2460 395
rect 2280 245 2375 295
rect 2425 245 2460 295
rect 2280 160 2460 245
rect 660 60 2460 160
rect 2790 55 2850 120
<< polycontact >>
rect 755 2075 805 2125
rect 2375 2075 2425 2125
rect 755 1925 805 1975
rect 755 1775 805 1825
rect 2375 1925 2425 1975
rect 2375 1775 2425 1825
rect 755 1625 805 1675
rect 2375 1625 2425 1675
rect 125 845 175 895
rect 695 845 745 895
rect 695 695 745 745
rect 2705 845 2755 895
rect 2375 695 2425 745
rect 695 545 745 595
rect 2375 545 2425 595
rect 695 395 745 445
rect 2375 395 2425 445
rect 695 245 745 295
rect 2375 245 2425 295
<< poly2 >>
rect 570 1330 720 1350
rect 570 1280 600 1330
rect 650 1280 720 1330
rect 570 1210 720 1280
rect 570 1160 600 1210
rect 650 1160 720 1210
rect 570 1140 720 1160
rect 2250 1330 2460 1350
rect 2250 1280 2360 1330
rect 2410 1280 2460 1330
rect 2250 1210 2460 1280
rect 2250 1160 2360 1210
rect 2410 1160 2460 1210
rect 2250 1140 2460 1160
<< poly2cap >>
rect 900 2035 2280 2130
rect 900 1985 1025 2035
rect 1075 1985 1175 2035
rect 1225 1985 1325 2035
rect 1375 1985 1475 2035
rect 1525 1985 1625 2035
rect 1675 1985 1775 2035
rect 1825 1985 1925 2035
rect 1975 1985 2075 2035
rect 2125 1985 2280 2035
rect 900 1795 2280 1985
rect 900 1745 1025 1795
rect 1075 1745 1175 1795
rect 1225 1745 1325 1795
rect 1375 1745 1475 1795
rect 1525 1745 1625 1795
rect 1675 1745 1775 1795
rect 1825 1745 1925 1795
rect 1975 1745 2075 1795
rect 2125 1745 2280 1795
rect 900 1650 2280 1745
rect 840 755 2280 860
rect 840 705 935 755
rect 985 705 1085 755
rect 1135 705 1235 755
rect 1285 705 1385 755
rect 1435 705 1535 755
rect 1585 705 1685 755
rect 1735 705 1835 755
rect 1885 705 1985 755
rect 2035 705 2135 755
rect 2185 705 2280 755
rect 840 595 2280 705
rect 840 545 935 595
rect 985 545 1085 595
rect 1135 545 1235 595
rect 1285 545 1385 595
rect 1435 545 1535 595
rect 1585 545 1685 595
rect 1735 545 1835 595
rect 1885 545 1985 595
rect 2035 545 2135 595
rect 2185 545 2280 595
rect 840 385 2280 545
rect 840 335 935 385
rect 985 335 1085 385
rect 1135 335 1235 385
rect 1285 335 1385 385
rect 1435 335 1535 385
rect 1585 335 1685 385
rect 1735 335 1835 385
rect 1885 335 1985 385
rect 2035 335 2135 385
rect 2185 335 2280 385
rect 840 160 2280 335
<< high_resist >>
rect 720 1350 2250 1450
rect 720 1040 2250 1140
<< poly2_high_resist >>
rect 720 1140 2250 1350
<< poly2contact >>
rect 600 1280 650 1330
rect 600 1160 650 1210
rect 2360 1280 2410 1330
rect 2360 1160 2410 1210
<< poly2capcontact >>
rect 1025 1985 1075 2035
rect 1175 1985 1225 2035
rect 1325 1985 1375 2035
rect 1475 1985 1525 2035
rect 1625 1985 1675 2035
rect 1775 1985 1825 2035
rect 1925 1985 1975 2035
rect 2075 1985 2125 2035
rect 1025 1745 1075 1795
rect 1175 1745 1225 1795
rect 1325 1745 1375 1795
rect 1475 1745 1525 1795
rect 1625 1745 1675 1795
rect 1775 1745 1825 1795
rect 1925 1745 1975 1795
rect 2075 1745 2125 1795
rect 935 705 985 755
rect 1085 705 1135 755
rect 1235 705 1285 755
rect 1385 705 1435 755
rect 1535 705 1585 755
rect 1685 705 1735 755
rect 1835 705 1885 755
rect 1985 705 2035 755
rect 2135 705 2185 755
rect 935 545 985 595
rect 1085 545 1135 595
rect 1235 545 1285 595
rect 1385 545 1435 595
rect 1535 545 1585 595
rect 1685 545 1735 595
rect 1835 545 1885 595
rect 1985 545 2035 595
rect 2135 545 2185 595
rect 935 335 985 385
rect 1085 335 1135 385
rect 1235 335 1285 385
rect 1385 335 1435 385
rect 1535 335 1585 385
rect 1685 335 1735 385
rect 1835 335 1885 385
rect 1985 335 2035 385
rect 2135 335 2185 385
<< metal1 >>
rect 0 2280 3060 2370
rect 60 2160 180 2280
rect 60 2125 300 2160
rect 60 2075 215 2125
rect 265 2075 300 2125
rect 60 1855 300 2075
rect 60 1805 215 1855
rect 265 1805 300 1855
rect 60 1770 300 1805
rect 720 2125 840 2190
rect 720 2075 755 2125
rect 805 2075 840 2125
rect 720 1975 840 2075
rect 720 1925 755 1975
rect 805 1925 840 1975
rect 720 1825 840 1925
rect 720 1775 755 1825
rect 805 1775 840 1825
rect 60 1525 180 1770
rect 720 1675 840 1775
rect 930 2035 2250 2280
rect 2640 2215 2760 2280
rect 930 1985 1025 2035
rect 1075 1985 1175 2035
rect 1225 1985 1325 2035
rect 1375 1985 1475 2035
rect 1525 1985 1625 2035
rect 1675 1985 1775 2035
rect 1825 1985 1925 2035
rect 1975 1985 2075 2035
rect 2125 1985 2250 2035
rect 930 1795 2250 1985
rect 930 1745 1025 1795
rect 1075 1745 1175 1795
rect 1225 1745 1325 1795
rect 1375 1745 1475 1795
rect 1525 1745 1625 1795
rect 1675 1745 1775 1795
rect 1825 1745 1925 1795
rect 1975 1745 2075 1795
rect 2125 1745 2250 1795
rect 930 1680 2250 1745
rect 2340 2125 2460 2190
rect 2340 2075 2375 2125
rect 2425 2075 2460 2125
rect 2340 1975 2460 2075
rect 2340 1925 2375 1975
rect 2425 1925 2460 1975
rect 2340 1825 2460 1925
rect 2340 1775 2375 1825
rect 2425 1775 2460 1825
rect 720 1625 755 1675
rect 805 1625 840 1675
rect 720 1620 840 1625
rect 2340 1675 2460 1775
rect 2340 1625 2375 1675
rect 2425 1625 2460 1675
rect 2340 1620 2460 1625
rect 60 1475 95 1525
rect 145 1475 180 1525
rect 60 1315 180 1475
rect 60 1265 95 1315
rect 145 1265 180 1315
rect 60 1135 180 1265
rect 60 1085 95 1135
rect 145 1085 180 1135
rect 60 1050 180 1085
rect 300 1525 420 1560
rect 300 1475 335 1525
rect 385 1475 420 1525
rect 720 1500 2460 1620
rect 300 1350 420 1475
rect 300 1330 690 1350
rect 300 1315 600 1330
rect 300 1265 335 1315
rect 385 1280 600 1315
rect 650 1280 690 1330
rect 385 1265 690 1280
rect 300 1210 690 1265
rect 300 1160 600 1210
rect 650 1160 690 1210
rect 300 1140 690 1160
rect 2310 1330 2460 1500
rect 2310 1280 2360 1330
rect 2410 1280 2460 1330
rect 2310 1210 2460 1280
rect 2310 1160 2360 1210
rect 2410 1160 2460 1210
rect 2640 2165 2675 2215
rect 2725 2165 2760 2215
rect 2640 2035 2760 2165
rect 2640 1985 2675 2035
rect 2725 1985 2760 2035
rect 2640 1885 2760 1985
rect 2640 1835 2675 1885
rect 2725 1835 2760 1885
rect 2640 1735 2760 1835
rect 2640 1685 2675 1735
rect 2725 1685 2760 1735
rect 2640 1585 2760 1685
rect 2640 1535 2675 1585
rect 2725 1535 2760 1585
rect 2640 1435 2760 1535
rect 2640 1385 2675 1435
rect 2725 1385 2760 1435
rect 2640 1285 2760 1385
rect 2640 1235 2675 1285
rect 2725 1235 2760 1285
rect 2640 1200 2760 1235
rect 2880 2155 3000 2190
rect 2880 2105 2915 2155
rect 2965 2105 3000 2155
rect 2880 2005 3000 2105
rect 2880 1955 2915 2005
rect 2965 1955 3000 2005
rect 2880 1825 3000 1955
rect 2880 1775 2915 1825
rect 2965 1775 3000 1825
rect 2880 1645 3000 1775
rect 2880 1595 2915 1645
rect 2965 1595 3000 1645
rect 2880 1465 3000 1595
rect 2880 1415 2915 1465
rect 2965 1415 3000 1465
rect 2880 1285 3000 1415
rect 2880 1235 2915 1285
rect 2965 1235 3000 1285
rect 300 1135 420 1140
rect 300 1085 335 1135
rect 385 1085 420 1135
rect 90 895 210 930
rect 90 845 125 895
rect 175 845 210 895
rect 90 810 210 845
rect 60 655 180 690
rect 60 605 95 655
rect 145 605 180 655
rect 60 505 180 605
rect 60 455 95 505
rect 145 455 180 505
rect 60 270 180 455
rect 300 655 420 1085
rect 2310 1110 2460 1160
rect 2880 1135 3000 1235
rect 2310 990 2790 1110
rect 300 605 335 655
rect 385 605 420 655
rect 300 505 420 605
rect 300 455 335 505
rect 385 455 420 505
rect 300 420 420 455
rect 660 895 2460 990
rect 660 845 695 895
rect 745 870 2460 895
rect 745 845 780 870
rect 660 745 780 845
rect 660 695 695 745
rect 745 695 780 745
rect 660 595 780 695
rect 660 545 695 595
rect 745 545 780 595
rect 660 445 780 545
rect 660 395 695 445
rect 745 395 780 445
rect 660 295 780 395
rect 60 205 300 270
rect 60 155 215 205
rect 265 155 300 205
rect 660 245 695 295
rect 745 245 780 295
rect 660 180 780 245
rect 870 755 2250 780
rect 870 705 935 755
rect 985 705 1085 755
rect 1135 705 1235 755
rect 1285 705 1385 755
rect 1435 705 1535 755
rect 1585 705 1685 755
rect 1735 705 1835 755
rect 1885 705 1985 755
rect 2035 705 2135 755
rect 2185 705 2250 755
rect 870 595 2250 705
rect 870 545 935 595
rect 985 545 1085 595
rect 1135 545 1235 595
rect 1285 545 1385 595
rect 1435 545 1535 595
rect 1585 545 1685 595
rect 1735 545 1835 595
rect 1885 545 1985 595
rect 2035 545 2135 595
rect 2185 545 2250 595
rect 870 385 2250 545
rect 870 335 935 385
rect 985 335 1085 385
rect 1135 335 1235 385
rect 1285 335 1385 385
rect 1435 335 1535 385
rect 1585 335 1685 385
rect 1735 335 1835 385
rect 1885 335 1985 385
rect 2035 335 2135 385
rect 2185 335 2250 385
rect 60 90 300 155
rect 870 90 2250 335
rect 2340 745 2460 870
rect 2670 895 2790 990
rect 2670 845 2705 895
rect 2755 845 2790 895
rect 2670 810 2790 845
rect 2880 1085 2915 1135
rect 2965 1085 3000 1135
rect 2340 695 2375 745
rect 2425 695 2460 745
rect 2340 595 2460 695
rect 2340 545 2375 595
rect 2425 545 2460 595
rect 2340 445 2460 545
rect 2340 395 2375 445
rect 2425 395 2460 445
rect 2340 295 2460 395
rect 2340 245 2375 295
rect 2425 245 2460 295
rect 2340 180 2460 245
rect 2640 655 2760 690
rect 2640 605 2675 655
rect 2725 605 2760 655
rect 2640 505 2760 605
rect 2640 455 2675 505
rect 2725 455 2760 505
rect 2640 355 2760 455
rect 2640 305 2675 355
rect 2725 305 2760 355
rect 2640 205 2760 305
rect 2640 155 2675 205
rect 2725 155 2760 205
rect 2880 655 3000 1085
rect 2880 605 2915 655
rect 2965 605 3000 655
rect 2880 445 3000 605
rect 2880 395 2915 445
rect 2965 395 3000 445
rect 2880 265 3000 395
rect 2880 215 2915 265
rect 2965 215 3000 265
rect 2880 180 3000 215
rect 2640 90 2760 155
rect 0 0 3060 90
<< labels >>
flabel metal1 s 330 780 330 780 2 FreeSans 400 0 0 0 n1
flabel metal1 s 150 870 150 870 2 FreeSans 400 0 0 0 a
port 2 ne
flabel metal1 s 30 2340 30 2340 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 30 30 30 30 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 2940 810 2940 810 2 FreeSans 400 0 0 0 z
port 1 ne
flabel poly2_high_resist s 1320 1260 1320 1260 2 FreeSans 400 0 0 0 r0
flabel metal1 s 2370 1380 2370 1380 2 FreeSans 400 0 0 0 n2
<< end >>
