`celldefine
module fill2 ();
endmodule
`endcelldefine
