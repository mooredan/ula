magic
tech scmos
magscale 1 2
timestamp 1572801172
<< error_p >>
rect 2 1332 10 1334
rect 2 1328 4 1332
rect 8 1328 10 1332
rect 2 1326 10 1328
rect 14 1332 22 1334
rect 14 1328 16 1332
rect 20 1328 22 1332
rect 14 1326 22 1328
rect 24 1332 32 1334
rect 24 1328 26 1332
rect 30 1328 32 1332
rect 24 1326 32 1328
rect 34 1332 42 1334
rect 34 1328 36 1332
rect 40 1328 42 1332
rect 34 1326 42 1328
rect 44 1332 52 1334
rect 44 1328 46 1332
rect 50 1328 52 1332
rect 44 1326 52 1328
rect 54 1332 62 1334
rect 54 1328 56 1332
rect 60 1328 62 1332
rect 54 1326 62 1328
rect 64 1332 72 1334
rect 64 1328 66 1332
rect 70 1328 72 1332
rect 64 1326 72 1328
rect 74 1332 82 1334
rect 74 1328 76 1332
rect 80 1328 82 1332
rect 74 1326 82 1328
rect 84 1332 92 1334
rect 84 1328 86 1332
rect 90 1328 92 1332
rect 84 1326 92 1328
rect 94 1332 102 1334
rect 94 1328 96 1332
rect 100 1328 102 1332
rect 94 1326 102 1328
rect 104 1332 112 1334
rect 104 1328 106 1332
rect 110 1328 112 1332
rect 104 1326 112 1328
rect 114 1332 122 1334
rect 114 1328 116 1332
rect 120 1328 122 1332
rect 114 1326 122 1328
rect 124 1332 132 1334
rect 124 1328 126 1332
rect 130 1328 132 1332
rect 124 1326 132 1328
rect 134 1332 142 1334
rect 134 1328 136 1332
rect 140 1328 142 1332
rect 134 1326 142 1328
rect 144 1332 152 1334
rect 144 1328 146 1332
rect 150 1328 152 1332
rect 144 1326 152 1328
rect 154 1332 162 1334
rect 154 1328 156 1332
rect 160 1328 162 1332
rect 154 1326 162 1328
rect 164 1332 172 1334
rect 164 1328 166 1332
rect 170 1328 172 1332
rect 164 1326 172 1328
rect 174 1332 182 1334
rect 174 1328 176 1332
rect 180 1328 182 1332
rect 174 1326 182 1328
rect 184 1332 192 1334
rect 184 1328 186 1332
rect 190 1328 192 1332
rect 184 1326 192 1328
rect 194 1332 202 1334
rect 194 1328 196 1332
rect 200 1328 202 1332
rect 194 1326 202 1328
rect 204 1332 212 1334
rect 204 1328 206 1332
rect 210 1328 212 1332
rect 204 1326 212 1328
rect 214 1332 222 1334
rect 214 1328 216 1332
rect 220 1328 222 1332
rect 214 1326 222 1328
rect 224 1332 232 1334
rect 224 1328 226 1332
rect 230 1328 232 1332
rect 224 1326 232 1328
rect 368 1332 376 1334
rect 368 1328 370 1332
rect 374 1328 376 1332
rect 368 1326 376 1328
rect 378 1332 386 1334
rect 378 1328 380 1332
rect 384 1328 386 1332
rect 378 1326 386 1328
rect 388 1332 396 1334
rect 388 1328 390 1332
rect 394 1328 396 1332
rect 388 1326 396 1328
rect 398 1332 406 1334
rect 398 1328 400 1332
rect 404 1328 406 1332
rect 398 1326 406 1328
rect 408 1332 416 1334
rect 408 1328 410 1332
rect 414 1328 416 1332
rect 408 1326 416 1328
rect 418 1332 426 1334
rect 418 1328 420 1332
rect 424 1328 426 1332
rect 418 1326 426 1328
rect 428 1332 436 1334
rect 428 1328 430 1332
rect 434 1328 436 1332
rect 428 1326 436 1328
rect 438 1332 446 1334
rect 438 1328 440 1332
rect 444 1328 446 1332
rect 438 1326 446 1328
rect 448 1332 456 1334
rect 448 1328 450 1332
rect 454 1328 456 1332
rect 448 1326 456 1328
rect 458 1332 466 1334
rect 458 1328 460 1332
rect 464 1328 466 1332
rect 458 1326 466 1328
rect 468 1332 476 1334
rect 468 1328 470 1332
rect 474 1328 476 1332
rect 468 1326 476 1328
rect 478 1332 486 1334
rect 478 1328 480 1332
rect 484 1328 486 1332
rect 478 1326 486 1328
rect 488 1332 496 1334
rect 488 1328 490 1332
rect 494 1328 496 1332
rect 488 1326 496 1328
rect 498 1332 506 1334
rect 498 1328 500 1332
rect 504 1328 506 1332
rect 498 1326 506 1328
rect 508 1332 516 1334
rect 508 1328 510 1332
rect 514 1328 516 1332
rect 508 1326 516 1328
rect 518 1332 526 1334
rect 518 1328 520 1332
rect 524 1328 526 1332
rect 518 1326 526 1328
rect 528 1332 536 1334
rect 528 1328 530 1332
rect 534 1328 536 1332
rect 528 1326 536 1328
rect 538 1332 546 1334
rect 538 1328 540 1332
rect 544 1328 546 1332
rect 538 1326 546 1328
rect 548 1332 556 1334
rect 548 1328 550 1332
rect 554 1328 556 1332
rect 548 1326 556 1328
rect 558 1332 566 1334
rect 558 1328 560 1332
rect 564 1328 566 1332
rect 558 1326 566 1328
rect 568 1332 576 1334
rect 568 1328 570 1332
rect 574 1328 576 1332
rect 568 1326 576 1328
rect 580 1330 588 1332
rect 580 1326 582 1330
rect 586 1326 588 1330
rect 580 1324 588 1326
rect 590 1330 598 1332
rect 590 1326 592 1330
rect 596 1326 598 1330
rect 590 1324 598 1326
rect 2 1322 10 1324
rect 2 1318 4 1322
rect 8 1318 10 1322
rect 2 1316 10 1318
rect 14 1322 22 1324
rect 14 1318 16 1322
rect 20 1318 22 1322
rect 14 1316 22 1318
rect 24 1322 32 1324
rect 24 1318 26 1322
rect 30 1318 32 1322
rect 24 1316 32 1318
rect 34 1322 42 1324
rect 34 1318 36 1322
rect 40 1318 42 1322
rect 34 1316 42 1318
rect 44 1322 52 1324
rect 44 1318 46 1322
rect 50 1318 52 1322
rect 44 1316 52 1318
rect 54 1322 62 1324
rect 54 1318 56 1322
rect 60 1318 62 1322
rect 54 1316 62 1318
rect 64 1322 72 1324
rect 64 1318 66 1322
rect 70 1318 72 1322
rect 64 1316 72 1318
rect 74 1322 82 1324
rect 74 1318 76 1322
rect 80 1318 82 1322
rect 74 1316 82 1318
rect 84 1322 92 1324
rect 84 1318 86 1322
rect 90 1318 92 1322
rect 84 1316 92 1318
rect 94 1322 102 1324
rect 94 1318 96 1322
rect 100 1318 102 1322
rect 94 1316 102 1318
rect 104 1322 112 1324
rect 104 1318 106 1322
rect 110 1318 112 1322
rect 104 1316 112 1318
rect 114 1322 122 1324
rect 114 1318 116 1322
rect 120 1318 122 1322
rect 114 1316 122 1318
rect 124 1322 132 1324
rect 124 1318 126 1322
rect 130 1318 132 1322
rect 124 1316 132 1318
rect 134 1322 142 1324
rect 134 1318 136 1322
rect 140 1318 142 1322
rect 134 1316 142 1318
rect 144 1322 152 1324
rect 144 1318 146 1322
rect 150 1318 152 1322
rect 144 1316 152 1318
rect 154 1322 162 1324
rect 154 1318 156 1322
rect 160 1318 162 1322
rect 154 1316 162 1318
rect 164 1322 172 1324
rect 164 1318 166 1322
rect 170 1318 172 1322
rect 164 1316 172 1318
rect 174 1322 182 1324
rect 174 1318 176 1322
rect 180 1318 182 1322
rect 174 1316 182 1318
rect 184 1322 192 1324
rect 184 1318 186 1322
rect 190 1318 192 1322
rect 184 1316 192 1318
rect 194 1322 202 1324
rect 194 1318 196 1322
rect 200 1318 202 1322
rect 194 1316 202 1318
rect 204 1322 212 1324
rect 204 1318 206 1322
rect 210 1318 212 1322
rect 204 1316 212 1318
rect 214 1322 222 1324
rect 214 1318 216 1322
rect 220 1318 222 1322
rect 214 1316 222 1318
rect 224 1322 232 1324
rect 224 1318 226 1322
rect 230 1318 232 1322
rect 224 1316 232 1318
rect 368 1322 376 1324
rect 368 1318 370 1322
rect 374 1318 376 1322
rect 368 1316 376 1318
rect 378 1322 386 1324
rect 378 1318 380 1322
rect 384 1318 386 1322
rect 378 1316 386 1318
rect 388 1322 396 1324
rect 388 1318 390 1322
rect 394 1318 396 1322
rect 388 1316 396 1318
rect 398 1322 406 1324
rect 398 1318 400 1322
rect 404 1318 406 1322
rect 398 1316 406 1318
rect 408 1322 416 1324
rect 408 1318 410 1322
rect 414 1318 416 1322
rect 408 1316 416 1318
rect 418 1322 426 1324
rect 418 1318 420 1322
rect 424 1318 426 1322
rect 418 1316 426 1318
rect 428 1322 436 1324
rect 428 1318 430 1322
rect 434 1318 436 1322
rect 428 1316 436 1318
rect 438 1322 446 1324
rect 438 1318 440 1322
rect 444 1318 446 1322
rect 438 1316 446 1318
rect 448 1322 456 1324
rect 448 1318 450 1322
rect 454 1318 456 1322
rect 448 1316 456 1318
rect 458 1322 466 1324
rect 458 1318 460 1322
rect 464 1318 466 1322
rect 458 1316 466 1318
rect 468 1322 476 1324
rect 468 1318 470 1322
rect 474 1318 476 1322
rect 468 1316 476 1318
rect 478 1322 486 1324
rect 478 1318 480 1322
rect 484 1318 486 1322
rect 478 1316 486 1318
rect 488 1322 496 1324
rect 488 1318 490 1322
rect 494 1318 496 1322
rect 488 1316 496 1318
rect 498 1322 506 1324
rect 498 1318 500 1322
rect 504 1318 506 1322
rect 498 1316 506 1318
rect 508 1322 516 1324
rect 508 1318 510 1322
rect 514 1318 516 1322
rect 508 1316 516 1318
rect 518 1322 526 1324
rect 518 1318 520 1322
rect 524 1318 526 1322
rect 518 1316 526 1318
rect 528 1322 536 1324
rect 528 1318 530 1322
rect 534 1318 536 1322
rect 528 1316 536 1318
rect 538 1322 546 1324
rect 538 1318 540 1322
rect 544 1318 546 1322
rect 538 1316 546 1318
rect 548 1322 556 1324
rect 548 1318 550 1322
rect 554 1318 556 1322
rect 548 1316 556 1318
rect 558 1322 566 1324
rect 558 1318 560 1322
rect 564 1318 566 1322
rect 558 1316 566 1318
rect 568 1322 576 1324
rect 568 1318 570 1322
rect 574 1318 576 1322
rect 568 1316 576 1318
rect 580 1320 588 1322
rect 580 1316 582 1320
rect 586 1316 588 1320
rect 580 1314 588 1316
rect 590 1320 598 1322
rect 590 1316 592 1320
rect 596 1316 598 1320
rect 590 1314 598 1316
rect 2 1312 10 1314
rect 2 1308 4 1312
rect 8 1308 10 1312
rect 2 1306 10 1308
rect 12 1312 20 1314
rect 12 1308 14 1312
rect 18 1308 20 1312
rect 580 1310 588 1312
rect 374 1308 382 1310
rect 12 1306 20 1308
rect 28 1306 36 1308
rect 2 1302 10 1304
rect 2 1298 4 1302
rect 8 1298 10 1302
rect 2 1296 10 1298
rect 12 1302 20 1304
rect 12 1298 14 1302
rect 18 1298 20 1302
rect 28 1302 30 1306
rect 34 1302 36 1306
rect 28 1300 36 1302
rect 38 1306 46 1308
rect 38 1302 40 1306
rect 44 1302 46 1306
rect 38 1300 46 1302
rect 48 1306 56 1308
rect 48 1302 50 1306
rect 54 1302 56 1306
rect 48 1300 56 1302
rect 58 1306 66 1308
rect 58 1302 60 1306
rect 64 1302 66 1306
rect 58 1300 66 1302
rect 68 1306 76 1308
rect 68 1302 70 1306
rect 74 1302 76 1306
rect 68 1300 76 1302
rect 78 1306 86 1308
rect 78 1302 80 1306
rect 84 1302 86 1306
rect 78 1300 86 1302
rect 88 1306 96 1308
rect 88 1302 90 1306
rect 94 1302 96 1306
rect 88 1300 96 1302
rect 98 1306 106 1308
rect 98 1302 100 1306
rect 104 1302 106 1306
rect 98 1300 106 1302
rect 108 1306 116 1308
rect 108 1302 110 1306
rect 114 1302 116 1306
rect 108 1300 116 1302
rect 118 1306 126 1308
rect 118 1302 120 1306
rect 124 1302 126 1306
rect 118 1300 126 1302
rect 128 1306 136 1308
rect 128 1302 130 1306
rect 134 1302 136 1306
rect 128 1300 136 1302
rect 138 1306 146 1308
rect 138 1302 140 1306
rect 144 1302 146 1306
rect 138 1300 146 1302
rect 148 1306 156 1308
rect 148 1302 150 1306
rect 154 1302 156 1306
rect 148 1300 156 1302
rect 158 1306 166 1308
rect 158 1302 160 1306
rect 164 1302 166 1306
rect 158 1300 166 1302
rect 168 1306 176 1308
rect 168 1302 170 1306
rect 174 1302 176 1306
rect 168 1300 176 1302
rect 178 1306 186 1308
rect 178 1302 180 1306
rect 184 1302 186 1306
rect 178 1300 186 1302
rect 188 1306 196 1308
rect 188 1302 190 1306
rect 194 1302 196 1306
rect 188 1300 196 1302
rect 198 1306 206 1308
rect 198 1302 200 1306
rect 204 1302 206 1306
rect 198 1300 206 1302
rect 208 1306 216 1308
rect 208 1302 210 1306
rect 214 1302 216 1306
rect 208 1300 216 1302
rect 218 1306 226 1308
rect 218 1302 220 1306
rect 224 1302 226 1306
rect 374 1304 376 1308
rect 380 1304 382 1308
rect 374 1302 382 1304
rect 384 1308 392 1310
rect 384 1304 386 1308
rect 390 1304 392 1308
rect 384 1302 392 1304
rect 394 1308 402 1310
rect 394 1304 396 1308
rect 400 1304 402 1308
rect 394 1302 402 1304
rect 404 1308 412 1310
rect 404 1304 406 1308
rect 410 1304 412 1308
rect 404 1302 412 1304
rect 414 1308 422 1310
rect 414 1304 416 1308
rect 420 1304 422 1308
rect 414 1302 422 1304
rect 424 1308 432 1310
rect 424 1304 426 1308
rect 430 1304 432 1308
rect 424 1302 432 1304
rect 434 1308 442 1310
rect 434 1304 436 1308
rect 440 1304 442 1308
rect 434 1302 442 1304
rect 444 1308 452 1310
rect 444 1304 446 1308
rect 450 1304 452 1308
rect 444 1302 452 1304
rect 454 1308 462 1310
rect 454 1304 456 1308
rect 460 1304 462 1308
rect 454 1302 462 1304
rect 464 1308 472 1310
rect 464 1304 466 1308
rect 470 1304 472 1308
rect 464 1302 472 1304
rect 474 1308 482 1310
rect 474 1304 476 1308
rect 480 1304 482 1308
rect 474 1302 482 1304
rect 484 1308 492 1310
rect 484 1304 486 1308
rect 490 1304 492 1308
rect 484 1302 492 1304
rect 494 1308 502 1310
rect 494 1304 496 1308
rect 500 1304 502 1308
rect 494 1302 502 1304
rect 504 1308 512 1310
rect 504 1304 506 1308
rect 510 1304 512 1308
rect 504 1302 512 1304
rect 514 1308 522 1310
rect 514 1304 516 1308
rect 520 1304 522 1308
rect 514 1302 522 1304
rect 524 1308 532 1310
rect 524 1304 526 1308
rect 530 1304 532 1308
rect 524 1302 532 1304
rect 534 1308 542 1310
rect 534 1304 536 1308
rect 540 1304 542 1308
rect 534 1302 542 1304
rect 544 1308 552 1310
rect 544 1304 546 1308
rect 550 1304 552 1308
rect 544 1302 552 1304
rect 554 1308 562 1310
rect 554 1304 556 1308
rect 560 1304 562 1308
rect 554 1302 562 1304
rect 564 1308 572 1310
rect 564 1304 566 1308
rect 570 1304 572 1308
rect 580 1306 582 1310
rect 586 1306 588 1310
rect 580 1304 588 1306
rect 590 1310 598 1312
rect 590 1306 592 1310
rect 596 1306 598 1310
rect 590 1304 598 1306
rect 564 1302 572 1304
rect 218 1300 226 1302
rect 580 1300 588 1302
rect 564 1298 572 1300
rect 12 1296 20 1298
rect 28 1296 36 1298
rect 2 1292 10 1294
rect 2 1288 4 1292
rect 8 1288 10 1292
rect 2 1286 10 1288
rect 12 1292 20 1294
rect 12 1288 14 1292
rect 18 1288 20 1292
rect 28 1292 30 1296
rect 34 1292 36 1296
rect 564 1294 566 1298
rect 570 1294 572 1298
rect 580 1296 582 1300
rect 586 1296 588 1300
rect 580 1294 588 1296
rect 590 1300 598 1302
rect 590 1296 592 1300
rect 596 1296 598 1300
rect 590 1294 598 1296
rect 28 1290 36 1292
rect 296 1292 304 1294
rect 564 1292 572 1294
rect 40 1288 48 1290
rect 12 1286 20 1288
rect 28 1286 36 1288
rect 2 1282 10 1284
rect 2 1278 4 1282
rect 8 1278 10 1282
rect 2 1276 10 1278
rect 12 1282 20 1284
rect 12 1278 14 1282
rect 18 1278 20 1282
rect 28 1282 30 1286
rect 34 1282 36 1286
rect 40 1284 42 1288
rect 46 1284 48 1288
rect 40 1282 48 1284
rect 50 1288 58 1290
rect 50 1284 52 1288
rect 56 1284 58 1288
rect 50 1282 58 1284
rect 60 1288 68 1290
rect 60 1284 62 1288
rect 66 1284 68 1288
rect 60 1282 68 1284
rect 70 1288 78 1290
rect 70 1284 72 1288
rect 76 1284 78 1288
rect 70 1282 78 1284
rect 80 1288 88 1290
rect 80 1284 82 1288
rect 86 1284 88 1288
rect 80 1282 88 1284
rect 90 1288 98 1290
rect 90 1284 92 1288
rect 96 1284 98 1288
rect 90 1282 98 1284
rect 100 1288 108 1290
rect 100 1284 102 1288
rect 106 1284 108 1288
rect 100 1282 108 1284
rect 112 1288 120 1290
rect 112 1284 114 1288
rect 118 1284 120 1288
rect 112 1282 120 1284
rect 122 1288 130 1290
rect 122 1284 124 1288
rect 128 1284 130 1288
rect 122 1282 130 1284
rect 132 1288 140 1290
rect 132 1284 134 1288
rect 138 1284 140 1288
rect 132 1282 140 1284
rect 142 1288 150 1290
rect 142 1284 144 1288
rect 148 1284 150 1288
rect 142 1282 150 1284
rect 152 1288 160 1290
rect 152 1284 154 1288
rect 158 1284 160 1288
rect 152 1282 160 1284
rect 162 1288 170 1290
rect 162 1284 164 1288
rect 168 1284 170 1288
rect 162 1282 170 1284
rect 172 1288 180 1290
rect 172 1284 174 1288
rect 178 1284 180 1288
rect 172 1282 180 1284
rect 182 1288 190 1290
rect 182 1284 184 1288
rect 188 1284 190 1288
rect 182 1282 190 1284
rect 192 1288 200 1290
rect 192 1284 194 1288
rect 198 1284 200 1288
rect 192 1282 200 1284
rect 202 1288 210 1290
rect 202 1284 204 1288
rect 208 1284 210 1288
rect 202 1282 210 1284
rect 212 1288 220 1290
rect 212 1284 214 1288
rect 218 1284 220 1288
rect 212 1282 220 1284
rect 222 1288 230 1290
rect 222 1284 224 1288
rect 228 1284 230 1288
rect 296 1288 298 1292
rect 302 1288 304 1292
rect 580 1290 588 1292
rect 296 1286 304 1288
rect 366 1288 374 1290
rect 366 1284 368 1288
rect 372 1284 374 1288
rect 222 1282 230 1284
rect 296 1282 304 1284
rect 366 1282 374 1284
rect 376 1288 384 1290
rect 376 1284 378 1288
rect 382 1284 384 1288
rect 376 1282 384 1284
rect 386 1288 394 1290
rect 386 1284 388 1288
rect 392 1284 394 1288
rect 386 1282 394 1284
rect 396 1288 404 1290
rect 396 1284 398 1288
rect 402 1284 404 1288
rect 396 1282 404 1284
rect 406 1288 414 1290
rect 406 1284 408 1288
rect 412 1284 414 1288
rect 406 1282 414 1284
rect 416 1288 424 1290
rect 416 1284 418 1288
rect 422 1284 424 1288
rect 416 1282 424 1284
rect 426 1288 434 1290
rect 426 1284 428 1288
rect 432 1284 434 1288
rect 426 1282 434 1284
rect 436 1288 444 1290
rect 436 1284 438 1288
rect 442 1284 444 1288
rect 436 1282 444 1284
rect 446 1288 454 1290
rect 446 1284 448 1288
rect 452 1284 454 1288
rect 446 1282 454 1284
rect 456 1288 464 1290
rect 456 1284 458 1288
rect 462 1284 464 1288
rect 456 1282 464 1284
rect 466 1288 474 1290
rect 466 1284 468 1288
rect 472 1284 474 1288
rect 466 1282 474 1284
rect 476 1288 484 1290
rect 476 1284 478 1288
rect 482 1284 484 1288
rect 476 1282 484 1284
rect 488 1288 496 1290
rect 488 1284 490 1288
rect 494 1284 496 1288
rect 488 1282 496 1284
rect 498 1288 506 1290
rect 498 1284 500 1288
rect 504 1284 506 1288
rect 498 1282 506 1284
rect 508 1288 516 1290
rect 508 1284 510 1288
rect 514 1284 516 1288
rect 508 1282 516 1284
rect 518 1288 526 1290
rect 518 1284 520 1288
rect 524 1284 526 1288
rect 518 1282 526 1284
rect 528 1288 536 1290
rect 528 1284 530 1288
rect 534 1284 536 1288
rect 528 1282 536 1284
rect 542 1288 550 1290
rect 542 1284 544 1288
rect 548 1284 550 1288
rect 542 1282 550 1284
rect 552 1288 560 1290
rect 552 1284 554 1288
rect 558 1284 560 1288
rect 552 1282 560 1284
rect 564 1288 572 1290
rect 564 1284 566 1288
rect 570 1284 572 1288
rect 580 1286 582 1290
rect 586 1286 588 1290
rect 580 1284 588 1286
rect 590 1290 598 1292
rect 590 1286 592 1290
rect 596 1286 598 1290
rect 590 1284 598 1286
rect 564 1282 572 1284
rect 28 1280 36 1282
rect 40 1278 48 1280
rect 12 1276 20 1278
rect 28 1276 36 1278
rect 2 1272 10 1274
rect 2 1268 4 1272
rect 8 1268 10 1272
rect 2 1266 10 1268
rect 12 1272 20 1274
rect 12 1268 14 1272
rect 18 1268 20 1272
rect 28 1272 30 1276
rect 34 1272 36 1276
rect 40 1274 42 1278
rect 46 1274 48 1278
rect 40 1272 48 1274
rect 50 1278 58 1280
rect 50 1274 52 1278
rect 56 1274 58 1278
rect 50 1272 58 1274
rect 60 1278 68 1280
rect 60 1274 62 1278
rect 66 1274 68 1278
rect 60 1272 68 1274
rect 70 1278 78 1280
rect 70 1274 72 1278
rect 76 1274 78 1278
rect 70 1272 78 1274
rect 80 1278 88 1280
rect 80 1274 82 1278
rect 86 1274 88 1278
rect 80 1272 88 1274
rect 90 1278 98 1280
rect 90 1274 92 1278
rect 96 1274 98 1278
rect 90 1272 98 1274
rect 100 1278 108 1280
rect 100 1274 102 1278
rect 106 1274 108 1278
rect 100 1272 108 1274
rect 112 1278 120 1280
rect 112 1274 114 1278
rect 118 1274 120 1278
rect 112 1272 120 1274
rect 122 1278 130 1280
rect 122 1274 124 1278
rect 128 1274 130 1278
rect 122 1272 130 1274
rect 132 1278 140 1280
rect 132 1274 134 1278
rect 138 1274 140 1278
rect 132 1272 140 1274
rect 142 1278 150 1280
rect 142 1274 144 1278
rect 148 1274 150 1278
rect 142 1272 150 1274
rect 152 1278 160 1280
rect 152 1274 154 1278
rect 158 1274 160 1278
rect 152 1272 160 1274
rect 162 1278 170 1280
rect 162 1274 164 1278
rect 168 1274 170 1278
rect 162 1272 170 1274
rect 172 1278 180 1280
rect 172 1274 174 1278
rect 178 1274 180 1278
rect 172 1272 180 1274
rect 182 1278 190 1280
rect 182 1274 184 1278
rect 188 1274 190 1278
rect 182 1272 190 1274
rect 192 1278 200 1280
rect 192 1274 194 1278
rect 198 1274 200 1278
rect 192 1272 200 1274
rect 202 1278 210 1280
rect 202 1274 204 1278
rect 208 1274 210 1278
rect 202 1272 210 1274
rect 212 1278 220 1280
rect 212 1274 214 1278
rect 218 1274 220 1278
rect 212 1272 220 1274
rect 222 1278 230 1280
rect 222 1274 224 1278
rect 228 1274 230 1278
rect 296 1278 298 1282
rect 302 1278 304 1282
rect 580 1280 588 1282
rect 296 1276 304 1278
rect 366 1278 374 1280
rect 366 1274 368 1278
rect 372 1274 374 1278
rect 222 1272 230 1274
rect 296 1272 304 1274
rect 366 1272 374 1274
rect 376 1278 384 1280
rect 376 1274 378 1278
rect 382 1274 384 1278
rect 376 1272 384 1274
rect 386 1278 394 1280
rect 386 1274 388 1278
rect 392 1274 394 1278
rect 386 1272 394 1274
rect 396 1278 404 1280
rect 396 1274 398 1278
rect 402 1274 404 1278
rect 396 1272 404 1274
rect 406 1278 414 1280
rect 406 1274 408 1278
rect 412 1274 414 1278
rect 406 1272 414 1274
rect 416 1278 424 1280
rect 416 1274 418 1278
rect 422 1274 424 1278
rect 416 1272 424 1274
rect 426 1278 434 1280
rect 426 1274 428 1278
rect 432 1274 434 1278
rect 426 1272 434 1274
rect 436 1278 444 1280
rect 436 1274 438 1278
rect 442 1274 444 1278
rect 436 1272 444 1274
rect 446 1278 454 1280
rect 446 1274 448 1278
rect 452 1274 454 1278
rect 446 1272 454 1274
rect 456 1278 464 1280
rect 456 1274 458 1278
rect 462 1274 464 1278
rect 456 1272 464 1274
rect 466 1278 474 1280
rect 466 1274 468 1278
rect 472 1274 474 1278
rect 466 1272 474 1274
rect 476 1278 484 1280
rect 476 1274 478 1278
rect 482 1274 484 1278
rect 476 1272 484 1274
rect 488 1278 496 1280
rect 488 1274 490 1278
rect 494 1274 496 1278
rect 488 1272 496 1274
rect 498 1278 506 1280
rect 498 1274 500 1278
rect 504 1274 506 1278
rect 498 1272 506 1274
rect 508 1278 516 1280
rect 508 1274 510 1278
rect 514 1274 516 1278
rect 508 1272 516 1274
rect 518 1278 526 1280
rect 518 1274 520 1278
rect 524 1274 526 1278
rect 518 1272 526 1274
rect 528 1278 536 1280
rect 528 1274 530 1278
rect 534 1274 536 1278
rect 528 1272 536 1274
rect 542 1278 550 1280
rect 542 1274 544 1278
rect 548 1274 550 1278
rect 542 1272 550 1274
rect 552 1278 560 1280
rect 552 1274 554 1278
rect 558 1274 560 1278
rect 552 1272 560 1274
rect 564 1278 572 1280
rect 564 1274 566 1278
rect 570 1274 572 1278
rect 580 1276 582 1280
rect 586 1276 588 1280
rect 580 1274 588 1276
rect 590 1280 598 1282
rect 590 1276 592 1280
rect 596 1276 598 1280
rect 590 1274 598 1276
rect 564 1272 572 1274
rect 28 1270 36 1272
rect 40 1268 48 1270
rect 12 1266 20 1268
rect 28 1266 36 1268
rect 2 1262 10 1264
rect 2 1258 4 1262
rect 8 1258 10 1262
rect 2 1256 10 1258
rect 12 1262 20 1264
rect 12 1258 14 1262
rect 18 1258 20 1262
rect 28 1262 30 1266
rect 34 1262 36 1266
rect 40 1264 42 1268
rect 46 1264 48 1268
rect 40 1262 48 1264
rect 50 1268 58 1270
rect 50 1264 52 1268
rect 56 1264 58 1268
rect 50 1262 58 1264
rect 60 1268 68 1270
rect 60 1264 62 1268
rect 66 1264 68 1268
rect 60 1262 68 1264
rect 70 1268 78 1270
rect 70 1264 72 1268
rect 76 1264 78 1268
rect 70 1262 78 1264
rect 80 1268 88 1270
rect 80 1264 82 1268
rect 86 1264 88 1268
rect 80 1262 88 1264
rect 90 1268 98 1270
rect 90 1264 92 1268
rect 96 1264 98 1268
rect 90 1262 98 1264
rect 100 1268 108 1270
rect 100 1264 102 1268
rect 106 1264 108 1268
rect 100 1262 108 1264
rect 112 1268 120 1270
rect 112 1264 114 1268
rect 118 1264 120 1268
rect 112 1262 120 1264
rect 122 1268 130 1270
rect 122 1264 124 1268
rect 128 1264 130 1268
rect 122 1262 130 1264
rect 132 1268 140 1270
rect 132 1264 134 1268
rect 138 1264 140 1268
rect 132 1262 140 1264
rect 142 1268 150 1270
rect 142 1264 144 1268
rect 148 1264 150 1268
rect 142 1262 150 1264
rect 152 1268 160 1270
rect 152 1264 154 1268
rect 158 1264 160 1268
rect 152 1262 160 1264
rect 162 1268 170 1270
rect 162 1264 164 1268
rect 168 1264 170 1268
rect 162 1262 170 1264
rect 172 1268 180 1270
rect 172 1264 174 1268
rect 178 1264 180 1268
rect 172 1262 180 1264
rect 182 1268 190 1270
rect 182 1264 184 1268
rect 188 1264 190 1268
rect 182 1262 190 1264
rect 192 1268 200 1270
rect 192 1264 194 1268
rect 198 1264 200 1268
rect 192 1262 200 1264
rect 202 1268 210 1270
rect 202 1264 204 1268
rect 208 1264 210 1268
rect 202 1262 210 1264
rect 212 1268 220 1270
rect 212 1264 214 1268
rect 218 1264 220 1268
rect 212 1262 220 1264
rect 222 1268 230 1270
rect 222 1264 224 1268
rect 228 1264 230 1268
rect 296 1268 298 1272
rect 302 1268 304 1272
rect 580 1270 588 1272
rect 296 1266 304 1268
rect 366 1268 374 1270
rect 366 1264 368 1268
rect 372 1264 374 1268
rect 222 1262 230 1264
rect 296 1262 304 1264
rect 366 1262 374 1264
rect 376 1268 384 1270
rect 376 1264 378 1268
rect 382 1264 384 1268
rect 376 1262 384 1264
rect 386 1268 394 1270
rect 386 1264 388 1268
rect 392 1264 394 1268
rect 386 1262 394 1264
rect 396 1268 404 1270
rect 396 1264 398 1268
rect 402 1264 404 1268
rect 396 1262 404 1264
rect 406 1268 414 1270
rect 406 1264 408 1268
rect 412 1264 414 1268
rect 406 1262 414 1264
rect 416 1268 424 1270
rect 416 1264 418 1268
rect 422 1264 424 1268
rect 416 1262 424 1264
rect 426 1268 434 1270
rect 426 1264 428 1268
rect 432 1264 434 1268
rect 426 1262 434 1264
rect 436 1268 444 1270
rect 436 1264 438 1268
rect 442 1264 444 1268
rect 436 1262 444 1264
rect 446 1268 454 1270
rect 446 1264 448 1268
rect 452 1264 454 1268
rect 446 1262 454 1264
rect 456 1268 464 1270
rect 456 1264 458 1268
rect 462 1264 464 1268
rect 456 1262 464 1264
rect 466 1268 474 1270
rect 466 1264 468 1268
rect 472 1264 474 1268
rect 466 1262 474 1264
rect 476 1268 484 1270
rect 476 1264 478 1268
rect 482 1264 484 1268
rect 476 1262 484 1264
rect 488 1268 496 1270
rect 488 1264 490 1268
rect 494 1264 496 1268
rect 488 1262 496 1264
rect 498 1268 506 1270
rect 498 1264 500 1268
rect 504 1264 506 1268
rect 498 1262 506 1264
rect 508 1268 516 1270
rect 508 1264 510 1268
rect 514 1264 516 1268
rect 508 1262 516 1264
rect 518 1268 526 1270
rect 518 1264 520 1268
rect 524 1264 526 1268
rect 518 1262 526 1264
rect 528 1268 536 1270
rect 528 1264 530 1268
rect 534 1264 536 1268
rect 528 1262 536 1264
rect 542 1268 550 1270
rect 542 1264 544 1268
rect 548 1264 550 1268
rect 542 1262 550 1264
rect 552 1268 560 1270
rect 552 1264 554 1268
rect 558 1264 560 1268
rect 552 1262 560 1264
rect 564 1268 572 1270
rect 564 1264 566 1268
rect 570 1264 572 1268
rect 580 1266 582 1270
rect 586 1266 588 1270
rect 580 1264 588 1266
rect 590 1270 598 1272
rect 590 1266 592 1270
rect 596 1266 598 1270
rect 590 1264 598 1266
rect 564 1262 572 1264
rect 28 1260 36 1262
rect 40 1258 48 1260
rect 12 1256 20 1258
rect 28 1256 36 1258
rect 2 1252 10 1254
rect 2 1248 4 1252
rect 8 1248 10 1252
rect 2 1246 10 1248
rect 12 1252 20 1254
rect 12 1248 14 1252
rect 18 1248 20 1252
rect 28 1252 30 1256
rect 34 1252 36 1256
rect 40 1254 42 1258
rect 46 1254 48 1258
rect 40 1252 48 1254
rect 50 1258 58 1260
rect 50 1254 52 1258
rect 56 1254 58 1258
rect 296 1258 298 1262
rect 302 1258 304 1262
rect 580 1260 588 1262
rect 296 1256 304 1258
rect 542 1258 550 1260
rect 542 1254 544 1258
rect 548 1254 550 1258
rect 50 1252 58 1254
rect 296 1252 304 1254
rect 542 1252 550 1254
rect 552 1258 560 1260
rect 552 1254 554 1258
rect 558 1254 560 1258
rect 552 1252 560 1254
rect 564 1258 572 1260
rect 564 1254 566 1258
rect 570 1254 572 1258
rect 580 1256 582 1260
rect 586 1256 588 1260
rect 580 1254 588 1256
rect 590 1260 598 1262
rect 590 1256 592 1260
rect 596 1256 598 1260
rect 590 1254 598 1256
rect 564 1252 572 1254
rect 28 1250 36 1252
rect 40 1248 48 1250
rect 12 1246 20 1248
rect 28 1246 36 1248
rect 2 1242 10 1244
rect 2 1238 4 1242
rect 8 1238 10 1242
rect 2 1236 10 1238
rect 12 1242 20 1244
rect 12 1238 14 1242
rect 18 1238 20 1242
rect 28 1242 30 1246
rect 34 1242 36 1246
rect 40 1244 42 1248
rect 46 1244 48 1248
rect 40 1242 48 1244
rect 50 1248 58 1250
rect 50 1244 52 1248
rect 56 1244 58 1248
rect 50 1242 58 1244
rect 64 1249 72 1251
rect 64 1245 66 1249
rect 70 1245 72 1249
rect 296 1248 298 1252
rect 302 1248 304 1252
rect 580 1250 588 1252
rect 296 1246 304 1248
rect 528 1248 536 1250
rect 64 1243 72 1245
rect 528 1244 530 1248
rect 534 1244 536 1248
rect 84 1242 92 1244
rect 28 1240 36 1242
rect 40 1238 48 1240
rect 12 1236 20 1238
rect 28 1236 36 1238
rect 2 1232 10 1234
rect 2 1228 4 1232
rect 8 1228 10 1232
rect 2 1226 10 1228
rect 12 1232 20 1234
rect 12 1228 14 1232
rect 18 1228 20 1232
rect 28 1232 30 1236
rect 34 1232 36 1236
rect 40 1234 42 1238
rect 46 1234 48 1238
rect 40 1232 48 1234
rect 50 1238 58 1240
rect 50 1234 52 1238
rect 56 1234 58 1238
rect 84 1238 86 1242
rect 90 1238 92 1242
rect 84 1236 92 1238
rect 94 1242 102 1244
rect 94 1238 96 1242
rect 100 1238 102 1242
rect 94 1236 102 1238
rect 104 1242 112 1244
rect 104 1238 106 1242
rect 110 1238 112 1242
rect 104 1236 112 1238
rect 114 1242 122 1244
rect 114 1238 116 1242
rect 120 1238 122 1242
rect 114 1236 122 1238
rect 124 1242 132 1244
rect 124 1238 126 1242
rect 130 1238 132 1242
rect 124 1236 132 1238
rect 134 1242 142 1244
rect 134 1238 136 1242
rect 140 1238 142 1242
rect 134 1236 142 1238
rect 144 1242 152 1244
rect 144 1238 146 1242
rect 150 1238 152 1242
rect 144 1236 152 1238
rect 154 1242 162 1244
rect 154 1238 156 1242
rect 160 1238 162 1242
rect 154 1236 162 1238
rect 164 1242 172 1244
rect 164 1238 166 1242
rect 170 1238 172 1242
rect 164 1236 172 1238
rect 174 1242 182 1244
rect 174 1238 176 1242
rect 180 1238 182 1242
rect 174 1236 182 1238
rect 184 1242 192 1244
rect 184 1238 186 1242
rect 190 1238 192 1242
rect 184 1236 192 1238
rect 194 1242 202 1244
rect 194 1238 196 1242
rect 200 1238 202 1242
rect 194 1236 202 1238
rect 204 1242 212 1244
rect 204 1238 206 1242
rect 210 1238 212 1242
rect 204 1236 212 1238
rect 214 1242 222 1244
rect 214 1238 216 1242
rect 220 1238 222 1242
rect 214 1236 222 1238
rect 224 1242 232 1244
rect 224 1238 226 1242
rect 230 1238 232 1242
rect 224 1236 232 1238
rect 296 1242 304 1244
rect 296 1238 298 1242
rect 302 1238 304 1242
rect 296 1236 304 1238
rect 368 1242 376 1244
rect 368 1238 370 1242
rect 374 1238 376 1242
rect 368 1236 376 1238
rect 378 1242 386 1244
rect 378 1238 380 1242
rect 384 1238 386 1242
rect 378 1236 386 1238
rect 388 1242 396 1244
rect 388 1238 390 1242
rect 394 1238 396 1242
rect 388 1236 396 1238
rect 398 1242 406 1244
rect 398 1238 400 1242
rect 404 1238 406 1242
rect 398 1236 406 1238
rect 408 1242 416 1244
rect 408 1238 410 1242
rect 414 1238 416 1242
rect 408 1236 416 1238
rect 418 1242 426 1244
rect 418 1238 420 1242
rect 424 1238 426 1242
rect 418 1236 426 1238
rect 428 1242 436 1244
rect 428 1238 430 1242
rect 434 1238 436 1242
rect 428 1236 436 1238
rect 438 1242 446 1244
rect 438 1238 440 1242
rect 444 1238 446 1242
rect 438 1236 446 1238
rect 448 1242 456 1244
rect 448 1238 450 1242
rect 454 1238 456 1242
rect 448 1236 456 1238
rect 458 1242 466 1244
rect 458 1238 460 1242
rect 464 1238 466 1242
rect 458 1236 466 1238
rect 468 1242 476 1244
rect 468 1238 470 1242
rect 474 1238 476 1242
rect 468 1236 476 1238
rect 478 1242 486 1244
rect 478 1238 480 1242
rect 484 1238 486 1242
rect 478 1236 486 1238
rect 488 1242 496 1244
rect 488 1238 490 1242
rect 494 1238 496 1242
rect 488 1236 496 1238
rect 498 1242 506 1244
rect 498 1238 500 1242
rect 504 1238 506 1242
rect 498 1236 506 1238
rect 508 1242 516 1244
rect 528 1242 536 1244
rect 542 1248 550 1250
rect 542 1244 544 1248
rect 548 1244 550 1248
rect 542 1242 550 1244
rect 552 1248 560 1250
rect 552 1244 554 1248
rect 558 1244 560 1248
rect 552 1242 560 1244
rect 564 1248 572 1250
rect 564 1244 566 1248
rect 570 1244 572 1248
rect 580 1246 582 1250
rect 586 1246 588 1250
rect 580 1244 588 1246
rect 590 1250 598 1252
rect 590 1246 592 1250
rect 596 1246 598 1250
rect 590 1244 598 1246
rect 564 1242 572 1244
rect 508 1238 510 1242
rect 514 1238 516 1242
rect 580 1240 588 1242
rect 508 1236 516 1238
rect 542 1238 550 1240
rect 542 1234 544 1238
rect 548 1234 550 1238
rect 50 1232 58 1234
rect 28 1230 36 1232
rect 82 1231 90 1233
rect 40 1228 48 1230
rect 12 1226 20 1228
rect 28 1226 36 1228
rect 2 1222 10 1224
rect 2 1218 4 1222
rect 8 1218 10 1222
rect 2 1216 10 1218
rect 12 1222 20 1224
rect 12 1218 14 1222
rect 18 1218 20 1222
rect 28 1222 30 1226
rect 34 1222 36 1226
rect 40 1224 42 1228
rect 46 1224 48 1228
rect 40 1222 48 1224
rect 50 1228 58 1230
rect 50 1224 52 1228
rect 56 1224 58 1228
rect 50 1222 58 1224
rect 64 1226 72 1228
rect 64 1222 66 1226
rect 70 1222 72 1226
rect 82 1227 84 1231
rect 88 1227 90 1231
rect 82 1225 90 1227
rect 92 1231 100 1233
rect 92 1227 94 1231
rect 98 1227 100 1231
rect 92 1225 100 1227
rect 296 1232 304 1234
rect 542 1232 550 1234
rect 552 1238 560 1240
rect 552 1234 554 1238
rect 558 1234 560 1238
rect 552 1232 560 1234
rect 564 1238 572 1240
rect 564 1234 566 1238
rect 570 1234 572 1238
rect 580 1236 582 1240
rect 586 1236 588 1240
rect 580 1234 588 1236
rect 590 1240 598 1242
rect 590 1236 592 1240
rect 596 1236 598 1240
rect 590 1234 598 1236
rect 564 1232 572 1234
rect 296 1228 298 1232
rect 302 1228 304 1232
rect 580 1230 588 1232
rect 296 1226 304 1228
rect 498 1227 506 1229
rect 28 1220 36 1222
rect 64 1220 72 1222
rect 82 1221 90 1223
rect 40 1218 48 1220
rect 12 1216 20 1218
rect 28 1216 36 1218
rect 2 1212 10 1214
rect 2 1208 4 1212
rect 8 1208 10 1212
rect 2 1206 10 1208
rect 12 1212 20 1214
rect 12 1208 14 1212
rect 18 1208 20 1212
rect 28 1212 30 1216
rect 34 1212 36 1216
rect 40 1214 42 1218
rect 46 1214 48 1218
rect 40 1212 48 1214
rect 50 1218 58 1220
rect 50 1214 52 1218
rect 56 1214 58 1218
rect 50 1212 58 1214
rect 64 1216 72 1218
rect 64 1212 66 1216
rect 70 1212 72 1216
rect 82 1217 84 1221
rect 88 1217 90 1221
rect 82 1215 90 1217
rect 92 1221 100 1223
rect 92 1217 94 1221
rect 98 1217 100 1221
rect 92 1215 100 1217
rect 296 1222 304 1224
rect 296 1218 298 1222
rect 302 1218 304 1222
rect 498 1223 500 1227
rect 504 1223 506 1227
rect 498 1221 506 1223
rect 508 1227 516 1229
rect 508 1223 510 1227
rect 514 1223 516 1227
rect 542 1228 550 1230
rect 508 1221 516 1223
rect 528 1223 536 1225
rect 528 1219 530 1223
rect 534 1219 536 1223
rect 542 1224 544 1228
rect 548 1224 550 1228
rect 542 1222 550 1224
rect 552 1228 560 1230
rect 552 1224 554 1228
rect 558 1224 560 1228
rect 552 1222 560 1224
rect 564 1228 572 1230
rect 564 1224 566 1228
rect 570 1224 572 1228
rect 580 1226 582 1230
rect 586 1226 588 1230
rect 580 1224 588 1226
rect 590 1230 598 1232
rect 590 1226 592 1230
rect 596 1226 598 1230
rect 590 1224 598 1226
rect 564 1222 572 1224
rect 580 1220 588 1222
rect 296 1216 304 1218
rect 498 1217 506 1219
rect 112 1214 120 1216
rect 28 1210 36 1212
rect 64 1210 72 1212
rect 82 1211 90 1213
rect 40 1208 48 1210
rect 12 1206 20 1208
rect 28 1206 36 1208
rect 2 1202 10 1204
rect 2 1198 4 1202
rect 8 1198 10 1202
rect 2 1196 10 1198
rect 12 1202 20 1204
rect 12 1198 14 1202
rect 18 1198 20 1202
rect 28 1202 30 1206
rect 34 1202 36 1206
rect 40 1204 42 1208
rect 46 1204 48 1208
rect 40 1202 48 1204
rect 50 1208 58 1210
rect 50 1204 52 1208
rect 56 1204 58 1208
rect 50 1202 58 1204
rect 64 1206 72 1208
rect 64 1202 66 1206
rect 70 1202 72 1206
rect 82 1207 84 1211
rect 88 1207 90 1211
rect 82 1205 90 1207
rect 92 1211 100 1213
rect 92 1207 94 1211
rect 98 1207 100 1211
rect 112 1210 114 1214
rect 118 1210 120 1214
rect 112 1208 120 1210
rect 122 1214 130 1216
rect 122 1210 124 1214
rect 128 1210 130 1214
rect 122 1208 130 1210
rect 132 1214 140 1216
rect 132 1210 134 1214
rect 138 1210 140 1214
rect 132 1208 140 1210
rect 142 1214 150 1216
rect 142 1210 144 1214
rect 148 1210 150 1214
rect 142 1208 150 1210
rect 152 1214 160 1216
rect 152 1210 154 1214
rect 158 1210 160 1214
rect 152 1208 160 1210
rect 162 1214 170 1216
rect 162 1210 164 1214
rect 168 1210 170 1214
rect 162 1208 170 1210
rect 172 1214 180 1216
rect 172 1210 174 1214
rect 178 1210 180 1214
rect 172 1208 180 1210
rect 182 1214 190 1216
rect 182 1210 184 1214
rect 188 1210 190 1214
rect 182 1208 190 1210
rect 192 1214 200 1216
rect 192 1210 194 1214
rect 198 1210 200 1214
rect 192 1208 200 1210
rect 202 1214 210 1216
rect 202 1210 204 1214
rect 208 1210 210 1214
rect 202 1208 210 1210
rect 212 1214 220 1216
rect 212 1210 214 1214
rect 218 1210 220 1214
rect 212 1208 220 1210
rect 222 1214 230 1216
rect 222 1210 224 1214
rect 228 1210 230 1214
rect 222 1208 230 1210
rect 232 1214 240 1216
rect 360 1214 368 1216
rect 232 1210 234 1214
rect 238 1210 240 1214
rect 232 1208 240 1210
rect 296 1212 304 1214
rect 296 1208 298 1212
rect 302 1208 304 1212
rect 360 1210 362 1214
rect 366 1210 368 1214
rect 360 1208 368 1210
rect 370 1214 378 1216
rect 370 1210 372 1214
rect 376 1210 378 1214
rect 370 1208 378 1210
rect 380 1214 388 1216
rect 380 1210 382 1214
rect 386 1210 388 1214
rect 380 1208 388 1210
rect 390 1214 398 1216
rect 390 1210 392 1214
rect 396 1210 398 1214
rect 390 1208 398 1210
rect 400 1214 408 1216
rect 400 1210 402 1214
rect 406 1210 408 1214
rect 400 1208 408 1210
rect 410 1214 418 1216
rect 410 1210 412 1214
rect 416 1210 418 1214
rect 410 1208 418 1210
rect 420 1214 428 1216
rect 420 1210 422 1214
rect 426 1210 428 1214
rect 420 1208 428 1210
rect 430 1214 438 1216
rect 430 1210 432 1214
rect 436 1210 438 1214
rect 430 1208 438 1210
rect 440 1214 448 1216
rect 440 1210 442 1214
rect 446 1210 448 1214
rect 440 1208 448 1210
rect 450 1214 458 1216
rect 450 1210 452 1214
rect 456 1210 458 1214
rect 450 1208 458 1210
rect 460 1214 468 1216
rect 460 1210 462 1214
rect 466 1210 468 1214
rect 460 1208 468 1210
rect 470 1214 478 1216
rect 470 1210 472 1214
rect 476 1210 478 1214
rect 470 1208 478 1210
rect 480 1214 488 1216
rect 480 1210 482 1214
rect 486 1210 488 1214
rect 498 1213 500 1217
rect 504 1213 506 1217
rect 498 1211 506 1213
rect 508 1217 516 1219
rect 528 1217 536 1219
rect 542 1218 550 1220
rect 508 1213 510 1217
rect 514 1213 516 1217
rect 508 1211 516 1213
rect 528 1213 536 1215
rect 480 1208 488 1210
rect 528 1209 530 1213
rect 534 1209 536 1213
rect 542 1214 544 1218
rect 548 1214 550 1218
rect 542 1212 550 1214
rect 552 1218 560 1220
rect 552 1214 554 1218
rect 558 1214 560 1218
rect 552 1212 560 1214
rect 564 1218 572 1220
rect 564 1214 566 1218
rect 570 1214 572 1218
rect 580 1216 582 1220
rect 586 1216 588 1220
rect 580 1214 588 1216
rect 590 1220 598 1222
rect 590 1216 592 1220
rect 596 1216 598 1220
rect 590 1214 598 1216
rect 564 1212 572 1214
rect 580 1210 588 1212
rect 92 1205 100 1207
rect 296 1206 304 1208
rect 498 1207 506 1209
rect 112 1204 120 1206
rect 28 1200 36 1202
rect 64 1200 72 1202
rect 82 1201 90 1203
rect 40 1198 48 1200
rect 12 1196 20 1198
rect 28 1196 36 1198
rect 2 1192 10 1194
rect 2 1188 4 1192
rect 8 1188 10 1192
rect 2 1186 10 1188
rect 12 1192 20 1194
rect 12 1188 14 1192
rect 18 1188 20 1192
rect 28 1192 30 1196
rect 34 1192 36 1196
rect 40 1194 42 1198
rect 46 1194 48 1198
rect 40 1192 48 1194
rect 50 1198 58 1200
rect 50 1194 52 1198
rect 56 1194 58 1198
rect 50 1192 58 1194
rect 64 1196 72 1198
rect 64 1192 66 1196
rect 70 1192 72 1196
rect 82 1197 84 1201
rect 88 1197 90 1201
rect 82 1195 90 1197
rect 92 1201 100 1203
rect 92 1197 94 1201
rect 98 1197 100 1201
rect 112 1200 114 1204
rect 118 1200 120 1204
rect 112 1198 120 1200
rect 122 1204 130 1206
rect 122 1200 124 1204
rect 128 1200 130 1204
rect 122 1198 130 1200
rect 132 1204 140 1206
rect 132 1200 134 1204
rect 138 1200 140 1204
rect 132 1198 140 1200
rect 142 1204 150 1206
rect 142 1200 144 1204
rect 148 1200 150 1204
rect 142 1198 150 1200
rect 152 1204 160 1206
rect 152 1200 154 1204
rect 158 1200 160 1204
rect 152 1198 160 1200
rect 162 1204 170 1206
rect 162 1200 164 1204
rect 168 1200 170 1204
rect 162 1198 170 1200
rect 172 1204 180 1206
rect 172 1200 174 1204
rect 178 1200 180 1204
rect 172 1198 180 1200
rect 182 1204 190 1206
rect 182 1200 184 1204
rect 188 1200 190 1204
rect 182 1198 190 1200
rect 192 1204 200 1206
rect 192 1200 194 1204
rect 198 1200 200 1204
rect 192 1198 200 1200
rect 202 1204 210 1206
rect 202 1200 204 1204
rect 208 1200 210 1204
rect 202 1198 210 1200
rect 212 1204 220 1206
rect 212 1200 214 1204
rect 218 1200 220 1204
rect 212 1198 220 1200
rect 222 1204 230 1206
rect 222 1200 224 1204
rect 228 1200 230 1204
rect 222 1198 230 1200
rect 232 1204 240 1206
rect 360 1204 368 1206
rect 232 1200 234 1204
rect 238 1200 240 1204
rect 232 1198 240 1200
rect 296 1202 304 1204
rect 296 1198 298 1202
rect 302 1198 304 1202
rect 360 1200 362 1204
rect 366 1200 368 1204
rect 360 1198 368 1200
rect 370 1204 378 1206
rect 370 1200 372 1204
rect 376 1200 378 1204
rect 370 1198 378 1200
rect 380 1204 388 1206
rect 380 1200 382 1204
rect 386 1200 388 1204
rect 380 1198 388 1200
rect 390 1204 398 1206
rect 390 1200 392 1204
rect 396 1200 398 1204
rect 390 1198 398 1200
rect 400 1204 408 1206
rect 400 1200 402 1204
rect 406 1200 408 1204
rect 400 1198 408 1200
rect 410 1204 418 1206
rect 410 1200 412 1204
rect 416 1200 418 1204
rect 410 1198 418 1200
rect 420 1204 428 1206
rect 420 1200 422 1204
rect 426 1200 428 1204
rect 420 1198 428 1200
rect 430 1204 438 1206
rect 430 1200 432 1204
rect 436 1200 438 1204
rect 430 1198 438 1200
rect 440 1204 448 1206
rect 440 1200 442 1204
rect 446 1200 448 1204
rect 440 1198 448 1200
rect 450 1204 458 1206
rect 450 1200 452 1204
rect 456 1200 458 1204
rect 450 1198 458 1200
rect 460 1204 468 1206
rect 460 1200 462 1204
rect 466 1200 468 1204
rect 460 1198 468 1200
rect 470 1204 478 1206
rect 470 1200 472 1204
rect 476 1200 478 1204
rect 470 1198 478 1200
rect 480 1204 488 1206
rect 480 1200 482 1204
rect 486 1200 488 1204
rect 498 1203 500 1207
rect 504 1203 506 1207
rect 498 1201 506 1203
rect 508 1207 516 1209
rect 528 1207 536 1209
rect 542 1208 550 1210
rect 508 1203 510 1207
rect 514 1203 516 1207
rect 508 1201 516 1203
rect 528 1203 536 1205
rect 480 1198 488 1200
rect 528 1199 530 1203
rect 534 1199 536 1203
rect 542 1204 544 1208
rect 548 1204 550 1208
rect 542 1202 550 1204
rect 552 1208 560 1210
rect 552 1204 554 1208
rect 558 1204 560 1208
rect 552 1202 560 1204
rect 564 1208 572 1210
rect 564 1204 566 1208
rect 570 1204 572 1208
rect 580 1206 582 1210
rect 586 1206 588 1210
rect 580 1204 588 1206
rect 590 1210 598 1212
rect 590 1206 592 1210
rect 596 1206 598 1210
rect 590 1204 598 1206
rect 564 1202 572 1204
rect 580 1200 588 1202
rect 92 1195 100 1197
rect 296 1196 304 1198
rect 498 1197 506 1199
rect 28 1190 36 1192
rect 64 1190 72 1192
rect 82 1191 90 1193
rect 40 1188 48 1190
rect 12 1186 20 1188
rect 28 1186 36 1188
rect 2 1182 10 1184
rect 2 1178 4 1182
rect 8 1178 10 1182
rect 2 1176 10 1178
rect 12 1182 20 1184
rect 12 1178 14 1182
rect 18 1178 20 1182
rect 28 1182 30 1186
rect 34 1182 36 1186
rect 40 1184 42 1188
rect 46 1184 48 1188
rect 40 1182 48 1184
rect 50 1188 58 1190
rect 50 1184 52 1188
rect 56 1184 58 1188
rect 82 1187 84 1191
rect 88 1187 90 1191
rect 82 1185 90 1187
rect 92 1191 100 1193
rect 92 1187 94 1191
rect 98 1187 100 1191
rect 92 1185 100 1187
rect 296 1192 304 1194
rect 296 1188 298 1192
rect 302 1188 304 1192
rect 498 1193 500 1197
rect 504 1193 506 1197
rect 498 1191 506 1193
rect 508 1197 516 1199
rect 528 1197 536 1199
rect 542 1198 550 1200
rect 508 1193 510 1197
rect 514 1193 516 1197
rect 508 1191 516 1193
rect 528 1193 536 1195
rect 528 1189 530 1193
rect 534 1189 536 1193
rect 542 1194 544 1198
rect 548 1194 550 1198
rect 542 1192 550 1194
rect 552 1198 560 1200
rect 552 1194 554 1198
rect 558 1194 560 1198
rect 552 1192 560 1194
rect 564 1198 572 1200
rect 564 1194 566 1198
rect 570 1194 572 1198
rect 580 1196 582 1200
rect 586 1196 588 1200
rect 580 1194 588 1196
rect 590 1200 598 1202
rect 590 1196 592 1200
rect 596 1196 598 1200
rect 590 1194 598 1196
rect 564 1192 572 1194
rect 580 1190 588 1192
rect 296 1186 304 1188
rect 498 1187 506 1189
rect 50 1182 58 1184
rect 296 1182 304 1184
rect 28 1180 36 1182
rect 40 1178 48 1180
rect 12 1176 20 1178
rect 28 1176 36 1178
rect 2 1172 10 1174
rect 2 1168 4 1172
rect 8 1168 10 1172
rect 2 1166 10 1168
rect 12 1172 20 1174
rect 12 1168 14 1172
rect 18 1168 20 1172
rect 28 1172 30 1176
rect 34 1172 36 1176
rect 40 1174 42 1178
rect 46 1174 48 1178
rect 40 1172 48 1174
rect 50 1178 58 1180
rect 50 1174 52 1178
rect 56 1174 58 1178
rect 50 1172 58 1174
rect 64 1177 72 1179
rect 64 1173 66 1177
rect 70 1173 72 1177
rect 28 1170 36 1172
rect 64 1171 72 1173
rect 84 1178 92 1180
rect 84 1174 86 1178
rect 90 1174 92 1178
rect 84 1172 92 1174
rect 94 1178 102 1180
rect 94 1174 96 1178
rect 100 1174 102 1178
rect 94 1172 102 1174
rect 104 1178 112 1180
rect 104 1174 106 1178
rect 110 1174 112 1178
rect 104 1172 112 1174
rect 114 1178 122 1180
rect 114 1174 116 1178
rect 120 1174 122 1178
rect 114 1172 122 1174
rect 124 1178 132 1180
rect 124 1174 126 1178
rect 130 1174 132 1178
rect 124 1172 132 1174
rect 134 1178 142 1180
rect 134 1174 136 1178
rect 140 1174 142 1178
rect 134 1172 142 1174
rect 144 1178 152 1180
rect 144 1174 146 1178
rect 150 1174 152 1178
rect 144 1172 152 1174
rect 154 1178 162 1180
rect 154 1174 156 1178
rect 160 1174 162 1178
rect 154 1172 162 1174
rect 164 1178 172 1180
rect 164 1174 166 1178
rect 170 1174 172 1178
rect 164 1172 172 1174
rect 174 1178 182 1180
rect 174 1174 176 1178
rect 180 1174 182 1178
rect 174 1172 182 1174
rect 184 1178 192 1180
rect 184 1174 186 1178
rect 190 1174 192 1178
rect 184 1172 192 1174
rect 194 1178 202 1180
rect 194 1174 196 1178
rect 200 1174 202 1178
rect 194 1172 202 1174
rect 204 1178 212 1180
rect 204 1174 206 1178
rect 210 1174 212 1178
rect 204 1172 212 1174
rect 214 1178 222 1180
rect 214 1174 216 1178
rect 220 1174 222 1178
rect 214 1172 222 1174
rect 224 1178 232 1180
rect 224 1174 226 1178
rect 230 1174 232 1178
rect 296 1178 298 1182
rect 302 1178 304 1182
rect 498 1183 500 1187
rect 504 1183 506 1187
rect 498 1181 506 1183
rect 508 1187 516 1189
rect 528 1187 536 1189
rect 542 1188 550 1190
rect 508 1183 510 1187
rect 514 1183 516 1187
rect 508 1181 516 1183
rect 542 1184 544 1188
rect 548 1184 550 1188
rect 542 1182 550 1184
rect 552 1188 560 1190
rect 552 1184 554 1188
rect 558 1184 560 1188
rect 552 1182 560 1184
rect 564 1188 572 1190
rect 564 1184 566 1188
rect 570 1184 572 1188
rect 580 1186 582 1190
rect 586 1186 588 1190
rect 580 1184 588 1186
rect 590 1190 598 1192
rect 590 1186 592 1190
rect 596 1186 598 1190
rect 590 1184 598 1186
rect 564 1182 572 1184
rect 580 1180 588 1182
rect 542 1178 550 1180
rect 296 1176 304 1178
rect 368 1176 376 1178
rect 224 1172 232 1174
rect 296 1172 304 1174
rect 40 1168 48 1170
rect 12 1166 20 1168
rect 28 1166 36 1168
rect 2 1162 10 1164
rect 2 1158 4 1162
rect 8 1158 10 1162
rect 2 1156 10 1158
rect 12 1162 20 1164
rect 12 1158 14 1162
rect 18 1158 20 1162
rect 28 1162 30 1166
rect 34 1162 36 1166
rect 40 1164 42 1168
rect 46 1164 48 1168
rect 40 1162 48 1164
rect 50 1168 58 1170
rect 50 1164 52 1168
rect 56 1164 58 1168
rect 50 1162 58 1164
rect 64 1167 72 1169
rect 64 1163 66 1167
rect 70 1163 72 1167
rect 296 1168 298 1172
rect 302 1168 304 1172
rect 368 1172 370 1176
rect 374 1172 376 1176
rect 368 1170 376 1172
rect 378 1176 386 1178
rect 378 1172 380 1176
rect 384 1172 386 1176
rect 378 1170 386 1172
rect 388 1176 396 1178
rect 388 1172 390 1176
rect 394 1172 396 1176
rect 388 1170 396 1172
rect 398 1176 406 1178
rect 398 1172 400 1176
rect 404 1172 406 1176
rect 398 1170 406 1172
rect 408 1176 416 1178
rect 408 1172 410 1176
rect 414 1172 416 1176
rect 408 1170 416 1172
rect 418 1176 426 1178
rect 418 1172 420 1176
rect 424 1172 426 1176
rect 418 1170 426 1172
rect 428 1176 436 1178
rect 428 1172 430 1176
rect 434 1172 436 1176
rect 428 1170 436 1172
rect 438 1176 446 1178
rect 438 1172 440 1176
rect 444 1172 446 1176
rect 438 1170 446 1172
rect 448 1176 456 1178
rect 448 1172 450 1176
rect 454 1172 456 1176
rect 448 1170 456 1172
rect 458 1176 466 1178
rect 458 1172 460 1176
rect 464 1172 466 1176
rect 458 1170 466 1172
rect 468 1176 476 1178
rect 468 1172 470 1176
rect 474 1172 476 1176
rect 468 1170 476 1172
rect 478 1176 486 1178
rect 478 1172 480 1176
rect 484 1172 486 1176
rect 478 1170 486 1172
rect 488 1176 496 1178
rect 488 1172 490 1176
rect 494 1172 496 1176
rect 488 1170 496 1172
rect 498 1176 506 1178
rect 498 1172 500 1176
rect 504 1172 506 1176
rect 498 1170 506 1172
rect 508 1176 516 1178
rect 508 1172 510 1176
rect 514 1172 516 1176
rect 508 1170 516 1172
rect 528 1174 536 1176
rect 528 1170 530 1174
rect 534 1170 536 1174
rect 542 1174 544 1178
rect 548 1174 550 1178
rect 542 1172 550 1174
rect 552 1178 560 1180
rect 552 1174 554 1178
rect 558 1174 560 1178
rect 552 1172 560 1174
rect 564 1178 572 1180
rect 564 1174 566 1178
rect 570 1174 572 1178
rect 580 1176 582 1180
rect 586 1176 588 1180
rect 580 1174 588 1176
rect 590 1180 598 1182
rect 590 1176 592 1180
rect 596 1176 598 1180
rect 590 1174 598 1176
rect 564 1172 572 1174
rect 580 1170 588 1172
rect 528 1168 536 1170
rect 542 1168 550 1170
rect 296 1166 304 1168
rect 528 1164 536 1166
rect 28 1160 36 1162
rect 64 1161 72 1163
rect 296 1162 304 1164
rect 40 1158 48 1160
rect 12 1156 20 1158
rect 28 1156 36 1158
rect 2 1152 10 1154
rect 2 1148 4 1152
rect 8 1148 10 1152
rect 2 1146 10 1148
rect 12 1152 20 1154
rect 12 1148 14 1152
rect 18 1148 20 1152
rect 28 1152 30 1156
rect 34 1152 36 1156
rect 40 1154 42 1158
rect 46 1154 48 1158
rect 40 1152 48 1154
rect 50 1158 58 1160
rect 50 1154 52 1158
rect 56 1154 58 1158
rect 50 1152 58 1154
rect 64 1157 72 1159
rect 64 1153 66 1157
rect 70 1153 72 1157
rect 296 1158 298 1162
rect 302 1158 304 1162
rect 528 1160 530 1164
rect 534 1160 536 1164
rect 542 1164 544 1168
rect 548 1164 550 1168
rect 542 1162 550 1164
rect 552 1168 560 1170
rect 552 1164 554 1168
rect 558 1164 560 1168
rect 552 1162 560 1164
rect 564 1168 572 1170
rect 564 1164 566 1168
rect 570 1164 572 1168
rect 580 1166 582 1170
rect 586 1166 588 1170
rect 580 1164 588 1166
rect 590 1170 598 1172
rect 590 1166 592 1170
rect 596 1166 598 1170
rect 590 1164 598 1166
rect 564 1162 572 1164
rect 580 1160 588 1162
rect 528 1158 536 1160
rect 542 1158 550 1160
rect 296 1156 304 1158
rect 528 1154 536 1156
rect 28 1150 36 1152
rect 64 1151 72 1153
rect 296 1152 304 1154
rect 83 1150 91 1152
rect 40 1148 48 1150
rect 12 1146 20 1148
rect 28 1146 36 1148
rect 2 1142 10 1144
rect 2 1138 4 1142
rect 8 1138 10 1142
rect 2 1136 10 1138
rect 12 1142 20 1144
rect 12 1138 14 1142
rect 18 1138 20 1142
rect 28 1142 30 1146
rect 34 1142 36 1146
rect 40 1144 42 1148
rect 46 1144 48 1148
rect 40 1142 48 1144
rect 50 1148 58 1150
rect 50 1144 52 1148
rect 56 1144 58 1148
rect 50 1142 58 1144
rect 64 1147 72 1149
rect 64 1143 66 1147
rect 70 1143 72 1147
rect 83 1146 85 1150
rect 89 1146 91 1150
rect 83 1144 91 1146
rect 93 1150 101 1152
rect 93 1146 95 1150
rect 99 1146 101 1150
rect 93 1144 101 1146
rect 103 1150 111 1152
rect 103 1146 105 1150
rect 109 1146 111 1150
rect 103 1144 111 1146
rect 113 1150 121 1152
rect 113 1146 115 1150
rect 119 1146 121 1150
rect 113 1144 121 1146
rect 123 1150 131 1152
rect 123 1146 125 1150
rect 129 1146 131 1150
rect 123 1144 131 1146
rect 133 1150 141 1152
rect 133 1146 135 1150
rect 139 1146 141 1150
rect 133 1144 141 1146
rect 143 1150 151 1152
rect 143 1146 145 1150
rect 149 1146 151 1150
rect 143 1144 151 1146
rect 153 1150 161 1152
rect 153 1146 155 1150
rect 159 1146 161 1150
rect 153 1144 161 1146
rect 163 1150 171 1152
rect 163 1146 165 1150
rect 169 1146 171 1150
rect 163 1144 171 1146
rect 173 1150 181 1152
rect 173 1146 175 1150
rect 179 1146 181 1150
rect 173 1144 181 1146
rect 183 1150 191 1152
rect 183 1146 185 1150
rect 189 1146 191 1150
rect 183 1144 191 1146
rect 193 1150 201 1152
rect 193 1146 195 1150
rect 199 1146 201 1150
rect 193 1144 201 1146
rect 203 1150 211 1152
rect 203 1146 205 1150
rect 209 1146 211 1150
rect 203 1144 211 1146
rect 213 1150 221 1152
rect 213 1146 215 1150
rect 219 1146 221 1150
rect 213 1144 221 1146
rect 223 1150 231 1152
rect 223 1146 225 1150
rect 229 1146 231 1150
rect 296 1148 298 1152
rect 302 1148 304 1152
rect 296 1146 304 1148
rect 368 1150 376 1152
rect 368 1146 370 1150
rect 374 1146 376 1150
rect 223 1144 231 1146
rect 368 1144 376 1146
rect 378 1150 386 1152
rect 378 1146 380 1150
rect 384 1146 386 1150
rect 378 1144 386 1146
rect 388 1150 396 1152
rect 388 1146 390 1150
rect 394 1146 396 1150
rect 388 1144 396 1146
rect 398 1150 406 1152
rect 398 1146 400 1150
rect 404 1146 406 1150
rect 398 1144 406 1146
rect 408 1150 416 1152
rect 408 1146 410 1150
rect 414 1146 416 1150
rect 408 1144 416 1146
rect 418 1150 426 1152
rect 418 1146 420 1150
rect 424 1146 426 1150
rect 418 1144 426 1146
rect 428 1150 436 1152
rect 428 1146 430 1150
rect 434 1146 436 1150
rect 428 1144 436 1146
rect 438 1150 446 1152
rect 438 1146 440 1150
rect 444 1146 446 1150
rect 438 1144 446 1146
rect 448 1150 456 1152
rect 448 1146 450 1150
rect 454 1146 456 1150
rect 448 1144 456 1146
rect 458 1150 466 1152
rect 458 1146 460 1150
rect 464 1146 466 1150
rect 458 1144 466 1146
rect 468 1150 476 1152
rect 468 1146 470 1150
rect 474 1146 476 1150
rect 468 1144 476 1146
rect 478 1150 486 1152
rect 478 1146 480 1150
rect 484 1146 486 1150
rect 478 1144 486 1146
rect 488 1150 496 1152
rect 488 1146 490 1150
rect 494 1146 496 1150
rect 488 1144 496 1146
rect 498 1150 506 1152
rect 498 1146 500 1150
rect 504 1146 506 1150
rect 498 1144 506 1146
rect 508 1150 516 1152
rect 508 1146 510 1150
rect 514 1146 516 1150
rect 528 1150 530 1154
rect 534 1150 536 1154
rect 542 1154 544 1158
rect 548 1154 550 1158
rect 542 1152 550 1154
rect 552 1158 560 1160
rect 552 1154 554 1158
rect 558 1154 560 1158
rect 552 1152 560 1154
rect 564 1158 572 1160
rect 564 1154 566 1158
rect 570 1154 572 1158
rect 580 1156 582 1160
rect 586 1156 588 1160
rect 580 1154 588 1156
rect 590 1160 598 1162
rect 590 1156 592 1160
rect 596 1156 598 1160
rect 590 1154 598 1156
rect 564 1152 572 1154
rect 580 1150 588 1152
rect 528 1148 536 1150
rect 542 1148 550 1150
rect 508 1144 516 1146
rect 528 1144 536 1146
rect 28 1140 36 1142
rect 64 1141 72 1143
rect 296 1142 304 1144
rect 40 1138 48 1140
rect 12 1136 20 1138
rect 28 1136 36 1138
rect 2 1132 10 1134
rect 2 1128 4 1132
rect 8 1128 10 1132
rect 2 1126 10 1128
rect 12 1132 20 1134
rect 12 1128 14 1132
rect 18 1128 20 1132
rect 28 1132 30 1136
rect 34 1132 36 1136
rect 40 1134 42 1138
rect 46 1134 48 1138
rect 40 1132 48 1134
rect 50 1138 58 1140
rect 50 1134 52 1138
rect 56 1134 58 1138
rect 50 1132 58 1134
rect 64 1137 72 1139
rect 64 1133 66 1137
rect 70 1133 72 1137
rect 28 1130 36 1132
rect 64 1131 72 1133
rect 83 1138 91 1140
rect 83 1134 85 1138
rect 89 1134 91 1138
rect 83 1132 91 1134
rect 93 1138 101 1140
rect 93 1134 95 1138
rect 99 1134 101 1138
rect 93 1132 101 1134
rect 103 1138 111 1140
rect 103 1134 105 1138
rect 109 1134 111 1138
rect 103 1132 111 1134
rect 113 1138 121 1140
rect 113 1134 115 1138
rect 119 1134 121 1138
rect 113 1132 121 1134
rect 123 1138 131 1140
rect 123 1134 125 1138
rect 129 1134 131 1138
rect 123 1132 131 1134
rect 133 1138 141 1140
rect 133 1134 135 1138
rect 139 1134 141 1138
rect 133 1132 141 1134
rect 143 1138 151 1140
rect 143 1134 145 1138
rect 149 1134 151 1138
rect 143 1132 151 1134
rect 153 1138 161 1140
rect 153 1134 155 1138
rect 159 1134 161 1138
rect 153 1132 161 1134
rect 163 1138 171 1140
rect 163 1134 165 1138
rect 169 1134 171 1138
rect 163 1132 171 1134
rect 173 1138 181 1140
rect 173 1134 175 1138
rect 179 1134 181 1138
rect 173 1132 181 1134
rect 183 1138 191 1140
rect 183 1134 185 1138
rect 189 1134 191 1138
rect 183 1132 191 1134
rect 193 1138 201 1140
rect 193 1134 195 1138
rect 199 1134 201 1138
rect 193 1132 201 1134
rect 203 1138 211 1140
rect 203 1134 205 1138
rect 209 1134 211 1138
rect 203 1132 211 1134
rect 213 1138 221 1140
rect 213 1134 215 1138
rect 219 1134 221 1138
rect 213 1132 221 1134
rect 223 1138 231 1140
rect 223 1134 225 1138
rect 229 1134 231 1138
rect 296 1138 298 1142
rect 302 1138 304 1142
rect 528 1140 530 1144
rect 534 1140 536 1144
rect 542 1144 544 1148
rect 548 1144 550 1148
rect 542 1142 550 1144
rect 552 1148 560 1150
rect 552 1144 554 1148
rect 558 1144 560 1148
rect 552 1142 560 1144
rect 564 1148 572 1150
rect 564 1144 566 1148
rect 570 1144 572 1148
rect 580 1146 582 1150
rect 586 1146 588 1150
rect 580 1144 588 1146
rect 590 1150 598 1152
rect 590 1146 592 1150
rect 596 1146 598 1150
rect 590 1144 598 1146
rect 564 1142 572 1144
rect 580 1140 588 1142
rect 296 1136 304 1138
rect 368 1138 376 1140
rect 368 1134 370 1138
rect 374 1134 376 1138
rect 223 1132 231 1134
rect 296 1132 304 1134
rect 368 1132 376 1134
rect 378 1138 386 1140
rect 378 1134 380 1138
rect 384 1134 386 1138
rect 378 1132 386 1134
rect 388 1138 396 1140
rect 388 1134 390 1138
rect 394 1134 396 1138
rect 388 1132 396 1134
rect 398 1138 406 1140
rect 398 1134 400 1138
rect 404 1134 406 1138
rect 398 1132 406 1134
rect 408 1138 416 1140
rect 408 1134 410 1138
rect 414 1134 416 1138
rect 408 1132 416 1134
rect 418 1138 426 1140
rect 418 1134 420 1138
rect 424 1134 426 1138
rect 418 1132 426 1134
rect 428 1138 436 1140
rect 428 1134 430 1138
rect 434 1134 436 1138
rect 428 1132 436 1134
rect 438 1138 446 1140
rect 438 1134 440 1138
rect 444 1134 446 1138
rect 438 1132 446 1134
rect 448 1138 456 1140
rect 448 1134 450 1138
rect 454 1134 456 1138
rect 448 1132 456 1134
rect 458 1138 466 1140
rect 458 1134 460 1138
rect 464 1134 466 1138
rect 458 1132 466 1134
rect 468 1138 476 1140
rect 468 1134 470 1138
rect 474 1134 476 1138
rect 468 1132 476 1134
rect 478 1138 486 1140
rect 478 1134 480 1138
rect 484 1134 486 1138
rect 478 1132 486 1134
rect 488 1138 496 1140
rect 488 1134 490 1138
rect 494 1134 496 1138
rect 488 1132 496 1134
rect 498 1138 506 1140
rect 498 1134 500 1138
rect 504 1134 506 1138
rect 498 1132 506 1134
rect 508 1138 516 1140
rect 528 1138 536 1140
rect 542 1138 550 1140
rect 508 1134 510 1138
rect 514 1134 516 1138
rect 508 1132 516 1134
rect 528 1134 536 1136
rect 40 1128 48 1130
rect 12 1126 20 1128
rect 28 1126 36 1128
rect 2 1122 10 1124
rect 2 1118 4 1122
rect 8 1118 10 1122
rect 2 1116 10 1118
rect 12 1122 20 1124
rect 12 1118 14 1122
rect 18 1118 20 1122
rect 28 1122 30 1126
rect 34 1122 36 1126
rect 40 1124 42 1128
rect 46 1124 48 1128
rect 40 1122 48 1124
rect 50 1128 58 1130
rect 50 1124 52 1128
rect 56 1124 58 1128
rect 50 1122 58 1124
rect 64 1127 72 1129
rect 64 1123 66 1127
rect 70 1123 72 1127
rect 296 1128 298 1132
rect 302 1128 304 1132
rect 528 1130 530 1134
rect 534 1130 536 1134
rect 542 1134 544 1138
rect 548 1134 550 1138
rect 542 1132 550 1134
rect 552 1138 560 1140
rect 552 1134 554 1138
rect 558 1134 560 1138
rect 552 1132 560 1134
rect 564 1138 572 1140
rect 564 1134 566 1138
rect 570 1134 572 1138
rect 580 1136 582 1140
rect 586 1136 588 1140
rect 580 1134 588 1136
rect 590 1140 598 1142
rect 590 1136 592 1140
rect 596 1136 598 1140
rect 590 1134 598 1136
rect 564 1132 572 1134
rect 580 1130 588 1132
rect 528 1128 536 1130
rect 542 1128 550 1130
rect 296 1126 304 1128
rect 528 1124 536 1126
rect 28 1120 36 1122
rect 64 1121 72 1123
rect 296 1122 304 1124
rect 40 1118 48 1120
rect 12 1116 20 1118
rect 28 1116 36 1118
rect 2 1112 10 1114
rect 2 1108 4 1112
rect 8 1108 10 1112
rect 2 1106 10 1108
rect 12 1112 20 1114
rect 12 1108 14 1112
rect 18 1108 20 1112
rect 28 1112 30 1116
rect 34 1112 36 1116
rect 40 1114 42 1118
rect 46 1114 48 1118
rect 40 1112 48 1114
rect 50 1118 58 1120
rect 50 1114 52 1118
rect 56 1114 58 1118
rect 50 1112 58 1114
rect 64 1117 72 1119
rect 64 1113 66 1117
rect 70 1113 72 1117
rect 296 1118 298 1122
rect 302 1118 304 1122
rect 528 1120 530 1124
rect 534 1120 536 1124
rect 542 1124 544 1128
rect 548 1124 550 1128
rect 542 1122 550 1124
rect 552 1128 560 1130
rect 552 1124 554 1128
rect 558 1124 560 1128
rect 552 1122 560 1124
rect 564 1128 572 1130
rect 564 1124 566 1128
rect 570 1124 572 1128
rect 580 1126 582 1130
rect 586 1126 588 1130
rect 580 1124 588 1126
rect 590 1130 598 1132
rect 590 1126 592 1130
rect 596 1126 598 1130
rect 590 1124 598 1126
rect 564 1122 572 1124
rect 580 1120 588 1122
rect 528 1118 536 1120
rect 542 1118 550 1120
rect 296 1116 304 1118
rect 528 1114 536 1116
rect 28 1110 36 1112
rect 64 1111 72 1113
rect 84 1111 92 1113
rect 40 1108 48 1110
rect 12 1106 20 1108
rect 28 1106 36 1108
rect 2 1102 10 1104
rect 2 1098 4 1102
rect 8 1098 10 1102
rect 2 1096 10 1098
rect 12 1102 20 1104
rect 12 1098 14 1102
rect 18 1098 20 1102
rect 28 1102 30 1106
rect 34 1102 36 1106
rect 40 1104 42 1108
rect 46 1104 48 1108
rect 40 1102 48 1104
rect 50 1108 58 1110
rect 50 1104 52 1108
rect 56 1104 58 1108
rect 84 1107 86 1111
rect 90 1107 92 1111
rect 84 1105 92 1107
rect 94 1111 102 1113
rect 94 1107 96 1111
rect 100 1107 102 1111
rect 94 1105 102 1107
rect 104 1111 112 1113
rect 104 1107 106 1111
rect 110 1107 112 1111
rect 104 1105 112 1107
rect 114 1111 122 1113
rect 114 1107 116 1111
rect 120 1107 122 1111
rect 114 1105 122 1107
rect 124 1111 132 1113
rect 124 1107 126 1111
rect 130 1107 132 1111
rect 124 1105 132 1107
rect 134 1111 142 1113
rect 134 1107 136 1111
rect 140 1107 142 1111
rect 134 1105 142 1107
rect 144 1111 152 1113
rect 144 1107 146 1111
rect 150 1107 152 1111
rect 144 1105 152 1107
rect 154 1111 162 1113
rect 154 1107 156 1111
rect 160 1107 162 1111
rect 154 1105 162 1107
rect 164 1111 172 1113
rect 164 1107 166 1111
rect 170 1107 172 1111
rect 164 1105 172 1107
rect 174 1111 182 1113
rect 174 1107 176 1111
rect 180 1107 182 1111
rect 174 1105 182 1107
rect 184 1111 192 1113
rect 184 1107 186 1111
rect 190 1107 192 1111
rect 184 1105 192 1107
rect 194 1111 202 1113
rect 194 1107 196 1111
rect 200 1107 202 1111
rect 194 1105 202 1107
rect 204 1111 212 1113
rect 204 1107 206 1111
rect 210 1107 212 1111
rect 204 1105 212 1107
rect 214 1111 222 1113
rect 214 1107 216 1111
rect 220 1107 222 1111
rect 214 1105 222 1107
rect 224 1111 232 1113
rect 224 1107 226 1111
rect 230 1107 232 1111
rect 224 1105 232 1107
rect 296 1112 304 1114
rect 296 1108 298 1112
rect 302 1108 304 1112
rect 296 1106 304 1108
rect 368 1112 376 1114
rect 368 1108 370 1112
rect 374 1108 376 1112
rect 368 1106 376 1108
rect 378 1112 386 1114
rect 378 1108 380 1112
rect 384 1108 386 1112
rect 378 1106 386 1108
rect 388 1112 396 1114
rect 388 1108 390 1112
rect 394 1108 396 1112
rect 388 1106 396 1108
rect 398 1112 406 1114
rect 398 1108 400 1112
rect 404 1108 406 1112
rect 398 1106 406 1108
rect 408 1112 416 1114
rect 408 1108 410 1112
rect 414 1108 416 1112
rect 408 1106 416 1108
rect 418 1112 426 1114
rect 418 1108 420 1112
rect 424 1108 426 1112
rect 418 1106 426 1108
rect 428 1112 436 1114
rect 428 1108 430 1112
rect 434 1108 436 1112
rect 428 1106 436 1108
rect 438 1112 446 1114
rect 438 1108 440 1112
rect 444 1108 446 1112
rect 438 1106 446 1108
rect 448 1112 456 1114
rect 448 1108 450 1112
rect 454 1108 456 1112
rect 448 1106 456 1108
rect 458 1112 466 1114
rect 458 1108 460 1112
rect 464 1108 466 1112
rect 458 1106 466 1108
rect 468 1112 476 1114
rect 468 1108 470 1112
rect 474 1108 476 1112
rect 468 1106 476 1108
rect 478 1112 486 1114
rect 478 1108 480 1112
rect 484 1108 486 1112
rect 478 1106 486 1108
rect 488 1112 496 1114
rect 488 1108 490 1112
rect 494 1108 496 1112
rect 488 1106 496 1108
rect 498 1112 506 1114
rect 498 1108 500 1112
rect 504 1108 506 1112
rect 498 1106 506 1108
rect 508 1112 516 1114
rect 508 1108 510 1112
rect 514 1108 516 1112
rect 528 1110 530 1114
rect 534 1110 536 1114
rect 542 1114 544 1118
rect 548 1114 550 1118
rect 542 1112 550 1114
rect 552 1118 560 1120
rect 552 1114 554 1118
rect 558 1114 560 1118
rect 552 1112 560 1114
rect 564 1118 572 1120
rect 564 1114 566 1118
rect 570 1114 572 1118
rect 580 1116 582 1120
rect 586 1116 588 1120
rect 580 1114 588 1116
rect 590 1120 598 1122
rect 590 1116 592 1120
rect 596 1116 598 1120
rect 590 1114 598 1116
rect 564 1112 572 1114
rect 580 1110 588 1112
rect 528 1108 536 1110
rect 542 1108 550 1110
rect 508 1106 516 1108
rect 542 1104 544 1108
rect 548 1104 550 1108
rect 50 1102 58 1104
rect 28 1100 36 1102
rect 84 1101 92 1103
rect 40 1098 48 1100
rect 12 1096 20 1098
rect 28 1096 36 1098
rect 2 1092 10 1094
rect 2 1088 4 1092
rect 8 1088 10 1092
rect 2 1086 10 1088
rect 12 1092 20 1094
rect 12 1088 14 1092
rect 18 1088 20 1092
rect 28 1092 30 1096
rect 34 1092 36 1096
rect 40 1094 42 1098
rect 46 1094 48 1098
rect 40 1092 48 1094
rect 50 1098 58 1100
rect 50 1094 52 1098
rect 56 1094 58 1098
rect 50 1092 58 1094
rect 64 1096 72 1098
rect 64 1092 66 1096
rect 70 1092 72 1096
rect 84 1097 86 1101
rect 90 1097 92 1101
rect 84 1095 92 1097
rect 94 1101 102 1103
rect 94 1097 96 1101
rect 100 1097 102 1101
rect 94 1095 102 1097
rect 296 1102 304 1104
rect 296 1098 298 1102
rect 302 1098 304 1102
rect 296 1096 304 1098
rect 498 1101 506 1103
rect 498 1097 500 1101
rect 504 1097 506 1101
rect 498 1095 506 1097
rect 508 1101 516 1103
rect 542 1102 550 1104
rect 552 1108 560 1110
rect 552 1104 554 1108
rect 558 1104 560 1108
rect 552 1102 560 1104
rect 564 1108 572 1110
rect 564 1104 566 1108
rect 570 1104 572 1108
rect 580 1106 582 1110
rect 586 1106 588 1110
rect 580 1104 588 1106
rect 590 1110 598 1112
rect 590 1106 592 1110
rect 596 1106 598 1110
rect 590 1104 598 1106
rect 564 1102 572 1104
rect 508 1097 510 1101
rect 514 1097 516 1101
rect 580 1100 588 1102
rect 542 1098 550 1100
rect 508 1095 516 1097
rect 528 1096 536 1098
rect 28 1090 36 1092
rect 64 1090 72 1092
rect 84 1091 92 1093
rect 40 1088 48 1090
rect 12 1086 20 1088
rect 28 1086 36 1088
rect 2 1082 10 1084
rect 2 1078 4 1082
rect 8 1078 10 1082
rect 2 1076 10 1078
rect 12 1082 20 1084
rect 12 1078 14 1082
rect 18 1078 20 1082
rect 28 1082 30 1086
rect 34 1082 36 1086
rect 40 1084 42 1088
rect 46 1084 48 1088
rect 40 1082 48 1084
rect 50 1088 58 1090
rect 50 1084 52 1088
rect 56 1084 58 1088
rect 50 1082 58 1084
rect 64 1086 72 1088
rect 64 1082 66 1086
rect 70 1082 72 1086
rect 84 1087 86 1091
rect 90 1087 92 1091
rect 84 1085 92 1087
rect 94 1091 102 1093
rect 94 1087 96 1091
rect 100 1087 102 1091
rect 296 1092 304 1094
rect 296 1088 298 1092
rect 302 1088 304 1092
rect 94 1085 102 1087
rect 112 1085 120 1087
rect 28 1080 36 1082
rect 64 1080 72 1082
rect 84 1081 92 1083
rect 40 1078 48 1080
rect 12 1076 20 1078
rect 28 1076 36 1078
rect 2 1072 10 1074
rect 2 1068 4 1072
rect 8 1068 10 1072
rect 2 1066 10 1068
rect 12 1072 20 1074
rect 12 1068 14 1072
rect 18 1068 20 1072
rect 28 1072 30 1076
rect 34 1072 36 1076
rect 40 1074 42 1078
rect 46 1074 48 1078
rect 40 1072 48 1074
rect 50 1078 58 1080
rect 50 1074 52 1078
rect 56 1074 58 1078
rect 50 1072 58 1074
rect 64 1076 72 1078
rect 64 1072 66 1076
rect 70 1072 72 1076
rect 84 1077 86 1081
rect 90 1077 92 1081
rect 84 1075 92 1077
rect 94 1081 102 1083
rect 94 1077 96 1081
rect 100 1077 102 1081
rect 112 1081 114 1085
rect 118 1081 120 1085
rect 112 1079 120 1081
rect 122 1085 130 1087
rect 122 1081 124 1085
rect 128 1081 130 1085
rect 122 1079 130 1081
rect 132 1085 140 1087
rect 132 1081 134 1085
rect 138 1081 140 1085
rect 132 1079 140 1081
rect 142 1085 150 1087
rect 142 1081 144 1085
rect 148 1081 150 1085
rect 142 1079 150 1081
rect 152 1085 160 1087
rect 152 1081 154 1085
rect 158 1081 160 1085
rect 152 1079 160 1081
rect 162 1085 170 1087
rect 162 1081 164 1085
rect 168 1081 170 1085
rect 162 1079 170 1081
rect 172 1085 180 1087
rect 172 1081 174 1085
rect 178 1081 180 1085
rect 172 1079 180 1081
rect 182 1085 190 1087
rect 182 1081 184 1085
rect 188 1081 190 1085
rect 182 1079 190 1081
rect 192 1085 200 1087
rect 192 1081 194 1085
rect 198 1081 200 1085
rect 192 1079 200 1081
rect 202 1085 210 1087
rect 202 1081 204 1085
rect 208 1081 210 1085
rect 202 1079 210 1081
rect 212 1085 220 1087
rect 212 1081 214 1085
rect 218 1081 220 1085
rect 212 1079 220 1081
rect 222 1085 230 1087
rect 222 1081 224 1085
rect 228 1081 230 1085
rect 222 1079 230 1081
rect 232 1085 240 1087
rect 296 1086 304 1088
rect 498 1091 506 1093
rect 498 1087 500 1091
rect 504 1087 506 1091
rect 232 1081 234 1085
rect 238 1081 240 1085
rect 360 1085 368 1087
rect 232 1079 240 1081
rect 296 1082 304 1084
rect 296 1078 298 1082
rect 302 1078 304 1082
rect 360 1081 362 1085
rect 366 1081 368 1085
rect 360 1079 368 1081
rect 370 1085 378 1087
rect 370 1081 372 1085
rect 376 1081 378 1085
rect 370 1079 378 1081
rect 380 1085 388 1087
rect 380 1081 382 1085
rect 386 1081 388 1085
rect 380 1079 388 1081
rect 390 1085 398 1087
rect 390 1081 392 1085
rect 396 1081 398 1085
rect 390 1079 398 1081
rect 400 1085 408 1087
rect 400 1081 402 1085
rect 406 1081 408 1085
rect 400 1079 408 1081
rect 410 1085 418 1087
rect 410 1081 412 1085
rect 416 1081 418 1085
rect 410 1079 418 1081
rect 420 1085 428 1087
rect 420 1081 422 1085
rect 426 1081 428 1085
rect 420 1079 428 1081
rect 430 1085 438 1087
rect 430 1081 432 1085
rect 436 1081 438 1085
rect 430 1079 438 1081
rect 440 1085 448 1087
rect 440 1081 442 1085
rect 446 1081 448 1085
rect 440 1079 448 1081
rect 450 1085 458 1087
rect 450 1081 452 1085
rect 456 1081 458 1085
rect 450 1079 458 1081
rect 460 1085 468 1087
rect 460 1081 462 1085
rect 466 1081 468 1085
rect 460 1079 468 1081
rect 470 1085 478 1087
rect 470 1081 472 1085
rect 476 1081 478 1085
rect 470 1079 478 1081
rect 480 1085 488 1087
rect 498 1085 506 1087
rect 508 1091 516 1093
rect 508 1087 510 1091
rect 514 1087 516 1091
rect 528 1092 530 1096
rect 534 1092 536 1096
rect 542 1094 544 1098
rect 548 1094 550 1098
rect 542 1092 550 1094
rect 552 1098 560 1100
rect 552 1094 554 1098
rect 558 1094 560 1098
rect 552 1092 560 1094
rect 564 1098 572 1100
rect 564 1094 566 1098
rect 570 1094 572 1098
rect 580 1096 582 1100
rect 586 1096 588 1100
rect 580 1094 588 1096
rect 590 1100 598 1102
rect 590 1096 592 1100
rect 596 1096 598 1100
rect 590 1094 598 1096
rect 564 1092 572 1094
rect 528 1090 536 1092
rect 580 1090 588 1092
rect 542 1088 550 1090
rect 508 1085 516 1087
rect 528 1086 536 1088
rect 480 1081 482 1085
rect 486 1081 488 1085
rect 480 1079 488 1081
rect 498 1081 506 1083
rect 94 1075 102 1077
rect 112 1075 120 1077
rect 28 1070 36 1072
rect 64 1070 72 1072
rect 84 1071 92 1073
rect 40 1068 48 1070
rect 12 1066 20 1068
rect 28 1066 36 1068
rect 2 1062 10 1064
rect 2 1058 4 1062
rect 8 1058 10 1062
rect 2 1056 10 1058
rect 12 1062 20 1064
rect 12 1058 14 1062
rect 18 1058 20 1062
rect 28 1062 30 1066
rect 34 1062 36 1066
rect 40 1064 42 1068
rect 46 1064 48 1068
rect 40 1062 48 1064
rect 50 1068 58 1070
rect 50 1064 52 1068
rect 56 1064 58 1068
rect 50 1062 58 1064
rect 64 1066 72 1068
rect 64 1062 66 1066
rect 70 1062 72 1066
rect 84 1067 86 1071
rect 90 1067 92 1071
rect 84 1065 92 1067
rect 94 1071 102 1073
rect 94 1067 96 1071
rect 100 1067 102 1071
rect 112 1071 114 1075
rect 118 1071 120 1075
rect 112 1069 120 1071
rect 122 1075 130 1077
rect 122 1071 124 1075
rect 128 1071 130 1075
rect 122 1069 130 1071
rect 132 1075 140 1077
rect 132 1071 134 1075
rect 138 1071 140 1075
rect 132 1069 140 1071
rect 142 1075 150 1077
rect 142 1071 144 1075
rect 148 1071 150 1075
rect 142 1069 150 1071
rect 152 1075 160 1077
rect 152 1071 154 1075
rect 158 1071 160 1075
rect 152 1069 160 1071
rect 162 1075 170 1077
rect 162 1071 164 1075
rect 168 1071 170 1075
rect 162 1069 170 1071
rect 172 1075 180 1077
rect 172 1071 174 1075
rect 178 1071 180 1075
rect 172 1069 180 1071
rect 182 1075 190 1077
rect 182 1071 184 1075
rect 188 1071 190 1075
rect 182 1069 190 1071
rect 192 1075 200 1077
rect 192 1071 194 1075
rect 198 1071 200 1075
rect 192 1069 200 1071
rect 202 1075 210 1077
rect 202 1071 204 1075
rect 208 1071 210 1075
rect 202 1069 210 1071
rect 212 1075 220 1077
rect 212 1071 214 1075
rect 218 1071 220 1075
rect 212 1069 220 1071
rect 222 1075 230 1077
rect 222 1071 224 1075
rect 228 1071 230 1075
rect 222 1069 230 1071
rect 232 1075 240 1077
rect 296 1076 304 1078
rect 498 1077 500 1081
rect 504 1077 506 1081
rect 232 1071 234 1075
rect 238 1071 240 1075
rect 360 1075 368 1077
rect 232 1069 240 1071
rect 296 1072 304 1074
rect 94 1065 102 1067
rect 296 1068 298 1072
rect 302 1068 304 1072
rect 360 1071 362 1075
rect 366 1071 368 1075
rect 360 1069 368 1071
rect 370 1075 378 1077
rect 370 1071 372 1075
rect 376 1071 378 1075
rect 370 1069 378 1071
rect 380 1075 388 1077
rect 380 1071 382 1075
rect 386 1071 388 1075
rect 380 1069 388 1071
rect 390 1075 398 1077
rect 390 1071 392 1075
rect 396 1071 398 1075
rect 390 1069 398 1071
rect 400 1075 408 1077
rect 400 1071 402 1075
rect 406 1071 408 1075
rect 400 1069 408 1071
rect 410 1075 418 1077
rect 410 1071 412 1075
rect 416 1071 418 1075
rect 410 1069 418 1071
rect 420 1075 428 1077
rect 420 1071 422 1075
rect 426 1071 428 1075
rect 420 1069 428 1071
rect 430 1075 438 1077
rect 430 1071 432 1075
rect 436 1071 438 1075
rect 430 1069 438 1071
rect 440 1075 448 1077
rect 440 1071 442 1075
rect 446 1071 448 1075
rect 440 1069 448 1071
rect 450 1075 458 1077
rect 450 1071 452 1075
rect 456 1071 458 1075
rect 450 1069 458 1071
rect 460 1075 468 1077
rect 460 1071 462 1075
rect 466 1071 468 1075
rect 460 1069 468 1071
rect 470 1075 478 1077
rect 470 1071 472 1075
rect 476 1071 478 1075
rect 470 1069 478 1071
rect 480 1075 488 1077
rect 498 1075 506 1077
rect 508 1081 516 1083
rect 508 1077 510 1081
rect 514 1077 516 1081
rect 528 1082 530 1086
rect 534 1082 536 1086
rect 542 1084 544 1088
rect 548 1084 550 1088
rect 542 1082 550 1084
rect 552 1088 560 1090
rect 552 1084 554 1088
rect 558 1084 560 1088
rect 552 1082 560 1084
rect 564 1088 572 1090
rect 564 1084 566 1088
rect 570 1084 572 1088
rect 580 1086 582 1090
rect 586 1086 588 1090
rect 580 1084 588 1086
rect 590 1090 598 1092
rect 590 1086 592 1090
rect 596 1086 598 1090
rect 590 1084 598 1086
rect 564 1082 572 1084
rect 528 1080 536 1082
rect 580 1080 588 1082
rect 542 1078 550 1080
rect 508 1075 516 1077
rect 528 1076 536 1078
rect 480 1071 482 1075
rect 486 1071 488 1075
rect 480 1069 488 1071
rect 498 1071 506 1073
rect 296 1066 304 1068
rect 498 1067 500 1071
rect 504 1067 506 1071
rect 498 1065 506 1067
rect 508 1071 516 1073
rect 508 1067 510 1071
rect 514 1067 516 1071
rect 528 1072 530 1076
rect 534 1072 536 1076
rect 542 1074 544 1078
rect 548 1074 550 1078
rect 542 1072 550 1074
rect 552 1078 560 1080
rect 552 1074 554 1078
rect 558 1074 560 1078
rect 552 1072 560 1074
rect 564 1078 572 1080
rect 564 1074 566 1078
rect 570 1074 572 1078
rect 580 1076 582 1080
rect 586 1076 588 1080
rect 580 1074 588 1076
rect 590 1080 598 1082
rect 590 1076 592 1080
rect 596 1076 598 1080
rect 590 1074 598 1076
rect 564 1072 572 1074
rect 528 1070 536 1072
rect 580 1070 588 1072
rect 542 1068 550 1070
rect 508 1065 516 1067
rect 528 1066 536 1068
rect 28 1060 36 1062
rect 64 1060 72 1062
rect 84 1061 92 1063
rect 40 1058 48 1060
rect 12 1056 20 1058
rect 28 1056 36 1058
rect 2 1052 10 1054
rect 2 1048 4 1052
rect 8 1048 10 1052
rect 2 1046 10 1048
rect 12 1052 20 1054
rect 12 1048 14 1052
rect 18 1048 20 1052
rect 28 1052 30 1056
rect 34 1052 36 1056
rect 40 1054 42 1058
rect 46 1054 48 1058
rect 40 1052 48 1054
rect 50 1058 58 1060
rect 50 1054 52 1058
rect 56 1054 58 1058
rect 84 1057 86 1061
rect 90 1057 92 1061
rect 84 1055 92 1057
rect 94 1061 102 1063
rect 94 1057 96 1061
rect 100 1057 102 1061
rect 94 1055 102 1057
rect 296 1062 304 1064
rect 296 1058 298 1062
rect 302 1058 304 1062
rect 296 1056 304 1058
rect 498 1061 506 1063
rect 498 1057 500 1061
rect 504 1057 506 1061
rect 498 1055 506 1057
rect 508 1061 516 1063
rect 508 1057 510 1061
rect 514 1057 516 1061
rect 528 1062 530 1066
rect 534 1062 536 1066
rect 542 1064 544 1068
rect 548 1064 550 1068
rect 542 1062 550 1064
rect 552 1068 560 1070
rect 552 1064 554 1068
rect 558 1064 560 1068
rect 552 1062 560 1064
rect 564 1068 572 1070
rect 564 1064 566 1068
rect 570 1064 572 1068
rect 580 1066 582 1070
rect 586 1066 588 1070
rect 580 1064 588 1066
rect 590 1070 598 1072
rect 590 1066 592 1070
rect 596 1066 598 1070
rect 590 1064 598 1066
rect 564 1062 572 1064
rect 528 1060 536 1062
rect 580 1060 588 1062
rect 508 1055 516 1057
rect 542 1058 550 1060
rect 542 1054 544 1058
rect 548 1054 550 1058
rect 50 1052 58 1054
rect 296 1052 304 1054
rect 542 1052 550 1054
rect 552 1058 560 1060
rect 552 1054 554 1058
rect 558 1054 560 1058
rect 552 1052 560 1054
rect 564 1058 572 1060
rect 564 1054 566 1058
rect 570 1054 572 1058
rect 580 1056 582 1060
rect 586 1056 588 1060
rect 580 1054 588 1056
rect 590 1060 598 1062
rect 590 1056 592 1060
rect 596 1056 598 1060
rect 590 1054 598 1056
rect 564 1052 572 1054
rect 28 1050 36 1052
rect 84 1050 92 1052
rect 40 1048 48 1050
rect 12 1046 20 1048
rect 28 1046 36 1048
rect 2 1042 10 1044
rect 2 1038 4 1042
rect 8 1038 10 1042
rect 2 1036 10 1038
rect 12 1042 20 1044
rect 12 1038 14 1042
rect 18 1038 20 1042
rect 28 1042 30 1046
rect 34 1042 36 1046
rect 40 1044 42 1048
rect 46 1044 48 1048
rect 40 1042 48 1044
rect 50 1048 58 1050
rect 50 1044 52 1048
rect 56 1044 58 1048
rect 50 1042 58 1044
rect 64 1047 72 1049
rect 64 1043 66 1047
rect 70 1043 72 1047
rect 84 1046 86 1050
rect 90 1046 92 1050
rect 84 1044 92 1046
rect 94 1050 102 1052
rect 94 1046 96 1050
rect 100 1046 102 1050
rect 94 1044 102 1046
rect 104 1050 112 1052
rect 104 1046 106 1050
rect 110 1046 112 1050
rect 104 1044 112 1046
rect 114 1050 122 1052
rect 114 1046 116 1050
rect 120 1046 122 1050
rect 114 1044 122 1046
rect 124 1050 132 1052
rect 124 1046 126 1050
rect 130 1046 132 1050
rect 124 1044 132 1046
rect 134 1050 142 1052
rect 134 1046 136 1050
rect 140 1046 142 1050
rect 134 1044 142 1046
rect 144 1050 152 1052
rect 144 1046 146 1050
rect 150 1046 152 1050
rect 144 1044 152 1046
rect 154 1050 162 1052
rect 154 1046 156 1050
rect 160 1046 162 1050
rect 154 1044 162 1046
rect 164 1050 172 1052
rect 164 1046 166 1050
rect 170 1046 172 1050
rect 164 1044 172 1046
rect 174 1050 182 1052
rect 174 1046 176 1050
rect 180 1046 182 1050
rect 174 1044 182 1046
rect 184 1050 192 1052
rect 184 1046 186 1050
rect 190 1046 192 1050
rect 184 1044 192 1046
rect 194 1050 202 1052
rect 194 1046 196 1050
rect 200 1046 202 1050
rect 194 1044 202 1046
rect 204 1050 212 1052
rect 204 1046 206 1050
rect 210 1046 212 1050
rect 204 1044 212 1046
rect 214 1050 222 1052
rect 214 1046 216 1050
rect 220 1046 222 1050
rect 214 1044 222 1046
rect 224 1050 232 1052
rect 224 1046 226 1050
rect 230 1046 232 1050
rect 296 1048 298 1052
rect 302 1048 304 1052
rect 296 1046 304 1048
rect 368 1050 376 1052
rect 368 1046 370 1050
rect 374 1046 376 1050
rect 224 1044 232 1046
rect 368 1044 376 1046
rect 378 1050 386 1052
rect 378 1046 380 1050
rect 384 1046 386 1050
rect 378 1044 386 1046
rect 388 1050 396 1052
rect 388 1046 390 1050
rect 394 1046 396 1050
rect 388 1044 396 1046
rect 398 1050 406 1052
rect 398 1046 400 1050
rect 404 1046 406 1050
rect 398 1044 406 1046
rect 408 1050 416 1052
rect 408 1046 410 1050
rect 414 1046 416 1050
rect 408 1044 416 1046
rect 418 1050 426 1052
rect 418 1046 420 1050
rect 424 1046 426 1050
rect 418 1044 426 1046
rect 428 1050 436 1052
rect 428 1046 430 1050
rect 434 1046 436 1050
rect 428 1044 436 1046
rect 438 1050 446 1052
rect 438 1046 440 1050
rect 444 1046 446 1050
rect 438 1044 446 1046
rect 448 1050 456 1052
rect 448 1046 450 1050
rect 454 1046 456 1050
rect 448 1044 456 1046
rect 458 1050 466 1052
rect 458 1046 460 1050
rect 464 1046 466 1050
rect 458 1044 466 1046
rect 468 1050 476 1052
rect 468 1046 470 1050
rect 474 1046 476 1050
rect 468 1044 476 1046
rect 478 1050 486 1052
rect 478 1046 480 1050
rect 484 1046 486 1050
rect 478 1044 486 1046
rect 488 1050 496 1052
rect 488 1046 490 1050
rect 494 1046 496 1050
rect 488 1044 496 1046
rect 498 1050 506 1052
rect 498 1046 500 1050
rect 504 1046 506 1050
rect 498 1044 506 1046
rect 508 1050 516 1052
rect 580 1050 588 1052
rect 508 1046 510 1050
rect 514 1046 516 1050
rect 508 1044 516 1046
rect 528 1047 536 1049
rect 28 1040 36 1042
rect 64 1041 72 1043
rect 296 1042 304 1044
rect 40 1038 48 1040
rect 12 1036 20 1038
rect 28 1036 36 1038
rect 2 1032 10 1034
rect 2 1028 4 1032
rect 8 1028 10 1032
rect 2 1026 10 1028
rect 12 1032 20 1034
rect 12 1028 14 1032
rect 18 1028 20 1032
rect 28 1032 30 1036
rect 34 1032 36 1036
rect 40 1034 42 1038
rect 46 1034 48 1038
rect 40 1032 48 1034
rect 50 1038 58 1040
rect 50 1034 52 1038
rect 56 1034 58 1038
rect 50 1032 58 1034
rect 64 1037 72 1039
rect 64 1033 66 1037
rect 70 1033 72 1037
rect 296 1038 298 1042
rect 302 1038 304 1042
rect 528 1043 530 1047
rect 534 1043 536 1047
rect 528 1041 536 1043
rect 542 1048 550 1050
rect 542 1044 544 1048
rect 548 1044 550 1048
rect 542 1042 550 1044
rect 552 1048 560 1050
rect 552 1044 554 1048
rect 558 1044 560 1048
rect 552 1042 560 1044
rect 564 1048 572 1050
rect 564 1044 566 1048
rect 570 1044 572 1048
rect 580 1046 582 1050
rect 586 1046 588 1050
rect 580 1044 588 1046
rect 590 1050 598 1052
rect 590 1046 592 1050
rect 596 1046 598 1050
rect 590 1044 598 1046
rect 564 1042 572 1044
rect 580 1040 588 1042
rect 296 1036 304 1038
rect 528 1037 536 1039
rect 28 1030 36 1032
rect 64 1031 72 1033
rect 296 1032 304 1034
rect 40 1028 48 1030
rect 12 1026 20 1028
rect 28 1026 36 1028
rect 2 1022 10 1024
rect 2 1018 4 1022
rect 8 1018 10 1022
rect 2 1016 10 1018
rect 12 1022 20 1024
rect 12 1018 14 1022
rect 18 1018 20 1022
rect 28 1022 30 1026
rect 34 1022 36 1026
rect 40 1024 42 1028
rect 46 1024 48 1028
rect 40 1022 48 1024
rect 50 1028 58 1030
rect 50 1024 52 1028
rect 56 1024 58 1028
rect 50 1022 58 1024
rect 64 1027 72 1029
rect 64 1023 66 1027
rect 70 1023 72 1027
rect 296 1028 298 1032
rect 302 1028 304 1032
rect 528 1033 530 1037
rect 534 1033 536 1037
rect 528 1031 536 1033
rect 542 1038 550 1040
rect 542 1034 544 1038
rect 548 1034 550 1038
rect 542 1032 550 1034
rect 552 1038 560 1040
rect 552 1034 554 1038
rect 558 1034 560 1038
rect 552 1032 560 1034
rect 564 1038 572 1040
rect 564 1034 566 1038
rect 570 1034 572 1038
rect 580 1036 582 1040
rect 586 1036 588 1040
rect 580 1034 588 1036
rect 590 1040 598 1042
rect 590 1036 592 1040
rect 596 1036 598 1040
rect 590 1034 598 1036
rect 564 1032 572 1034
rect 580 1030 588 1032
rect 296 1026 304 1028
rect 528 1027 536 1029
rect 28 1020 36 1022
rect 64 1021 72 1023
rect 82 1022 90 1024
rect 40 1018 48 1020
rect 12 1016 20 1018
rect 28 1016 36 1018
rect 2 1012 10 1014
rect 2 1008 4 1012
rect 8 1008 10 1012
rect 2 1006 10 1008
rect 12 1012 20 1014
rect 12 1008 14 1012
rect 18 1008 20 1012
rect 28 1012 30 1016
rect 34 1012 36 1016
rect 40 1014 42 1018
rect 46 1014 48 1018
rect 40 1012 48 1014
rect 50 1018 58 1020
rect 50 1014 52 1018
rect 56 1014 58 1018
rect 50 1012 58 1014
rect 64 1017 72 1019
rect 64 1013 66 1017
rect 70 1013 72 1017
rect 82 1018 84 1022
rect 88 1018 90 1022
rect 82 1016 90 1018
rect 92 1022 100 1024
rect 92 1018 94 1022
rect 98 1018 100 1022
rect 92 1016 100 1018
rect 102 1022 110 1024
rect 102 1018 104 1022
rect 108 1018 110 1022
rect 102 1016 110 1018
rect 112 1022 120 1024
rect 112 1018 114 1022
rect 118 1018 120 1022
rect 112 1016 120 1018
rect 122 1022 130 1024
rect 122 1018 124 1022
rect 128 1018 130 1022
rect 122 1016 130 1018
rect 132 1022 140 1024
rect 132 1018 134 1022
rect 138 1018 140 1022
rect 132 1016 140 1018
rect 142 1022 150 1024
rect 142 1018 144 1022
rect 148 1018 150 1022
rect 142 1016 150 1018
rect 152 1022 160 1024
rect 152 1018 154 1022
rect 158 1018 160 1022
rect 152 1016 160 1018
rect 162 1022 170 1024
rect 162 1018 164 1022
rect 168 1018 170 1022
rect 162 1016 170 1018
rect 172 1022 180 1024
rect 172 1018 174 1022
rect 178 1018 180 1022
rect 172 1016 180 1018
rect 182 1022 190 1024
rect 182 1018 184 1022
rect 188 1018 190 1022
rect 182 1016 190 1018
rect 192 1022 200 1024
rect 192 1018 194 1022
rect 198 1018 200 1022
rect 192 1016 200 1018
rect 202 1022 210 1024
rect 202 1018 204 1022
rect 208 1018 210 1022
rect 202 1016 210 1018
rect 212 1022 220 1024
rect 212 1018 214 1022
rect 218 1018 220 1022
rect 212 1016 220 1018
rect 222 1022 230 1024
rect 222 1018 224 1022
rect 228 1018 230 1022
rect 222 1016 230 1018
rect 296 1022 304 1024
rect 296 1018 298 1022
rect 302 1018 304 1022
rect 296 1016 304 1018
rect 367 1022 375 1024
rect 367 1018 369 1022
rect 373 1018 375 1022
rect 367 1016 375 1018
rect 377 1022 385 1024
rect 377 1018 379 1022
rect 383 1018 385 1022
rect 377 1016 385 1018
rect 387 1022 395 1024
rect 387 1018 389 1022
rect 393 1018 395 1022
rect 387 1016 395 1018
rect 397 1022 405 1024
rect 397 1018 399 1022
rect 403 1018 405 1022
rect 397 1016 405 1018
rect 407 1022 415 1024
rect 407 1018 409 1022
rect 413 1018 415 1022
rect 407 1016 415 1018
rect 417 1022 425 1024
rect 417 1018 419 1022
rect 423 1018 425 1022
rect 417 1016 425 1018
rect 427 1022 435 1024
rect 427 1018 429 1022
rect 433 1018 435 1022
rect 427 1016 435 1018
rect 437 1022 445 1024
rect 437 1018 439 1022
rect 443 1018 445 1022
rect 437 1016 445 1018
rect 447 1022 455 1024
rect 447 1018 449 1022
rect 453 1018 455 1022
rect 447 1016 455 1018
rect 457 1022 465 1024
rect 457 1018 459 1022
rect 463 1018 465 1022
rect 457 1016 465 1018
rect 467 1022 475 1024
rect 467 1018 469 1022
rect 473 1018 475 1022
rect 467 1016 475 1018
rect 477 1022 485 1024
rect 477 1018 479 1022
rect 483 1018 485 1022
rect 477 1016 485 1018
rect 487 1022 495 1024
rect 487 1018 489 1022
rect 493 1018 495 1022
rect 487 1016 495 1018
rect 497 1022 505 1024
rect 497 1018 499 1022
rect 503 1018 505 1022
rect 497 1016 505 1018
rect 507 1022 515 1024
rect 507 1018 509 1022
rect 513 1018 515 1022
rect 528 1023 530 1027
rect 534 1023 536 1027
rect 528 1021 536 1023
rect 542 1028 550 1030
rect 542 1024 544 1028
rect 548 1024 550 1028
rect 542 1022 550 1024
rect 552 1028 560 1030
rect 552 1024 554 1028
rect 558 1024 560 1028
rect 552 1022 560 1024
rect 564 1028 572 1030
rect 564 1024 566 1028
rect 570 1024 572 1028
rect 580 1026 582 1030
rect 586 1026 588 1030
rect 580 1024 588 1026
rect 590 1030 598 1032
rect 590 1026 592 1030
rect 596 1026 598 1030
rect 590 1024 598 1026
rect 564 1022 572 1024
rect 580 1020 588 1022
rect 507 1016 515 1018
rect 528 1017 536 1019
rect 28 1010 36 1012
rect 64 1011 72 1013
rect 296 1012 304 1014
rect 528 1013 530 1017
rect 534 1013 536 1017
rect 82 1010 90 1012
rect 40 1008 48 1010
rect 12 1006 20 1008
rect 28 1006 36 1008
rect 2 1002 10 1004
rect 2 998 4 1002
rect 8 998 10 1002
rect 2 996 10 998
rect 12 1002 20 1004
rect 12 998 14 1002
rect 18 998 20 1002
rect 28 1002 30 1006
rect 34 1002 36 1006
rect 40 1004 42 1008
rect 46 1004 48 1008
rect 40 1002 48 1004
rect 50 1008 58 1010
rect 50 1004 52 1008
rect 56 1004 58 1008
rect 50 1002 58 1004
rect 64 1007 72 1009
rect 64 1003 66 1007
rect 70 1003 72 1007
rect 82 1006 84 1010
rect 88 1006 90 1010
rect 82 1004 90 1006
rect 92 1010 100 1012
rect 92 1006 94 1010
rect 98 1006 100 1010
rect 92 1004 100 1006
rect 102 1010 110 1012
rect 102 1006 104 1010
rect 108 1006 110 1010
rect 102 1004 110 1006
rect 112 1010 120 1012
rect 112 1006 114 1010
rect 118 1006 120 1010
rect 112 1004 120 1006
rect 122 1010 130 1012
rect 122 1006 124 1010
rect 128 1006 130 1010
rect 122 1004 130 1006
rect 132 1010 140 1012
rect 132 1006 134 1010
rect 138 1006 140 1010
rect 132 1004 140 1006
rect 142 1010 150 1012
rect 142 1006 144 1010
rect 148 1006 150 1010
rect 142 1004 150 1006
rect 152 1010 160 1012
rect 152 1006 154 1010
rect 158 1006 160 1010
rect 152 1004 160 1006
rect 162 1010 170 1012
rect 162 1006 164 1010
rect 168 1006 170 1010
rect 162 1004 170 1006
rect 172 1010 180 1012
rect 172 1006 174 1010
rect 178 1006 180 1010
rect 172 1004 180 1006
rect 182 1010 190 1012
rect 182 1006 184 1010
rect 188 1006 190 1010
rect 182 1004 190 1006
rect 192 1010 200 1012
rect 192 1006 194 1010
rect 198 1006 200 1010
rect 192 1004 200 1006
rect 202 1010 210 1012
rect 202 1006 204 1010
rect 208 1006 210 1010
rect 202 1004 210 1006
rect 212 1010 220 1012
rect 212 1006 214 1010
rect 218 1006 220 1010
rect 212 1004 220 1006
rect 222 1010 230 1012
rect 222 1006 224 1010
rect 228 1006 230 1010
rect 296 1008 298 1012
rect 302 1008 304 1012
rect 296 1006 304 1008
rect 367 1010 375 1012
rect 367 1006 369 1010
rect 373 1006 375 1010
rect 222 1004 230 1006
rect 367 1004 375 1006
rect 377 1010 385 1012
rect 377 1006 379 1010
rect 383 1006 385 1010
rect 377 1004 385 1006
rect 387 1010 395 1012
rect 387 1006 389 1010
rect 393 1006 395 1010
rect 387 1004 395 1006
rect 397 1010 405 1012
rect 397 1006 399 1010
rect 403 1006 405 1010
rect 397 1004 405 1006
rect 407 1010 415 1012
rect 407 1006 409 1010
rect 413 1006 415 1010
rect 407 1004 415 1006
rect 417 1010 425 1012
rect 417 1006 419 1010
rect 423 1006 425 1010
rect 417 1004 425 1006
rect 427 1010 435 1012
rect 427 1006 429 1010
rect 433 1006 435 1010
rect 427 1004 435 1006
rect 437 1010 445 1012
rect 437 1006 439 1010
rect 443 1006 445 1010
rect 437 1004 445 1006
rect 447 1010 455 1012
rect 447 1006 449 1010
rect 453 1006 455 1010
rect 447 1004 455 1006
rect 457 1010 465 1012
rect 457 1006 459 1010
rect 463 1006 465 1010
rect 457 1004 465 1006
rect 467 1010 475 1012
rect 467 1006 469 1010
rect 473 1006 475 1010
rect 467 1004 475 1006
rect 477 1010 485 1012
rect 477 1006 479 1010
rect 483 1006 485 1010
rect 477 1004 485 1006
rect 487 1010 495 1012
rect 487 1006 489 1010
rect 493 1006 495 1010
rect 487 1004 495 1006
rect 497 1010 505 1012
rect 497 1006 499 1010
rect 503 1006 505 1010
rect 497 1004 505 1006
rect 507 1010 515 1012
rect 528 1011 536 1013
rect 542 1018 550 1020
rect 542 1014 544 1018
rect 548 1014 550 1018
rect 542 1012 550 1014
rect 552 1018 560 1020
rect 552 1014 554 1018
rect 558 1014 560 1018
rect 552 1012 560 1014
rect 564 1018 572 1020
rect 564 1014 566 1018
rect 570 1014 572 1018
rect 580 1016 582 1020
rect 586 1016 588 1020
rect 580 1014 588 1016
rect 590 1020 598 1022
rect 590 1016 592 1020
rect 596 1016 598 1020
rect 590 1014 598 1016
rect 564 1012 572 1014
rect 580 1010 588 1012
rect 507 1006 509 1010
rect 513 1006 515 1010
rect 507 1004 515 1006
rect 528 1007 536 1009
rect 28 1000 36 1002
rect 64 1001 72 1003
rect 296 1002 304 1004
rect 40 998 48 1000
rect 12 996 20 998
rect 28 996 36 998
rect 2 992 10 994
rect 2 988 4 992
rect 8 988 10 992
rect 2 986 10 988
rect 12 992 20 994
rect 12 988 14 992
rect 18 988 20 992
rect 28 992 30 996
rect 34 992 36 996
rect 40 994 42 998
rect 46 994 48 998
rect 40 992 48 994
rect 50 998 58 1000
rect 50 994 52 998
rect 56 994 58 998
rect 50 992 58 994
rect 64 997 72 999
rect 64 993 66 997
rect 70 993 72 997
rect 296 998 298 1002
rect 302 998 304 1002
rect 528 1003 530 1007
rect 534 1003 536 1007
rect 528 1001 536 1003
rect 542 1008 550 1010
rect 542 1004 544 1008
rect 548 1004 550 1008
rect 542 1002 550 1004
rect 552 1008 560 1010
rect 552 1004 554 1008
rect 558 1004 560 1008
rect 552 1002 560 1004
rect 564 1008 572 1010
rect 564 1004 566 1008
rect 570 1004 572 1008
rect 580 1006 582 1010
rect 586 1006 588 1010
rect 580 1004 588 1006
rect 590 1010 598 1012
rect 590 1006 592 1010
rect 596 1006 598 1010
rect 590 1004 598 1006
rect 564 1002 572 1004
rect 580 1000 588 1002
rect 296 996 304 998
rect 528 997 536 999
rect 28 990 36 992
rect 64 991 72 993
rect 296 992 304 994
rect 40 988 48 990
rect 12 986 20 988
rect 28 986 36 988
rect 2 982 10 984
rect 2 978 4 982
rect 8 978 10 982
rect 2 976 10 978
rect 12 982 20 984
rect 12 978 14 982
rect 18 978 20 982
rect 28 982 30 986
rect 34 982 36 986
rect 40 984 42 988
rect 46 984 48 988
rect 40 982 48 984
rect 50 988 58 990
rect 50 984 52 988
rect 56 984 58 988
rect 50 982 58 984
rect 64 987 72 989
rect 64 983 66 987
rect 70 983 72 987
rect 296 988 298 992
rect 302 988 304 992
rect 528 993 530 997
rect 534 993 536 997
rect 528 991 536 993
rect 542 998 550 1000
rect 542 994 544 998
rect 548 994 550 998
rect 542 992 550 994
rect 552 998 560 1000
rect 552 994 554 998
rect 558 994 560 998
rect 552 992 560 994
rect 564 998 572 1000
rect 564 994 566 998
rect 570 994 572 998
rect 580 996 582 1000
rect 586 996 588 1000
rect 580 994 588 996
rect 590 1000 598 1002
rect 590 996 592 1000
rect 596 996 598 1000
rect 590 994 598 996
rect 564 992 572 994
rect 580 990 588 992
rect 296 986 304 988
rect 528 987 536 989
rect 28 980 36 982
rect 64 981 72 983
rect 84 984 92 986
rect 84 980 86 984
rect 90 980 92 984
rect 40 978 48 980
rect 12 976 20 978
rect 28 976 36 978
rect 2 972 10 974
rect 2 968 4 972
rect 8 968 10 972
rect 2 966 10 968
rect 12 972 20 974
rect 12 968 14 972
rect 18 968 20 972
rect 28 972 30 976
rect 34 972 36 976
rect 40 974 42 978
rect 46 974 48 978
rect 40 972 48 974
rect 50 978 58 980
rect 84 978 92 980
rect 94 984 102 986
rect 94 980 96 984
rect 100 980 102 984
rect 94 978 102 980
rect 104 984 112 986
rect 104 980 106 984
rect 110 980 112 984
rect 104 978 112 980
rect 114 984 122 986
rect 114 980 116 984
rect 120 980 122 984
rect 114 978 122 980
rect 124 984 132 986
rect 124 980 126 984
rect 130 980 132 984
rect 124 978 132 980
rect 134 984 142 986
rect 134 980 136 984
rect 140 980 142 984
rect 134 978 142 980
rect 144 984 152 986
rect 144 980 146 984
rect 150 980 152 984
rect 144 978 152 980
rect 154 984 162 986
rect 154 980 156 984
rect 160 980 162 984
rect 154 978 162 980
rect 164 984 172 986
rect 164 980 166 984
rect 170 980 172 984
rect 164 978 172 980
rect 174 984 182 986
rect 174 980 176 984
rect 180 980 182 984
rect 174 978 182 980
rect 184 984 192 986
rect 184 980 186 984
rect 190 980 192 984
rect 184 978 192 980
rect 194 984 202 986
rect 194 980 196 984
rect 200 980 202 984
rect 194 978 202 980
rect 204 984 212 986
rect 204 980 206 984
rect 210 980 212 984
rect 204 978 212 980
rect 214 984 222 986
rect 214 980 216 984
rect 220 980 222 984
rect 214 978 222 980
rect 224 984 232 986
rect 368 984 376 986
rect 224 980 226 984
rect 230 980 232 984
rect 224 978 232 980
rect 296 982 304 984
rect 296 978 298 982
rect 302 978 304 982
rect 368 980 370 984
rect 374 980 376 984
rect 368 978 376 980
rect 378 984 386 986
rect 378 980 380 984
rect 384 980 386 984
rect 378 978 386 980
rect 388 984 396 986
rect 388 980 390 984
rect 394 980 396 984
rect 388 978 396 980
rect 398 984 406 986
rect 398 980 400 984
rect 404 980 406 984
rect 398 978 406 980
rect 408 984 416 986
rect 408 980 410 984
rect 414 980 416 984
rect 408 978 416 980
rect 418 984 426 986
rect 418 980 420 984
rect 424 980 426 984
rect 418 978 426 980
rect 428 984 436 986
rect 428 980 430 984
rect 434 980 436 984
rect 428 978 436 980
rect 438 984 446 986
rect 438 980 440 984
rect 444 980 446 984
rect 438 978 446 980
rect 448 984 456 986
rect 448 980 450 984
rect 454 980 456 984
rect 448 978 456 980
rect 458 984 466 986
rect 458 980 460 984
rect 464 980 466 984
rect 458 978 466 980
rect 468 984 476 986
rect 468 980 470 984
rect 474 980 476 984
rect 468 978 476 980
rect 478 984 486 986
rect 478 980 480 984
rect 484 980 486 984
rect 478 978 486 980
rect 488 984 496 986
rect 488 980 490 984
rect 494 980 496 984
rect 488 978 496 980
rect 498 984 506 986
rect 498 980 500 984
rect 504 980 506 984
rect 498 978 506 980
rect 508 984 516 986
rect 508 980 510 984
rect 514 980 516 984
rect 528 983 530 987
rect 534 983 536 987
rect 528 981 536 983
rect 542 988 550 990
rect 542 984 544 988
rect 548 984 550 988
rect 542 982 550 984
rect 552 988 560 990
rect 552 984 554 988
rect 558 984 560 988
rect 552 982 560 984
rect 564 988 572 990
rect 564 984 566 988
rect 570 984 572 988
rect 580 986 582 990
rect 586 986 588 990
rect 580 984 588 986
rect 590 990 598 992
rect 590 986 592 990
rect 596 986 598 990
rect 590 984 598 986
rect 564 982 572 984
rect 580 980 588 982
rect 508 978 516 980
rect 542 978 550 980
rect 50 974 52 978
rect 56 974 58 978
rect 296 976 304 978
rect 50 972 58 974
rect 84 973 92 975
rect 28 970 36 972
rect 40 968 48 970
rect 12 966 20 968
rect 28 966 36 968
rect 2 962 10 964
rect 2 958 4 962
rect 8 958 10 962
rect 2 956 10 958
rect 12 962 20 964
rect 12 958 14 962
rect 18 958 20 962
rect 28 962 30 966
rect 34 962 36 966
rect 40 964 42 968
rect 46 964 48 968
rect 40 962 48 964
rect 50 968 58 970
rect 50 964 52 968
rect 56 964 58 968
rect 84 969 86 973
rect 90 969 92 973
rect 84 967 92 969
rect 94 973 102 975
rect 542 974 544 978
rect 548 974 550 978
rect 94 969 96 973
rect 100 969 102 973
rect 94 967 102 969
rect 296 972 304 974
rect 296 968 298 972
rect 302 968 304 972
rect 296 966 304 968
rect 500 972 508 974
rect 500 968 502 972
rect 506 968 508 972
rect 500 966 508 968
rect 510 972 518 974
rect 542 972 550 974
rect 552 978 560 980
rect 552 974 554 978
rect 558 974 560 978
rect 552 972 560 974
rect 564 978 572 980
rect 564 974 566 978
rect 570 974 572 978
rect 580 976 582 980
rect 586 976 588 980
rect 580 974 588 976
rect 590 980 598 982
rect 590 976 592 980
rect 596 976 598 980
rect 590 974 598 976
rect 564 972 572 974
rect 510 968 512 972
rect 516 968 518 972
rect 580 970 588 972
rect 542 968 550 970
rect 510 966 518 968
rect 528 966 536 968
rect 50 962 58 964
rect 84 963 92 965
rect 28 960 36 962
rect 64 960 72 962
rect 40 958 48 960
rect 12 956 20 958
rect 28 956 36 958
rect 2 952 10 954
rect 2 948 4 952
rect 8 948 10 952
rect 2 946 10 948
rect 12 952 20 954
rect 12 948 14 952
rect 18 948 20 952
rect 28 952 30 956
rect 34 952 36 956
rect 40 954 42 958
rect 46 954 48 958
rect 40 952 48 954
rect 50 958 58 960
rect 50 954 52 958
rect 56 954 58 958
rect 64 956 66 960
rect 70 956 72 960
rect 84 959 86 963
rect 90 959 92 963
rect 84 957 92 959
rect 94 963 102 965
rect 94 959 96 963
rect 100 959 102 963
rect 94 957 102 959
rect 296 962 304 964
rect 296 958 298 962
rect 302 958 304 962
rect 500 962 508 964
rect 500 958 502 962
rect 506 958 508 962
rect 64 954 72 956
rect 112 956 120 958
rect 50 952 58 954
rect 84 953 92 955
rect 28 950 36 952
rect 64 950 72 952
rect 40 948 48 950
rect 12 946 20 948
rect 28 946 36 948
rect 2 942 10 944
rect 2 938 4 942
rect 8 938 10 942
rect 2 936 10 938
rect 12 942 20 944
rect 12 938 14 942
rect 18 938 20 942
rect 28 942 30 946
rect 34 942 36 946
rect 40 944 42 948
rect 46 944 48 948
rect 40 942 48 944
rect 50 948 58 950
rect 50 944 52 948
rect 56 944 58 948
rect 64 946 66 950
rect 70 946 72 950
rect 84 949 86 953
rect 90 949 92 953
rect 84 947 92 949
rect 94 953 102 955
rect 94 949 96 953
rect 100 949 102 953
rect 112 952 114 956
rect 118 952 120 956
rect 112 950 120 952
rect 122 956 130 958
rect 122 952 124 956
rect 128 952 130 956
rect 122 950 130 952
rect 132 956 140 958
rect 132 952 134 956
rect 138 952 140 956
rect 132 950 140 952
rect 142 956 150 958
rect 142 952 144 956
rect 148 952 150 956
rect 142 950 150 952
rect 152 956 160 958
rect 152 952 154 956
rect 158 952 160 956
rect 152 950 160 952
rect 162 956 170 958
rect 162 952 164 956
rect 168 952 170 956
rect 162 950 170 952
rect 172 956 180 958
rect 172 952 174 956
rect 178 952 180 956
rect 172 950 180 952
rect 182 956 190 958
rect 182 952 184 956
rect 188 952 190 956
rect 182 950 190 952
rect 192 956 200 958
rect 192 952 194 956
rect 198 952 200 956
rect 192 950 200 952
rect 202 956 210 958
rect 202 952 204 956
rect 208 952 210 956
rect 202 950 210 952
rect 212 956 220 958
rect 212 952 214 956
rect 218 952 220 956
rect 212 950 220 952
rect 222 956 230 958
rect 222 952 224 956
rect 228 952 230 956
rect 222 950 230 952
rect 232 956 240 958
rect 296 956 304 958
rect 360 956 368 958
rect 232 952 234 956
rect 238 952 240 956
rect 232 950 240 952
rect 296 952 304 954
rect 94 947 102 949
rect 296 948 298 952
rect 302 948 304 952
rect 360 952 362 956
rect 366 952 368 956
rect 360 950 368 952
rect 370 956 378 958
rect 370 952 372 956
rect 376 952 378 956
rect 370 950 378 952
rect 380 956 388 958
rect 380 952 382 956
rect 386 952 388 956
rect 380 950 388 952
rect 390 956 398 958
rect 390 952 392 956
rect 396 952 398 956
rect 390 950 398 952
rect 400 956 408 958
rect 400 952 402 956
rect 406 952 408 956
rect 400 950 408 952
rect 410 956 418 958
rect 410 952 412 956
rect 416 952 418 956
rect 410 950 418 952
rect 420 956 428 958
rect 420 952 422 956
rect 426 952 428 956
rect 420 950 428 952
rect 430 956 438 958
rect 430 952 432 956
rect 436 952 438 956
rect 430 950 438 952
rect 440 956 448 958
rect 440 952 442 956
rect 446 952 448 956
rect 440 950 448 952
rect 450 956 458 958
rect 450 952 452 956
rect 456 952 458 956
rect 450 950 458 952
rect 460 956 468 958
rect 460 952 462 956
rect 466 952 468 956
rect 460 950 468 952
rect 470 956 478 958
rect 470 952 472 956
rect 476 952 478 956
rect 470 950 478 952
rect 480 956 488 958
rect 500 956 508 958
rect 510 962 518 964
rect 510 958 512 962
rect 516 958 518 962
rect 528 962 530 966
rect 534 962 536 966
rect 542 964 544 968
rect 548 964 550 968
rect 542 962 550 964
rect 552 968 560 970
rect 552 964 554 968
rect 558 964 560 968
rect 552 962 560 964
rect 564 968 572 970
rect 564 964 566 968
rect 570 964 572 968
rect 580 966 582 970
rect 586 966 588 970
rect 580 964 588 966
rect 590 970 598 972
rect 590 966 592 970
rect 596 966 598 970
rect 590 964 598 966
rect 564 962 572 964
rect 528 960 536 962
rect 580 960 588 962
rect 542 958 550 960
rect 510 956 518 958
rect 528 956 536 958
rect 480 952 482 956
rect 486 952 488 956
rect 480 950 488 952
rect 500 952 508 954
rect 500 948 502 952
rect 506 948 508 952
rect 64 944 72 946
rect 112 946 120 948
rect 50 942 58 944
rect 84 943 92 945
rect 28 940 36 942
rect 64 940 72 942
rect 40 938 48 940
rect 12 936 20 938
rect 28 936 36 938
rect 2 932 10 934
rect 2 928 4 932
rect 8 928 10 932
rect 2 926 10 928
rect 12 932 20 934
rect 12 928 14 932
rect 18 928 20 932
rect 28 932 30 936
rect 34 932 36 936
rect 40 934 42 938
rect 46 934 48 938
rect 40 932 48 934
rect 50 938 58 940
rect 50 934 52 938
rect 56 934 58 938
rect 64 936 66 940
rect 70 936 72 940
rect 84 939 86 943
rect 90 939 92 943
rect 84 937 92 939
rect 94 943 102 945
rect 94 939 96 943
rect 100 939 102 943
rect 112 942 114 946
rect 118 942 120 946
rect 112 940 120 942
rect 122 946 130 948
rect 122 942 124 946
rect 128 942 130 946
rect 122 940 130 942
rect 132 946 140 948
rect 132 942 134 946
rect 138 942 140 946
rect 132 940 140 942
rect 142 946 150 948
rect 142 942 144 946
rect 148 942 150 946
rect 142 940 150 942
rect 152 946 160 948
rect 152 942 154 946
rect 158 942 160 946
rect 152 940 160 942
rect 162 946 170 948
rect 162 942 164 946
rect 168 942 170 946
rect 162 940 170 942
rect 172 946 180 948
rect 172 942 174 946
rect 178 942 180 946
rect 172 940 180 942
rect 182 946 190 948
rect 182 942 184 946
rect 188 942 190 946
rect 182 940 190 942
rect 192 946 200 948
rect 192 942 194 946
rect 198 942 200 946
rect 192 940 200 942
rect 202 946 210 948
rect 202 942 204 946
rect 208 942 210 946
rect 202 940 210 942
rect 212 946 220 948
rect 212 942 214 946
rect 218 942 220 946
rect 212 940 220 942
rect 222 946 230 948
rect 222 942 224 946
rect 228 942 230 946
rect 222 940 230 942
rect 232 946 240 948
rect 296 946 304 948
rect 360 946 368 948
rect 232 942 234 946
rect 238 942 240 946
rect 232 940 240 942
rect 296 942 304 944
rect 94 937 102 939
rect 296 938 298 942
rect 302 938 304 942
rect 360 942 362 946
rect 366 942 368 946
rect 360 940 368 942
rect 370 946 378 948
rect 370 942 372 946
rect 376 942 378 946
rect 370 940 378 942
rect 380 946 388 948
rect 380 942 382 946
rect 386 942 388 946
rect 380 940 388 942
rect 390 946 398 948
rect 390 942 392 946
rect 396 942 398 946
rect 390 940 398 942
rect 400 946 408 948
rect 400 942 402 946
rect 406 942 408 946
rect 400 940 408 942
rect 410 946 418 948
rect 410 942 412 946
rect 416 942 418 946
rect 410 940 418 942
rect 420 946 428 948
rect 420 942 422 946
rect 426 942 428 946
rect 420 940 428 942
rect 430 946 438 948
rect 430 942 432 946
rect 436 942 438 946
rect 430 940 438 942
rect 440 946 448 948
rect 440 942 442 946
rect 446 942 448 946
rect 440 940 448 942
rect 450 946 458 948
rect 450 942 452 946
rect 456 942 458 946
rect 450 940 458 942
rect 460 946 468 948
rect 460 942 462 946
rect 466 942 468 946
rect 460 940 468 942
rect 470 946 478 948
rect 470 942 472 946
rect 476 942 478 946
rect 470 940 478 942
rect 480 946 488 948
rect 500 946 508 948
rect 510 952 518 954
rect 510 948 512 952
rect 516 948 518 952
rect 528 952 530 956
rect 534 952 536 956
rect 542 954 544 958
rect 548 954 550 958
rect 542 952 550 954
rect 552 958 560 960
rect 552 954 554 958
rect 558 954 560 958
rect 552 952 560 954
rect 564 958 572 960
rect 564 954 566 958
rect 570 954 572 958
rect 580 956 582 960
rect 586 956 588 960
rect 580 954 588 956
rect 590 960 598 962
rect 590 956 592 960
rect 596 956 598 960
rect 590 954 598 956
rect 564 952 572 954
rect 528 950 536 952
rect 580 950 588 952
rect 542 948 550 950
rect 510 946 518 948
rect 528 946 536 948
rect 480 942 482 946
rect 486 942 488 946
rect 480 940 488 942
rect 500 942 508 944
rect 296 936 304 938
rect 500 938 502 942
rect 506 938 508 942
rect 500 936 508 938
rect 510 942 518 944
rect 510 938 512 942
rect 516 938 518 942
rect 528 942 530 946
rect 534 942 536 946
rect 542 944 544 948
rect 548 944 550 948
rect 542 942 550 944
rect 552 948 560 950
rect 552 944 554 948
rect 558 944 560 948
rect 552 942 560 944
rect 564 948 572 950
rect 564 944 566 948
rect 570 944 572 948
rect 580 946 582 950
rect 586 946 588 950
rect 580 944 588 946
rect 590 950 598 952
rect 590 946 592 950
rect 596 946 598 950
rect 590 944 598 946
rect 564 942 572 944
rect 528 940 536 942
rect 580 940 588 942
rect 542 938 550 940
rect 510 936 518 938
rect 528 936 536 938
rect 64 934 72 936
rect 50 932 58 934
rect 84 933 92 935
rect 28 930 36 932
rect 64 930 72 932
rect 40 928 48 930
rect 12 926 20 928
rect 28 926 36 928
rect 2 922 10 924
rect 2 918 4 922
rect 8 918 10 922
rect 2 916 10 918
rect 12 922 20 924
rect 12 918 14 922
rect 18 918 20 922
rect 28 922 30 926
rect 34 922 36 926
rect 40 924 42 928
rect 46 924 48 928
rect 40 922 48 924
rect 50 928 58 930
rect 50 924 52 928
rect 56 924 58 928
rect 64 926 66 930
rect 70 926 72 930
rect 84 929 86 933
rect 90 929 92 933
rect 84 927 92 929
rect 94 933 102 935
rect 94 929 96 933
rect 100 929 102 933
rect 94 927 102 929
rect 296 932 304 934
rect 296 928 298 932
rect 302 928 304 932
rect 296 926 304 928
rect 500 932 508 934
rect 500 928 502 932
rect 506 928 508 932
rect 500 926 508 928
rect 510 932 518 934
rect 510 928 512 932
rect 516 928 518 932
rect 528 932 530 936
rect 534 932 536 936
rect 542 934 544 938
rect 548 934 550 938
rect 542 932 550 934
rect 552 938 560 940
rect 552 934 554 938
rect 558 934 560 938
rect 552 932 560 934
rect 564 938 572 940
rect 564 934 566 938
rect 570 934 572 938
rect 580 936 582 940
rect 586 936 588 940
rect 580 934 588 936
rect 590 940 598 942
rect 590 936 592 940
rect 596 936 598 940
rect 590 934 598 936
rect 564 932 572 934
rect 528 930 536 932
rect 580 930 588 932
rect 542 928 550 930
rect 510 926 518 928
rect 528 926 536 928
rect 64 924 72 926
rect 50 922 58 924
rect 296 922 304 924
rect 528 922 530 926
rect 534 922 536 926
rect 542 924 544 928
rect 548 924 550 928
rect 542 922 550 924
rect 552 928 560 930
rect 552 924 554 928
rect 558 924 560 928
rect 552 922 560 924
rect 564 928 572 930
rect 564 924 566 928
rect 570 924 572 928
rect 580 926 582 930
rect 586 926 588 930
rect 580 924 588 926
rect 590 930 598 932
rect 590 926 592 930
rect 596 926 598 930
rect 590 924 598 926
rect 564 922 572 924
rect 28 920 36 922
rect 64 920 72 922
rect 40 918 48 920
rect 12 916 20 918
rect 28 916 36 918
rect 2 912 10 914
rect 2 908 4 912
rect 8 908 10 912
rect 2 906 10 908
rect 12 912 20 914
rect 12 908 14 912
rect 18 908 20 912
rect 28 912 30 916
rect 34 912 36 916
rect 40 914 42 918
rect 46 914 48 918
rect 40 912 48 914
rect 50 918 58 920
rect 50 914 52 918
rect 56 914 58 918
rect 64 916 66 920
rect 70 916 72 920
rect 64 914 72 916
rect 82 920 90 922
rect 82 916 84 920
rect 88 916 90 920
rect 82 914 90 916
rect 92 920 100 922
rect 92 916 94 920
rect 98 916 100 920
rect 92 914 100 916
rect 102 920 110 922
rect 102 916 104 920
rect 108 916 110 920
rect 102 914 110 916
rect 112 920 120 922
rect 112 916 114 920
rect 118 916 120 920
rect 112 914 120 916
rect 122 920 130 922
rect 122 916 124 920
rect 128 916 130 920
rect 122 914 130 916
rect 132 920 140 922
rect 132 916 134 920
rect 138 916 140 920
rect 132 914 140 916
rect 142 920 150 922
rect 142 916 144 920
rect 148 916 150 920
rect 142 914 150 916
rect 152 920 160 922
rect 152 916 154 920
rect 158 916 160 920
rect 152 914 160 916
rect 162 920 170 922
rect 162 916 164 920
rect 168 916 170 920
rect 162 914 170 916
rect 172 920 180 922
rect 172 916 174 920
rect 178 916 180 920
rect 172 914 180 916
rect 182 920 190 922
rect 182 916 184 920
rect 188 916 190 920
rect 182 914 190 916
rect 192 920 200 922
rect 192 916 194 920
rect 198 916 200 920
rect 192 914 200 916
rect 202 920 210 922
rect 202 916 204 920
rect 208 916 210 920
rect 202 914 210 916
rect 212 920 220 922
rect 212 916 214 920
rect 218 916 220 920
rect 212 914 220 916
rect 222 920 230 922
rect 222 916 224 920
rect 228 916 230 920
rect 296 918 298 922
rect 302 918 304 922
rect 296 916 304 918
rect 370 920 378 922
rect 370 916 372 920
rect 376 916 378 920
rect 222 914 230 916
rect 370 914 378 916
rect 380 920 388 922
rect 380 916 382 920
rect 386 916 388 920
rect 380 914 388 916
rect 390 920 398 922
rect 390 916 392 920
rect 396 916 398 920
rect 390 914 398 916
rect 400 920 408 922
rect 400 916 402 920
rect 406 916 408 920
rect 400 914 408 916
rect 410 920 418 922
rect 410 916 412 920
rect 416 916 418 920
rect 410 914 418 916
rect 420 920 428 922
rect 420 916 422 920
rect 426 916 428 920
rect 420 914 428 916
rect 430 920 438 922
rect 430 916 432 920
rect 436 916 438 920
rect 430 914 438 916
rect 440 920 448 922
rect 440 916 442 920
rect 446 916 448 920
rect 440 914 448 916
rect 450 920 458 922
rect 450 916 452 920
rect 456 916 458 920
rect 450 914 458 916
rect 460 920 468 922
rect 460 916 462 920
rect 466 916 468 920
rect 460 914 468 916
rect 470 920 478 922
rect 470 916 472 920
rect 476 916 478 920
rect 470 914 478 916
rect 480 920 488 922
rect 480 916 482 920
rect 486 916 488 920
rect 480 914 488 916
rect 490 920 498 922
rect 490 916 492 920
rect 496 916 498 920
rect 490 914 498 916
rect 500 920 508 922
rect 500 916 502 920
rect 506 916 508 920
rect 500 914 508 916
rect 510 920 518 922
rect 528 920 536 922
rect 580 920 588 922
rect 510 916 512 920
rect 516 916 518 920
rect 542 918 550 920
rect 510 914 518 916
rect 528 916 536 918
rect 50 912 58 914
rect 296 912 304 914
rect 28 910 36 912
rect 64 910 72 912
rect 40 908 48 910
rect 12 906 20 908
rect 28 906 36 908
rect 2 902 10 904
rect 2 898 4 902
rect 8 898 10 902
rect 2 896 10 898
rect 12 902 20 904
rect 12 898 14 902
rect 18 898 20 902
rect 28 902 30 906
rect 34 902 36 906
rect 40 904 42 908
rect 46 904 48 908
rect 40 902 48 904
rect 50 908 58 910
rect 50 904 52 908
rect 56 904 58 908
rect 64 906 66 910
rect 70 906 72 910
rect 296 908 298 912
rect 302 908 304 912
rect 528 912 530 916
rect 534 912 536 916
rect 542 914 544 918
rect 548 914 550 918
rect 542 912 550 914
rect 552 918 560 920
rect 552 914 554 918
rect 558 914 560 918
rect 552 912 560 914
rect 564 918 572 920
rect 564 914 566 918
rect 570 914 572 918
rect 580 916 582 920
rect 586 916 588 920
rect 580 914 588 916
rect 590 920 598 922
rect 590 916 592 920
rect 596 916 598 920
rect 590 914 598 916
rect 564 912 572 914
rect 528 910 536 912
rect 580 910 588 912
rect 296 906 304 908
rect 542 908 550 910
rect 64 904 72 906
rect 542 904 544 908
rect 548 904 550 908
rect 50 902 58 904
rect 296 902 304 904
rect 542 902 550 904
rect 552 908 560 910
rect 552 904 554 908
rect 558 904 560 908
rect 552 902 560 904
rect 564 908 572 910
rect 564 904 566 908
rect 570 904 572 908
rect 580 906 582 910
rect 586 906 588 910
rect 580 904 588 906
rect 590 910 598 912
rect 590 906 592 910
rect 596 906 598 910
rect 590 904 598 906
rect 564 902 572 904
rect 28 900 36 902
rect 40 898 48 900
rect 12 896 20 898
rect 28 896 36 898
rect 2 892 10 894
rect 2 888 4 892
rect 8 888 10 892
rect 2 886 10 888
rect 12 892 20 894
rect 12 888 14 892
rect 18 888 20 892
rect 28 892 30 896
rect 34 892 36 896
rect 40 894 42 898
rect 46 894 48 898
rect 40 892 48 894
rect 50 898 58 900
rect 50 894 52 898
rect 56 894 58 898
rect 296 898 298 902
rect 302 898 304 902
rect 580 900 588 902
rect 296 896 304 898
rect 542 898 550 900
rect 542 894 544 898
rect 548 894 550 898
rect 50 892 58 894
rect 80 892 88 894
rect 28 890 36 892
rect 40 888 48 890
rect 12 886 20 888
rect 28 886 36 888
rect 2 882 10 884
rect 2 878 4 882
rect 8 878 10 882
rect 2 876 10 878
rect 12 882 20 884
rect 12 878 14 882
rect 18 878 20 882
rect 28 882 30 886
rect 34 882 36 886
rect 40 884 42 888
rect 46 884 48 888
rect 40 882 48 884
rect 50 888 58 890
rect 50 884 52 888
rect 56 884 58 888
rect 80 888 82 892
rect 86 888 88 892
rect 80 886 88 888
rect 91 892 99 894
rect 91 888 93 892
rect 97 888 99 892
rect 91 886 99 888
rect 102 892 110 894
rect 102 888 104 892
rect 108 888 110 892
rect 102 886 110 888
rect 113 892 121 894
rect 113 888 115 892
rect 119 888 121 892
rect 113 886 121 888
rect 123 892 131 894
rect 123 888 125 892
rect 129 888 131 892
rect 123 886 131 888
rect 133 892 141 894
rect 133 888 135 892
rect 139 888 141 892
rect 133 886 141 888
rect 143 892 151 894
rect 143 888 145 892
rect 149 888 151 892
rect 143 886 151 888
rect 153 892 161 894
rect 153 888 155 892
rect 159 888 161 892
rect 153 886 161 888
rect 163 892 171 894
rect 163 888 165 892
rect 169 888 171 892
rect 163 886 171 888
rect 173 892 181 894
rect 173 888 175 892
rect 179 888 181 892
rect 173 886 181 888
rect 183 892 191 894
rect 183 888 185 892
rect 189 888 191 892
rect 183 886 191 888
rect 193 892 201 894
rect 193 888 195 892
rect 199 888 201 892
rect 193 886 201 888
rect 203 892 211 894
rect 203 888 205 892
rect 209 888 211 892
rect 203 886 211 888
rect 213 892 221 894
rect 213 888 215 892
rect 219 888 221 892
rect 213 886 221 888
rect 223 892 231 894
rect 223 888 225 892
rect 229 888 231 892
rect 223 886 231 888
rect 296 892 304 894
rect 296 888 298 892
rect 302 888 304 892
rect 296 886 304 888
rect 369 892 377 894
rect 369 888 371 892
rect 375 888 377 892
rect 369 886 377 888
rect 379 892 387 894
rect 379 888 381 892
rect 385 888 387 892
rect 379 886 387 888
rect 389 892 397 894
rect 389 888 391 892
rect 395 888 397 892
rect 389 886 397 888
rect 399 892 407 894
rect 399 888 401 892
rect 405 888 407 892
rect 399 886 407 888
rect 409 892 417 894
rect 409 888 411 892
rect 415 888 417 892
rect 409 886 417 888
rect 419 892 427 894
rect 419 888 421 892
rect 425 888 427 892
rect 419 886 427 888
rect 429 892 437 894
rect 429 888 431 892
rect 435 888 437 892
rect 429 886 437 888
rect 439 892 447 894
rect 439 888 441 892
rect 445 888 447 892
rect 439 886 447 888
rect 449 892 457 894
rect 449 888 451 892
rect 455 888 457 892
rect 449 886 457 888
rect 459 892 467 894
rect 459 888 461 892
rect 465 888 467 892
rect 459 886 467 888
rect 469 892 477 894
rect 469 888 471 892
rect 475 888 477 892
rect 469 886 477 888
rect 479 892 487 894
rect 479 888 481 892
rect 485 888 487 892
rect 479 886 487 888
rect 490 892 498 894
rect 490 888 492 892
rect 496 888 498 892
rect 490 886 498 888
rect 501 892 509 894
rect 501 888 503 892
rect 507 888 509 892
rect 501 886 509 888
rect 512 892 520 894
rect 542 892 550 894
rect 552 898 560 900
rect 552 894 554 898
rect 558 894 560 898
rect 552 892 560 894
rect 564 898 572 900
rect 564 894 566 898
rect 570 894 572 898
rect 580 896 582 900
rect 586 896 588 900
rect 580 894 588 896
rect 590 900 598 902
rect 590 896 592 900
rect 596 896 598 900
rect 590 894 598 896
rect 564 892 572 894
rect 512 888 514 892
rect 518 888 520 892
rect 580 890 588 892
rect 512 886 520 888
rect 542 888 550 890
rect 542 884 544 888
rect 548 884 550 888
rect 50 882 58 884
rect 296 882 304 884
rect 542 882 550 884
rect 552 888 560 890
rect 552 884 554 888
rect 558 884 560 888
rect 552 882 560 884
rect 564 888 572 890
rect 564 884 566 888
rect 570 884 572 888
rect 580 886 582 890
rect 586 886 588 890
rect 580 884 588 886
rect 590 890 598 892
rect 590 886 592 890
rect 596 886 598 890
rect 590 884 598 886
rect 564 882 572 884
rect 28 880 36 882
rect 93 880 101 882
rect 12 876 20 878
rect 40 878 48 880
rect 40 874 42 878
rect 46 874 48 878
rect 2 872 10 874
rect 2 868 4 872
rect 8 868 10 872
rect 2 866 10 868
rect 12 872 20 874
rect 40 872 48 874
rect 50 878 58 880
rect 50 874 52 878
rect 56 874 58 878
rect 93 876 95 880
rect 99 876 101 880
rect 93 874 101 876
rect 103 880 111 882
rect 103 876 105 880
rect 109 876 111 880
rect 103 874 111 876
rect 113 880 121 882
rect 113 876 115 880
rect 119 876 121 880
rect 113 874 121 876
rect 123 880 131 882
rect 123 876 125 880
rect 129 876 131 880
rect 123 874 131 876
rect 133 880 141 882
rect 133 876 135 880
rect 139 876 141 880
rect 133 874 141 876
rect 143 880 151 882
rect 143 876 145 880
rect 149 876 151 880
rect 143 874 151 876
rect 153 880 161 882
rect 153 876 155 880
rect 159 876 161 880
rect 153 874 161 876
rect 163 880 171 882
rect 163 876 165 880
rect 169 876 171 880
rect 163 874 171 876
rect 173 880 181 882
rect 173 876 175 880
rect 179 876 181 880
rect 173 874 181 876
rect 183 880 191 882
rect 183 876 185 880
rect 189 876 191 880
rect 183 874 191 876
rect 193 880 201 882
rect 193 876 195 880
rect 199 876 201 880
rect 193 874 201 876
rect 203 880 211 882
rect 203 876 205 880
rect 209 876 211 880
rect 203 874 211 876
rect 213 880 221 882
rect 213 876 215 880
rect 219 876 221 880
rect 213 874 221 876
rect 223 880 231 882
rect 223 876 225 880
rect 229 876 231 880
rect 296 878 298 882
rect 302 878 304 882
rect 296 876 304 878
rect 369 880 377 882
rect 369 876 371 880
rect 375 876 377 880
rect 223 874 231 876
rect 369 874 377 876
rect 379 880 387 882
rect 379 876 381 880
rect 385 876 387 880
rect 379 874 387 876
rect 389 880 397 882
rect 389 876 391 880
rect 395 876 397 880
rect 389 874 397 876
rect 399 880 407 882
rect 399 876 401 880
rect 405 876 407 880
rect 399 874 407 876
rect 409 880 417 882
rect 409 876 411 880
rect 415 876 417 880
rect 409 874 417 876
rect 419 880 427 882
rect 419 876 421 880
rect 425 876 427 880
rect 419 874 427 876
rect 429 880 437 882
rect 429 876 431 880
rect 435 876 437 880
rect 429 874 437 876
rect 439 880 447 882
rect 439 876 441 880
rect 445 876 447 880
rect 439 874 447 876
rect 449 880 457 882
rect 449 876 451 880
rect 455 876 457 880
rect 449 874 457 876
rect 459 880 467 882
rect 459 876 461 880
rect 465 876 467 880
rect 459 874 467 876
rect 469 880 477 882
rect 469 876 471 880
rect 475 876 477 880
rect 469 874 477 876
rect 479 880 487 882
rect 479 876 481 880
rect 485 876 487 880
rect 479 874 487 876
rect 489 880 497 882
rect 489 876 491 880
rect 495 876 497 880
rect 489 874 497 876
rect 499 880 507 882
rect 580 880 588 882
rect 499 876 501 880
rect 505 876 507 880
rect 499 874 507 876
rect 542 878 550 880
rect 542 874 544 878
rect 548 874 550 878
rect 50 872 58 874
rect 296 872 304 874
rect 542 872 550 874
rect 552 878 560 880
rect 552 874 554 878
rect 558 874 560 878
rect 580 876 582 880
rect 586 876 588 880
rect 580 874 588 876
rect 590 880 598 882
rect 590 876 592 880
rect 596 876 598 880
rect 590 874 598 876
rect 552 872 560 874
rect 12 868 14 872
rect 18 868 20 872
rect 12 866 20 868
rect 40 868 48 870
rect 40 864 42 868
rect 46 864 48 868
rect 2 862 10 864
rect 2 858 4 862
rect 8 858 10 862
rect 2 856 10 858
rect 12 862 20 864
rect 40 862 48 864
rect 50 868 58 870
rect 50 864 52 868
rect 56 864 58 868
rect 50 862 58 864
rect 64 868 72 870
rect 64 864 66 868
rect 70 864 72 868
rect 64 862 72 864
rect 74 868 82 870
rect 74 864 76 868
rect 80 864 82 868
rect 74 862 82 864
rect 93 868 101 870
rect 93 864 95 868
rect 99 864 101 868
rect 93 862 101 864
rect 103 868 111 870
rect 103 864 105 868
rect 109 864 111 868
rect 103 862 111 864
rect 113 868 121 870
rect 113 864 115 868
rect 119 864 121 868
rect 113 862 121 864
rect 123 868 131 870
rect 123 864 125 868
rect 129 864 131 868
rect 123 862 131 864
rect 133 868 141 870
rect 133 864 135 868
rect 139 864 141 868
rect 133 862 141 864
rect 143 868 151 870
rect 143 864 145 868
rect 149 864 151 868
rect 143 862 151 864
rect 153 868 161 870
rect 153 864 155 868
rect 159 864 161 868
rect 153 862 161 864
rect 163 868 171 870
rect 163 864 165 868
rect 169 864 171 868
rect 163 862 171 864
rect 173 868 181 870
rect 173 864 175 868
rect 179 864 181 868
rect 173 862 181 864
rect 183 868 191 870
rect 183 864 185 868
rect 189 864 191 868
rect 183 862 191 864
rect 193 868 201 870
rect 193 864 195 868
rect 199 864 201 868
rect 193 862 201 864
rect 203 868 211 870
rect 203 864 205 868
rect 209 864 211 868
rect 203 862 211 864
rect 213 868 221 870
rect 213 864 215 868
rect 219 864 221 868
rect 213 862 221 864
rect 223 868 231 870
rect 223 864 225 868
rect 229 864 231 868
rect 296 868 298 872
rect 302 868 304 872
rect 580 870 588 872
rect 296 866 304 868
rect 369 868 377 870
rect 223 862 231 864
rect 369 864 371 868
rect 375 864 377 868
rect 369 862 377 864
rect 379 868 387 870
rect 379 864 381 868
rect 385 864 387 868
rect 379 862 387 864
rect 389 868 397 870
rect 389 864 391 868
rect 395 864 397 868
rect 389 862 397 864
rect 399 868 407 870
rect 399 864 401 868
rect 405 864 407 868
rect 399 862 407 864
rect 409 868 417 870
rect 409 864 411 868
rect 415 864 417 868
rect 409 862 417 864
rect 419 868 427 870
rect 419 864 421 868
rect 425 864 427 868
rect 419 862 427 864
rect 429 868 437 870
rect 429 864 431 868
rect 435 864 437 868
rect 429 862 437 864
rect 439 868 447 870
rect 439 864 441 868
rect 445 864 447 868
rect 439 862 447 864
rect 449 868 457 870
rect 449 864 451 868
rect 455 864 457 868
rect 449 862 457 864
rect 459 868 467 870
rect 459 864 461 868
rect 465 864 467 868
rect 459 862 467 864
rect 469 868 477 870
rect 469 864 471 868
rect 475 864 477 868
rect 469 862 477 864
rect 479 868 487 870
rect 479 864 481 868
rect 485 864 487 868
rect 479 862 487 864
rect 489 868 497 870
rect 489 864 491 868
rect 495 864 497 868
rect 489 862 497 864
rect 499 868 507 870
rect 499 864 501 868
rect 505 864 507 868
rect 499 862 507 864
rect 518 868 526 870
rect 518 864 520 868
rect 524 864 526 868
rect 518 862 526 864
rect 528 868 536 870
rect 528 864 530 868
rect 534 864 536 868
rect 528 862 536 864
rect 542 868 550 870
rect 542 864 544 868
rect 548 864 550 868
rect 542 862 550 864
rect 552 868 560 870
rect 552 864 554 868
rect 558 864 560 868
rect 580 866 582 870
rect 586 866 588 870
rect 580 864 588 866
rect 590 870 598 872
rect 590 866 592 870
rect 596 866 598 870
rect 590 864 598 866
rect 552 862 560 864
rect 12 858 14 862
rect 18 858 20 862
rect 12 856 20 858
rect 580 860 588 862
rect 580 856 582 860
rect 586 856 588 860
rect 580 854 588 856
rect 590 860 598 862
rect 590 856 592 860
rect 596 856 598 860
rect 590 854 598 856
rect 2 852 10 854
rect 2 848 4 852
rect 8 848 10 852
rect 2 846 10 848
rect 12 852 20 854
rect 12 848 14 852
rect 18 848 20 852
rect 580 850 588 852
rect 12 846 20 848
rect 30 848 38 850
rect 30 844 32 848
rect 36 844 38 848
rect 2 842 10 844
rect 2 838 4 842
rect 8 838 10 842
rect 2 836 10 838
rect 12 842 20 844
rect 30 842 38 844
rect 40 848 48 850
rect 40 844 42 848
rect 46 844 48 848
rect 40 842 48 844
rect 50 848 58 850
rect 50 844 52 848
rect 56 844 58 848
rect 50 842 58 844
rect 78 848 86 850
rect 78 844 80 848
rect 84 844 86 848
rect 78 842 86 844
rect 88 848 96 850
rect 88 844 90 848
rect 94 844 96 848
rect 88 842 96 844
rect 98 848 106 850
rect 98 844 100 848
rect 104 844 106 848
rect 98 842 106 844
rect 108 848 116 850
rect 108 844 110 848
rect 114 844 116 848
rect 108 842 116 844
rect 118 848 126 850
rect 118 844 120 848
rect 124 844 126 848
rect 118 842 126 844
rect 128 848 136 850
rect 128 844 130 848
rect 134 844 136 848
rect 128 842 136 844
rect 138 848 146 850
rect 138 844 140 848
rect 144 844 146 848
rect 138 842 146 844
rect 148 848 156 850
rect 148 844 150 848
rect 154 844 156 848
rect 148 842 156 844
rect 158 848 166 850
rect 158 844 160 848
rect 164 844 166 848
rect 158 842 166 844
rect 168 848 176 850
rect 168 844 170 848
rect 174 844 176 848
rect 168 842 176 844
rect 178 848 186 850
rect 178 844 180 848
rect 184 844 186 848
rect 178 842 186 844
rect 188 848 196 850
rect 188 844 190 848
rect 194 844 196 848
rect 188 842 196 844
rect 198 848 206 850
rect 198 844 200 848
rect 204 844 206 848
rect 198 842 206 844
rect 208 848 216 850
rect 208 844 210 848
rect 214 844 216 848
rect 208 842 216 844
rect 218 848 226 850
rect 218 844 220 848
rect 224 844 226 848
rect 218 842 226 844
rect 296 848 304 850
rect 296 844 298 848
rect 302 844 304 848
rect 296 842 304 844
rect 368 848 376 850
rect 368 844 370 848
rect 374 844 376 848
rect 368 842 376 844
rect 378 848 386 850
rect 378 844 380 848
rect 384 844 386 848
rect 378 842 386 844
rect 388 848 396 850
rect 388 844 390 848
rect 394 844 396 848
rect 388 842 396 844
rect 398 848 406 850
rect 398 844 400 848
rect 404 844 406 848
rect 398 842 406 844
rect 408 848 416 850
rect 408 844 410 848
rect 414 844 416 848
rect 408 842 416 844
rect 418 848 426 850
rect 418 844 420 848
rect 424 844 426 848
rect 418 842 426 844
rect 428 848 436 850
rect 428 844 430 848
rect 434 844 436 848
rect 428 842 436 844
rect 438 848 446 850
rect 438 844 440 848
rect 444 844 446 848
rect 438 842 446 844
rect 448 848 456 850
rect 448 844 450 848
rect 454 844 456 848
rect 448 842 456 844
rect 458 848 466 850
rect 458 844 460 848
rect 464 844 466 848
rect 458 842 466 844
rect 468 848 476 850
rect 468 844 470 848
rect 474 844 476 848
rect 468 842 476 844
rect 478 848 486 850
rect 478 844 480 848
rect 484 844 486 848
rect 478 842 486 844
rect 488 848 496 850
rect 488 844 490 848
rect 494 844 496 848
rect 488 842 496 844
rect 498 848 506 850
rect 498 844 500 848
rect 504 844 506 848
rect 498 842 506 844
rect 508 848 516 850
rect 508 844 510 848
rect 514 844 516 848
rect 508 842 516 844
rect 518 848 526 850
rect 518 844 520 848
rect 524 844 526 848
rect 518 842 526 844
rect 528 848 536 850
rect 528 844 530 848
rect 534 844 536 848
rect 528 842 536 844
rect 538 848 546 850
rect 538 844 540 848
rect 544 844 546 848
rect 538 842 546 844
rect 548 848 556 850
rect 548 844 550 848
rect 554 844 556 848
rect 548 842 556 844
rect 558 848 566 850
rect 558 844 560 848
rect 564 844 566 848
rect 558 842 566 844
rect 568 848 576 850
rect 568 844 570 848
rect 574 844 576 848
rect 580 846 582 850
rect 586 846 588 850
rect 580 844 588 846
rect 590 850 598 852
rect 590 846 592 850
rect 596 846 598 850
rect 590 844 598 846
rect 568 842 576 844
rect 12 838 14 842
rect 18 838 20 842
rect 580 840 588 842
rect 12 836 20 838
rect 30 837 38 839
rect 2 832 10 834
rect 2 828 4 832
rect 8 828 10 832
rect 2 826 10 828
rect 12 832 20 834
rect 12 828 14 832
rect 18 828 20 832
rect 30 833 32 837
rect 36 833 38 837
rect 30 831 38 833
rect 40 837 48 839
rect 40 833 42 837
rect 46 833 48 837
rect 40 831 48 833
rect 50 837 58 839
rect 50 833 52 837
rect 56 833 58 837
rect 50 831 58 833
rect 78 837 86 839
rect 78 833 80 837
rect 84 833 86 837
rect 78 831 86 833
rect 88 837 96 839
rect 88 833 90 837
rect 94 833 96 837
rect 88 831 96 833
rect 98 837 106 839
rect 98 833 100 837
rect 104 833 106 837
rect 98 831 106 833
rect 108 837 116 839
rect 108 833 110 837
rect 114 833 116 837
rect 108 831 116 833
rect 118 837 126 839
rect 118 833 120 837
rect 124 833 126 837
rect 118 831 126 833
rect 128 837 136 839
rect 128 833 130 837
rect 134 833 136 837
rect 128 831 136 833
rect 138 837 146 839
rect 138 833 140 837
rect 144 833 146 837
rect 138 831 146 833
rect 148 837 156 839
rect 148 833 150 837
rect 154 833 156 837
rect 148 831 156 833
rect 158 837 166 839
rect 158 833 160 837
rect 164 833 166 837
rect 158 831 166 833
rect 168 837 176 839
rect 168 833 170 837
rect 174 833 176 837
rect 168 831 176 833
rect 178 837 186 839
rect 178 833 180 837
rect 184 833 186 837
rect 178 831 186 833
rect 188 837 196 839
rect 188 833 190 837
rect 194 833 196 837
rect 188 831 196 833
rect 198 837 206 839
rect 198 833 200 837
rect 204 833 206 837
rect 198 831 206 833
rect 208 837 216 839
rect 208 833 210 837
rect 214 833 216 837
rect 208 831 216 833
rect 218 837 226 839
rect 218 833 220 837
rect 224 833 226 837
rect 218 831 226 833
rect 296 837 304 839
rect 296 833 298 837
rect 302 833 304 837
rect 296 831 304 833
rect 368 837 376 839
rect 368 833 370 837
rect 374 833 376 837
rect 368 831 376 833
rect 378 837 386 839
rect 378 833 380 837
rect 384 833 386 837
rect 378 831 386 833
rect 388 837 396 839
rect 388 833 390 837
rect 394 833 396 837
rect 388 831 396 833
rect 398 837 406 839
rect 398 833 400 837
rect 404 833 406 837
rect 398 831 406 833
rect 408 837 416 839
rect 408 833 410 837
rect 414 833 416 837
rect 408 831 416 833
rect 418 837 426 839
rect 418 833 420 837
rect 424 833 426 837
rect 418 831 426 833
rect 428 837 436 839
rect 428 833 430 837
rect 434 833 436 837
rect 428 831 436 833
rect 438 837 446 839
rect 438 833 440 837
rect 444 833 446 837
rect 438 831 446 833
rect 448 837 456 839
rect 448 833 450 837
rect 454 833 456 837
rect 448 831 456 833
rect 458 837 466 839
rect 458 833 460 837
rect 464 833 466 837
rect 458 831 466 833
rect 468 837 476 839
rect 468 833 470 837
rect 474 833 476 837
rect 468 831 476 833
rect 478 837 486 839
rect 478 833 480 837
rect 484 833 486 837
rect 478 831 486 833
rect 488 837 496 839
rect 488 833 490 837
rect 494 833 496 837
rect 488 831 496 833
rect 498 837 506 839
rect 498 833 500 837
rect 504 833 506 837
rect 498 831 506 833
rect 508 837 516 839
rect 508 833 510 837
rect 514 833 516 837
rect 508 831 516 833
rect 518 837 526 839
rect 518 833 520 837
rect 524 833 526 837
rect 518 831 526 833
rect 528 837 536 839
rect 528 833 530 837
rect 534 833 536 837
rect 528 831 536 833
rect 538 837 546 839
rect 538 833 540 837
rect 544 833 546 837
rect 538 831 546 833
rect 548 837 556 839
rect 548 833 550 837
rect 554 833 556 837
rect 548 831 556 833
rect 558 837 566 839
rect 558 833 560 837
rect 564 833 566 837
rect 558 831 566 833
rect 568 837 576 839
rect 568 833 570 837
rect 574 833 576 837
rect 580 836 582 840
rect 586 836 588 840
rect 580 834 588 836
rect 590 840 598 842
rect 590 836 592 840
rect 596 836 598 840
rect 590 834 598 836
rect 568 831 576 833
rect 580 830 588 832
rect 12 826 20 828
rect 30 827 38 829
rect 30 823 32 827
rect 36 823 38 827
rect 30 821 38 823
rect 40 827 48 829
rect 40 823 42 827
rect 46 823 48 827
rect 40 821 48 823
rect 50 827 58 829
rect 50 823 52 827
rect 56 823 58 827
rect 50 821 58 823
rect 78 827 86 829
rect 78 823 80 827
rect 84 823 86 827
rect 78 821 86 823
rect 88 827 96 829
rect 88 823 90 827
rect 94 823 96 827
rect 88 821 96 823
rect 98 827 106 829
rect 98 823 100 827
rect 104 823 106 827
rect 98 821 106 823
rect 108 827 116 829
rect 108 823 110 827
rect 114 823 116 827
rect 108 821 116 823
rect 118 827 126 829
rect 118 823 120 827
rect 124 823 126 827
rect 118 821 126 823
rect 128 827 136 829
rect 128 823 130 827
rect 134 823 136 827
rect 128 821 136 823
rect 138 827 146 829
rect 138 823 140 827
rect 144 823 146 827
rect 138 821 146 823
rect 148 827 156 829
rect 148 823 150 827
rect 154 823 156 827
rect 148 821 156 823
rect 158 827 166 829
rect 158 823 160 827
rect 164 823 166 827
rect 158 821 166 823
rect 168 827 176 829
rect 168 823 170 827
rect 174 823 176 827
rect 168 821 176 823
rect 178 827 186 829
rect 178 823 180 827
rect 184 823 186 827
rect 178 821 186 823
rect 188 827 196 829
rect 188 823 190 827
rect 194 823 196 827
rect 188 821 196 823
rect 198 827 206 829
rect 198 823 200 827
rect 204 823 206 827
rect 198 821 206 823
rect 208 827 216 829
rect 208 823 210 827
rect 214 823 216 827
rect 208 821 216 823
rect 218 827 226 829
rect 218 823 220 827
rect 224 823 226 827
rect 218 821 226 823
rect 296 827 304 829
rect 296 823 298 827
rect 302 823 304 827
rect 296 821 304 823
rect 368 827 376 829
rect 368 823 370 827
rect 374 823 376 827
rect 368 821 376 823
rect 378 827 386 829
rect 378 823 380 827
rect 384 823 386 827
rect 378 821 386 823
rect 388 827 396 829
rect 388 823 390 827
rect 394 823 396 827
rect 388 821 396 823
rect 398 827 406 829
rect 398 823 400 827
rect 404 823 406 827
rect 398 821 406 823
rect 408 827 416 829
rect 408 823 410 827
rect 414 823 416 827
rect 408 821 416 823
rect 418 827 426 829
rect 418 823 420 827
rect 424 823 426 827
rect 418 821 426 823
rect 428 827 436 829
rect 428 823 430 827
rect 434 823 436 827
rect 428 821 436 823
rect 438 827 446 829
rect 438 823 440 827
rect 444 823 446 827
rect 438 821 446 823
rect 448 827 456 829
rect 448 823 450 827
rect 454 823 456 827
rect 448 821 456 823
rect 458 827 466 829
rect 458 823 460 827
rect 464 823 466 827
rect 458 821 466 823
rect 468 827 476 829
rect 468 823 470 827
rect 474 823 476 827
rect 468 821 476 823
rect 478 827 486 829
rect 478 823 480 827
rect 484 823 486 827
rect 478 821 486 823
rect 488 827 496 829
rect 488 823 490 827
rect 494 823 496 827
rect 488 821 496 823
rect 498 827 506 829
rect 498 823 500 827
rect 504 823 506 827
rect 498 821 506 823
rect 508 827 516 829
rect 508 823 510 827
rect 514 823 516 827
rect 508 821 516 823
rect 518 827 526 829
rect 518 823 520 827
rect 524 823 526 827
rect 518 821 526 823
rect 528 827 536 829
rect 528 823 530 827
rect 534 823 536 827
rect 528 821 536 823
rect 538 827 546 829
rect 538 823 540 827
rect 544 823 546 827
rect 538 821 546 823
rect 548 827 556 829
rect 548 823 550 827
rect 554 823 556 827
rect 548 821 556 823
rect 558 827 566 829
rect 558 823 560 827
rect 564 823 566 827
rect 558 821 566 823
rect 568 827 576 829
rect 568 823 570 827
rect 574 823 576 827
rect 580 826 582 830
rect 586 826 588 830
rect 580 824 588 826
rect 590 830 598 832
rect 590 826 592 830
rect 596 826 598 830
rect 590 824 598 826
rect 568 821 576 823
rect 590 821 598 823
rect 14 816 22 818
rect 2 812 10 814
rect 2 808 4 812
rect 8 808 10 812
rect 14 812 16 816
rect 20 812 22 816
rect 14 810 22 812
rect 26 816 34 818
rect 26 812 28 816
rect 32 812 34 816
rect 26 810 34 812
rect 36 816 44 818
rect 36 812 38 816
rect 42 812 44 816
rect 36 810 44 812
rect 46 816 54 818
rect 46 812 48 816
rect 52 812 54 816
rect 46 810 54 812
rect 78 816 86 818
rect 78 812 80 816
rect 84 812 86 816
rect 78 810 86 812
rect 88 816 96 818
rect 88 812 90 816
rect 94 812 96 816
rect 88 810 96 812
rect 98 816 106 818
rect 98 812 100 816
rect 104 812 106 816
rect 98 810 106 812
rect 108 816 116 818
rect 108 812 110 816
rect 114 812 116 816
rect 108 810 116 812
rect 118 816 126 818
rect 118 812 120 816
rect 124 812 126 816
rect 118 810 126 812
rect 128 816 136 818
rect 128 812 130 816
rect 134 812 136 816
rect 128 810 136 812
rect 138 816 146 818
rect 138 812 140 816
rect 144 812 146 816
rect 138 810 146 812
rect 148 816 156 818
rect 148 812 150 816
rect 154 812 156 816
rect 148 810 156 812
rect 158 816 166 818
rect 158 812 160 816
rect 164 812 166 816
rect 158 810 166 812
rect 168 816 176 818
rect 168 812 170 816
rect 174 812 176 816
rect 168 810 176 812
rect 178 816 186 818
rect 178 812 180 816
rect 184 812 186 816
rect 178 810 186 812
rect 188 816 196 818
rect 188 812 190 816
rect 194 812 196 816
rect 188 810 196 812
rect 198 816 206 818
rect 198 812 200 816
rect 204 812 206 816
rect 198 810 206 812
rect 208 816 216 818
rect 208 812 210 816
rect 214 812 216 816
rect 590 817 592 821
rect 596 817 598 821
rect 590 815 598 817
rect 208 810 216 812
rect 590 811 598 813
rect 2 806 10 808
rect 14 806 22 808
rect 2 802 10 804
rect 2 798 4 802
rect 8 798 10 802
rect 14 802 16 806
rect 20 802 22 806
rect 14 800 22 802
rect 223 807 231 809
rect 223 803 225 807
rect 229 803 231 807
rect 223 801 231 803
rect 233 807 241 809
rect 233 803 235 807
rect 239 803 241 807
rect 233 801 241 803
rect 243 807 251 809
rect 243 803 245 807
rect 249 803 251 807
rect 243 801 251 803
rect 551 807 559 809
rect 551 803 553 807
rect 557 803 559 807
rect 551 801 559 803
rect 561 807 569 809
rect 561 803 563 807
rect 567 803 569 807
rect 561 801 569 803
rect 571 807 579 809
rect 571 803 573 807
rect 577 803 579 807
rect 590 807 592 811
rect 596 807 598 811
rect 590 805 598 807
rect 571 801 579 803
rect 590 801 598 803
rect 2 796 10 798
rect 14 796 22 798
rect 2 792 10 794
rect 2 788 4 792
rect 8 788 10 792
rect 14 792 16 796
rect 20 792 22 796
rect 14 790 22 792
rect 223 797 231 799
rect 223 793 225 797
rect 229 793 231 797
rect 223 791 231 793
rect 233 797 241 799
rect 233 793 235 797
rect 239 793 241 797
rect 233 791 241 793
rect 243 797 251 799
rect 243 793 245 797
rect 249 793 251 797
rect 243 791 251 793
rect 387 797 395 799
rect 387 793 389 797
rect 393 793 395 797
rect 387 791 395 793
rect 397 797 405 799
rect 397 793 399 797
rect 403 793 405 797
rect 397 791 405 793
rect 407 797 415 799
rect 407 793 409 797
rect 413 793 415 797
rect 407 791 415 793
rect 551 797 559 799
rect 551 793 553 797
rect 557 793 559 797
rect 551 791 559 793
rect 561 797 569 799
rect 561 793 563 797
rect 567 793 569 797
rect 561 791 569 793
rect 571 797 579 799
rect 571 793 573 797
rect 577 793 579 797
rect 590 797 592 801
rect 596 797 598 801
rect 590 795 598 797
rect 571 791 579 793
rect 590 791 598 793
rect 2 786 10 788
rect 387 787 395 789
rect 14 784 22 786
rect 2 782 10 784
rect 2 778 4 782
rect 8 778 10 782
rect 14 780 16 784
rect 20 780 22 784
rect 387 783 389 787
rect 393 783 395 787
rect 387 781 395 783
rect 397 787 405 789
rect 397 783 399 787
rect 403 783 405 787
rect 397 781 405 783
rect 407 787 415 789
rect 407 783 409 787
rect 413 783 415 787
rect 590 787 592 791
rect 596 787 598 791
rect 590 785 598 787
rect 407 781 415 783
rect 576 782 584 784
rect 14 778 22 780
rect 576 778 578 782
rect 582 778 584 782
rect 2 776 10 778
rect 50 776 58 778
rect 14 774 22 776
rect 2 772 10 774
rect 2 768 4 772
rect 8 768 10 772
rect 14 770 16 774
rect 20 770 22 774
rect 50 772 52 776
rect 56 772 58 776
rect 50 770 58 772
rect 60 776 68 778
rect 576 776 584 778
rect 590 781 598 783
rect 590 777 592 781
rect 596 777 598 781
rect 60 772 62 776
rect 66 772 68 776
rect 590 775 598 777
rect 60 770 68 772
rect 590 771 598 773
rect 14 768 22 770
rect 2 766 10 768
rect 590 767 592 771
rect 596 767 598 771
rect 14 764 22 766
rect 590 765 598 767
rect 2 762 10 764
rect 2 758 4 762
rect 8 758 10 762
rect 14 760 16 764
rect 20 760 22 764
rect 286 761 294 763
rect 14 758 22 760
rect 28 758 36 760
rect 2 756 10 758
rect 14 754 22 756
rect 2 752 10 754
rect 2 748 4 752
rect 8 748 10 752
rect 14 750 16 754
rect 20 750 22 754
rect 28 754 30 758
rect 34 754 36 758
rect 28 752 36 754
rect 44 758 52 760
rect 44 754 46 758
rect 50 754 52 758
rect 44 752 52 754
rect 60 756 68 758
rect 60 752 62 756
rect 66 752 68 756
rect 60 750 68 752
rect 78 757 86 759
rect 78 753 80 757
rect 84 753 86 757
rect 110 757 118 759
rect 78 751 86 753
rect 94 754 102 756
rect 94 750 96 754
rect 100 750 102 754
rect 110 753 112 757
rect 116 753 118 757
rect 142 757 150 759
rect 110 751 118 753
rect 126 754 134 756
rect 14 748 22 750
rect 28 748 36 750
rect 2 746 10 748
rect 14 744 22 746
rect 2 742 10 744
rect 2 738 4 742
rect 8 738 10 742
rect 14 740 16 744
rect 20 740 22 744
rect 28 744 30 748
rect 34 744 36 748
rect 28 742 36 744
rect 44 748 52 750
rect 44 744 46 748
rect 50 744 52 748
rect 44 742 52 744
rect 60 746 68 748
rect 60 742 62 746
rect 66 742 68 746
rect 60 740 68 742
rect 78 747 86 749
rect 94 748 102 750
rect 126 750 128 754
rect 132 750 134 754
rect 142 753 144 757
rect 148 753 150 757
rect 174 757 182 759
rect 142 751 150 753
rect 158 754 166 756
rect 78 743 80 747
rect 84 743 86 747
rect 110 747 118 749
rect 126 748 134 750
rect 158 750 160 754
rect 164 750 166 754
rect 174 753 176 757
rect 180 753 182 757
rect 206 758 214 760
rect 174 751 182 753
rect 190 754 198 756
rect 78 741 86 743
rect 94 744 102 746
rect 94 740 96 744
rect 100 740 102 744
rect 110 743 112 747
rect 116 743 118 747
rect 142 747 150 749
rect 158 748 166 750
rect 190 750 192 754
rect 196 750 198 754
rect 206 754 208 758
rect 212 754 214 758
rect 238 756 246 758
rect 270 756 278 758
rect 206 752 214 754
rect 222 754 230 756
rect 222 750 224 754
rect 228 750 230 754
rect 238 752 240 756
rect 244 752 246 756
rect 238 750 246 752
rect 254 754 262 756
rect 254 750 256 754
rect 260 750 262 754
rect 270 752 272 756
rect 276 752 278 756
rect 286 757 288 761
rect 292 757 294 761
rect 286 755 294 757
rect 302 762 310 764
rect 302 758 304 762
rect 308 758 310 762
rect 590 761 598 763
rect 302 756 310 758
rect 386 758 394 760
rect 386 754 388 758
rect 392 754 394 758
rect 386 752 394 754
rect 402 758 410 760
rect 402 754 404 758
rect 408 754 410 758
rect 402 752 410 754
rect 434 758 442 760
rect 434 754 436 758
rect 440 754 442 758
rect 434 752 442 754
rect 450 759 458 761
rect 450 755 452 759
rect 456 755 458 759
rect 450 753 458 755
rect 466 759 474 761
rect 466 755 468 759
rect 472 755 474 759
rect 466 753 474 755
rect 482 759 490 761
rect 482 755 484 759
rect 488 755 490 759
rect 482 753 490 755
rect 498 759 506 761
rect 498 755 500 759
rect 504 755 506 759
rect 498 753 506 755
rect 514 759 522 761
rect 514 755 516 759
rect 520 755 522 759
rect 514 753 522 755
rect 530 759 538 761
rect 530 755 532 759
rect 536 755 538 759
rect 530 753 538 755
rect 546 759 554 761
rect 546 755 548 759
rect 552 755 554 759
rect 546 753 554 755
rect 562 759 570 761
rect 562 755 564 759
rect 568 755 570 759
rect 562 753 570 755
rect 578 759 586 761
rect 578 755 580 759
rect 584 755 586 759
rect 590 757 592 761
rect 596 757 598 761
rect 590 755 598 757
rect 578 753 586 755
rect 270 750 278 752
rect 286 750 294 752
rect 110 741 118 743
rect 126 744 134 746
rect 14 738 22 740
rect 28 738 36 740
rect 2 736 10 738
rect 14 734 22 736
rect 2 732 10 734
rect 2 728 4 732
rect 8 728 10 732
rect 14 730 16 734
rect 20 730 22 734
rect 28 734 30 738
rect 34 734 36 738
rect 28 732 36 734
rect 44 738 52 740
rect 44 734 46 738
rect 50 734 52 738
rect 44 732 52 734
rect 60 736 68 738
rect 60 732 62 736
rect 66 732 68 736
rect 60 730 68 732
rect 78 737 86 739
rect 94 738 102 740
rect 126 740 128 744
rect 132 740 134 744
rect 142 743 144 747
rect 148 743 150 747
rect 174 747 182 749
rect 190 748 198 750
rect 206 748 214 750
rect 222 748 230 750
rect 254 748 262 750
rect 142 741 150 743
rect 158 744 166 746
rect 78 733 80 737
rect 84 733 86 737
rect 110 737 118 739
rect 126 738 134 740
rect 158 740 160 744
rect 164 740 166 744
rect 174 743 176 747
rect 180 743 182 747
rect 174 741 182 743
rect 190 744 198 746
rect 78 731 86 733
rect 94 734 102 736
rect 94 730 96 734
rect 100 730 102 734
rect 110 733 112 737
rect 116 733 118 737
rect 142 737 150 739
rect 158 738 166 740
rect 190 740 192 744
rect 196 740 198 744
rect 206 744 208 748
rect 212 744 214 748
rect 238 746 246 748
rect 270 746 278 748
rect 206 742 214 744
rect 222 744 230 746
rect 222 740 224 744
rect 228 740 230 744
rect 238 742 240 746
rect 244 742 246 746
rect 238 740 246 742
rect 254 744 262 746
rect 254 740 256 744
rect 260 740 262 744
rect 270 742 272 746
rect 276 742 278 746
rect 286 746 288 750
rect 292 746 294 750
rect 286 744 294 746
rect 302 750 310 752
rect 590 751 598 753
rect 302 746 304 750
rect 308 746 310 750
rect 302 744 310 746
rect 386 748 394 750
rect 386 744 388 748
rect 392 744 394 748
rect 386 742 394 744
rect 402 748 410 750
rect 434 748 442 750
rect 402 744 404 748
rect 408 744 410 748
rect 402 742 410 744
rect 418 746 426 748
rect 418 742 420 746
rect 424 742 426 746
rect 434 744 436 748
rect 440 744 442 748
rect 434 742 442 744
rect 450 749 458 751
rect 450 745 452 749
rect 456 745 458 749
rect 450 743 458 745
rect 466 749 474 751
rect 466 745 468 749
rect 472 745 474 749
rect 466 743 474 745
rect 482 749 490 751
rect 482 745 484 749
rect 488 745 490 749
rect 482 743 490 745
rect 498 749 506 751
rect 498 745 500 749
rect 504 745 506 749
rect 498 743 506 745
rect 514 749 522 751
rect 514 745 516 749
rect 520 745 522 749
rect 514 743 522 745
rect 530 749 538 751
rect 530 745 532 749
rect 536 745 538 749
rect 530 743 538 745
rect 546 749 554 751
rect 546 745 548 749
rect 552 745 554 749
rect 546 743 554 745
rect 562 749 570 751
rect 562 745 564 749
rect 568 745 570 749
rect 562 743 570 745
rect 578 749 586 751
rect 578 745 580 749
rect 584 745 586 749
rect 590 747 592 751
rect 596 747 598 751
rect 590 745 598 747
rect 578 743 586 745
rect 270 740 278 742
rect 110 731 118 733
rect 126 734 134 736
rect 14 728 22 730
rect 28 728 36 730
rect 2 726 10 728
rect 14 724 22 726
rect 2 722 10 724
rect 2 718 4 722
rect 8 718 10 722
rect 14 720 16 724
rect 20 720 22 724
rect 28 724 30 728
rect 34 724 36 728
rect 28 722 36 724
rect 44 728 52 730
rect 44 724 46 728
rect 50 724 52 728
rect 44 722 52 724
rect 60 726 68 728
rect 60 722 62 726
rect 66 722 68 726
rect 60 720 68 722
rect 78 727 86 729
rect 94 728 102 730
rect 126 730 128 734
rect 132 730 134 734
rect 142 733 144 737
rect 148 733 150 737
rect 174 737 182 739
rect 190 738 198 740
rect 206 738 214 740
rect 222 738 230 740
rect 254 738 262 740
rect 286 738 294 740
rect 142 731 150 733
rect 158 734 166 736
rect 78 723 80 727
rect 84 723 86 727
rect 110 727 118 729
rect 126 728 134 730
rect 158 730 160 734
rect 164 730 166 734
rect 174 733 176 737
rect 180 733 182 737
rect 174 731 182 733
rect 190 734 198 736
rect 78 721 86 723
rect 94 724 102 726
rect 94 720 96 724
rect 100 720 102 724
rect 110 723 112 727
rect 116 723 118 727
rect 142 727 150 729
rect 158 728 166 730
rect 190 730 192 734
rect 196 730 198 734
rect 206 734 208 738
rect 212 734 214 738
rect 238 736 246 738
rect 270 736 278 738
rect 206 732 214 734
rect 222 734 230 736
rect 222 730 224 734
rect 228 730 230 734
rect 238 732 240 736
rect 244 732 246 736
rect 238 730 246 732
rect 254 734 262 736
rect 254 730 256 734
rect 260 730 262 734
rect 270 732 272 736
rect 276 732 278 736
rect 286 734 288 738
rect 292 734 294 738
rect 286 732 294 734
rect 302 739 310 741
rect 418 740 426 742
rect 590 741 598 743
rect 302 735 304 739
rect 308 735 310 739
rect 302 733 310 735
rect 386 738 394 740
rect 386 734 388 738
rect 392 734 394 738
rect 386 732 394 734
rect 402 738 410 740
rect 434 738 442 740
rect 402 734 404 738
rect 408 734 410 738
rect 402 732 410 734
rect 418 736 426 738
rect 418 732 420 736
rect 424 732 426 736
rect 434 734 436 738
rect 440 734 442 738
rect 434 732 442 734
rect 450 739 458 741
rect 450 735 452 739
rect 456 735 458 739
rect 450 733 458 735
rect 466 739 474 741
rect 466 735 468 739
rect 472 735 474 739
rect 466 733 474 735
rect 482 739 490 741
rect 482 735 484 739
rect 488 735 490 739
rect 482 733 490 735
rect 498 739 506 741
rect 498 735 500 739
rect 504 735 506 739
rect 498 733 506 735
rect 514 739 522 741
rect 514 735 516 739
rect 520 735 522 739
rect 514 733 522 735
rect 530 739 538 741
rect 530 735 532 739
rect 536 735 538 739
rect 530 733 538 735
rect 546 739 554 741
rect 546 735 548 739
rect 552 735 554 739
rect 546 733 554 735
rect 562 739 570 741
rect 562 735 564 739
rect 568 735 570 739
rect 562 733 570 735
rect 578 739 586 741
rect 578 735 580 739
rect 584 735 586 739
rect 590 737 592 741
rect 596 737 598 741
rect 590 735 598 737
rect 578 733 586 735
rect 270 730 278 732
rect 418 730 426 732
rect 590 731 598 733
rect 110 721 118 723
rect 126 724 134 726
rect 14 718 22 720
rect 44 718 52 720
rect 94 718 102 720
rect 126 720 128 724
rect 132 720 134 724
rect 142 723 144 727
rect 148 723 150 727
rect 174 727 182 729
rect 190 728 198 730
rect 206 728 214 730
rect 222 728 230 730
rect 254 728 262 730
rect 386 728 394 730
rect 142 721 150 723
rect 158 724 166 726
rect 2 716 10 718
rect 14 714 22 716
rect 2 712 10 714
rect 2 708 4 712
rect 8 708 10 712
rect 14 710 16 714
rect 20 710 22 714
rect 44 714 46 718
rect 50 714 52 718
rect 44 712 52 714
rect 60 716 68 718
rect 110 717 118 719
rect 126 718 134 720
rect 158 720 160 724
rect 164 720 166 724
rect 174 723 176 727
rect 180 723 182 727
rect 174 721 182 723
rect 190 724 198 726
rect 60 712 62 716
rect 66 712 68 716
rect 60 710 68 712
rect 94 714 102 716
rect 94 710 96 714
rect 100 710 102 714
rect 110 713 112 717
rect 116 713 118 717
rect 142 717 150 719
rect 158 718 166 720
rect 190 720 192 724
rect 196 720 198 724
rect 206 724 208 728
rect 212 724 214 728
rect 238 726 246 728
rect 270 726 278 728
rect 206 722 214 724
rect 222 724 230 726
rect 222 720 224 724
rect 228 720 230 724
rect 238 722 240 726
rect 244 722 246 726
rect 238 720 246 722
rect 254 724 262 726
rect 254 720 256 724
rect 260 720 262 724
rect 270 722 272 726
rect 276 722 278 726
rect 270 720 278 722
rect 286 726 294 728
rect 286 722 288 726
rect 292 722 294 726
rect 286 720 294 722
rect 302 726 310 728
rect 302 722 304 726
rect 308 722 310 726
rect 386 724 388 728
rect 392 724 394 728
rect 386 722 394 724
rect 402 728 410 730
rect 434 728 442 730
rect 402 724 404 728
rect 408 724 410 728
rect 402 722 410 724
rect 418 726 426 728
rect 418 722 420 726
rect 424 722 426 726
rect 434 724 436 728
rect 440 724 442 728
rect 434 722 442 724
rect 450 729 458 731
rect 450 725 452 729
rect 456 725 458 729
rect 450 723 458 725
rect 466 729 474 731
rect 466 725 468 729
rect 472 725 474 729
rect 466 723 474 725
rect 482 729 490 731
rect 482 725 484 729
rect 488 725 490 729
rect 482 723 490 725
rect 498 729 506 731
rect 498 725 500 729
rect 504 725 506 729
rect 498 723 506 725
rect 514 729 522 731
rect 514 725 516 729
rect 520 725 522 729
rect 514 723 522 725
rect 530 729 538 731
rect 530 725 532 729
rect 536 725 538 729
rect 530 723 538 725
rect 546 729 554 731
rect 546 725 548 729
rect 552 725 554 729
rect 546 723 554 725
rect 562 729 570 731
rect 562 725 564 729
rect 568 725 570 729
rect 562 723 570 725
rect 578 729 586 731
rect 578 725 580 729
rect 584 725 586 729
rect 590 727 592 731
rect 596 727 598 731
rect 590 725 598 727
rect 578 723 586 725
rect 302 720 310 722
rect 418 720 426 722
rect 590 721 598 723
rect 110 711 118 713
rect 126 714 134 716
rect 14 708 22 710
rect 94 708 102 710
rect 126 710 128 714
rect 132 710 134 714
rect 142 713 144 717
rect 148 713 150 717
rect 174 717 182 719
rect 190 718 198 720
rect 206 718 214 720
rect 222 718 230 720
rect 254 718 262 720
rect 386 718 394 720
rect 142 711 150 713
rect 158 714 166 716
rect 126 708 134 710
rect 158 710 160 714
rect 164 710 166 714
rect 174 713 176 717
rect 180 713 182 717
rect 174 711 182 713
rect 190 714 198 716
rect 158 708 166 710
rect 190 710 192 714
rect 196 710 198 714
rect 206 714 208 718
rect 212 714 214 718
rect 270 716 278 718
rect 206 712 214 714
rect 222 714 230 716
rect 190 708 198 710
rect 222 710 224 714
rect 228 710 230 714
rect 222 708 230 710
rect 254 714 262 716
rect 254 710 256 714
rect 260 710 262 714
rect 270 712 272 716
rect 276 712 278 716
rect 270 710 278 712
rect 302 714 310 716
rect 302 710 304 714
rect 308 710 310 714
rect 386 714 388 718
rect 392 714 394 718
rect 386 712 394 714
rect 402 718 410 720
rect 402 714 404 718
rect 408 714 410 718
rect 434 718 442 720
rect 402 712 410 714
rect 418 715 426 717
rect 254 708 262 710
rect 302 708 310 710
rect 418 711 420 715
rect 424 711 426 715
rect 434 714 436 718
rect 440 714 442 718
rect 434 712 442 714
rect 450 719 458 721
rect 450 715 452 719
rect 456 715 458 719
rect 450 713 458 715
rect 466 719 474 721
rect 466 715 468 719
rect 472 715 474 719
rect 466 713 474 715
rect 482 719 490 721
rect 482 715 484 719
rect 488 715 490 719
rect 482 713 490 715
rect 498 719 506 721
rect 498 715 500 719
rect 504 715 506 719
rect 498 713 506 715
rect 514 719 522 721
rect 514 715 516 719
rect 520 715 522 719
rect 514 713 522 715
rect 530 719 538 721
rect 530 715 532 719
rect 536 715 538 719
rect 530 713 538 715
rect 546 719 554 721
rect 546 715 548 719
rect 552 715 554 719
rect 546 713 554 715
rect 562 719 570 721
rect 562 715 564 719
rect 568 715 570 719
rect 562 713 570 715
rect 578 719 586 721
rect 578 715 580 719
rect 584 715 586 719
rect 590 717 592 721
rect 596 717 598 721
rect 590 715 598 717
rect 578 713 586 715
rect 418 709 426 711
rect 590 711 598 713
rect 2 706 10 708
rect 590 707 592 711
rect 596 707 598 711
rect 590 705 598 707
rect 2 702 10 704
rect 580 703 588 705
rect 2 698 4 702
rect 8 698 10 702
rect 2 696 10 698
rect 18 700 26 702
rect 18 696 20 700
rect 24 696 26 700
rect 18 694 26 696
rect 50 700 58 702
rect 50 696 52 700
rect 56 696 58 700
rect 50 694 58 696
rect 104 699 112 701
rect 104 695 106 699
rect 110 695 112 699
rect 2 692 10 694
rect 2 688 4 692
rect 8 688 10 692
rect 2 686 10 688
rect 34 692 42 694
rect 104 693 112 695
rect 114 699 122 701
rect 114 695 116 699
rect 120 695 122 699
rect 114 693 122 695
rect 172 700 180 702
rect 172 696 174 700
rect 178 696 180 700
rect 172 694 180 696
rect 182 700 190 702
rect 182 696 184 700
rect 188 696 190 700
rect 182 694 190 696
rect 274 700 282 702
rect 274 696 276 700
rect 280 696 282 700
rect 198 693 214 695
rect 34 688 36 692
rect 40 688 42 692
rect 34 686 42 688
rect 76 691 84 693
rect 76 687 78 691
rect 82 687 84 691
rect 76 685 84 687
rect 90 691 98 693
rect 90 687 92 691
rect 96 687 98 691
rect 90 685 98 687
rect 128 691 136 693
rect 128 687 130 691
rect 134 687 136 691
rect 128 685 136 687
rect 138 691 146 693
rect 138 687 140 691
rect 144 687 146 691
rect 138 685 146 687
rect 148 691 156 693
rect 148 687 150 691
rect 154 687 156 691
rect 148 685 156 687
rect 158 691 166 693
rect 158 687 160 691
rect 164 687 166 691
rect 198 689 200 693
rect 204 689 208 693
rect 212 689 214 693
rect 198 687 214 689
rect 216 693 224 695
rect 216 689 218 693
rect 222 689 224 693
rect 216 687 224 689
rect 248 693 256 695
rect 248 689 250 693
rect 254 689 256 693
rect 248 687 256 689
rect 260 693 268 695
rect 274 694 282 696
rect 284 700 292 702
rect 284 696 286 700
rect 290 696 292 700
rect 284 694 292 696
rect 460 701 468 703
rect 460 697 462 701
rect 466 697 468 701
rect 460 695 468 697
rect 470 701 478 703
rect 470 697 472 701
rect 476 697 478 701
rect 470 695 478 697
rect 556 701 564 703
rect 556 697 558 701
rect 562 697 564 701
rect 556 695 564 697
rect 566 701 574 703
rect 566 697 568 701
rect 572 697 574 701
rect 580 699 582 703
rect 586 699 588 703
rect 580 697 588 699
rect 590 701 598 703
rect 590 697 592 701
rect 596 697 598 701
rect 566 695 574 697
rect 590 695 598 697
rect 260 689 262 693
rect 266 689 268 693
rect 260 687 268 689
rect 388 691 396 693
rect 388 687 390 691
rect 394 687 396 691
rect 158 685 166 687
rect 388 685 396 687
rect 398 691 406 693
rect 398 687 400 691
rect 404 687 406 691
rect 398 685 406 687
rect 408 691 416 693
rect 408 687 410 691
rect 414 687 416 691
rect 408 685 416 687
rect 418 691 426 693
rect 418 687 420 691
rect 424 687 426 691
rect 418 685 426 687
rect 446 692 454 694
rect 446 688 448 692
rect 452 688 454 692
rect 446 686 454 688
rect 484 691 492 693
rect 484 687 486 691
rect 490 687 492 691
rect 484 685 492 687
rect 494 691 502 693
rect 494 687 496 691
rect 500 687 502 691
rect 494 685 502 687
rect 504 691 512 693
rect 504 687 506 691
rect 510 687 512 691
rect 504 685 512 687
rect 514 691 522 693
rect 514 687 516 691
rect 520 687 522 691
rect 514 685 522 687
rect 542 690 550 692
rect 542 686 544 690
rect 548 686 550 690
rect 542 684 550 686
rect 580 691 588 693
rect 580 687 582 691
rect 586 687 588 691
rect 580 685 588 687
rect 590 691 598 693
rect 590 687 592 691
rect 596 687 598 691
rect 590 685 598 687
rect 388 679 396 681
rect 40 676 48 678
rect 40 672 42 676
rect 46 672 48 676
rect 40 670 48 672
rect 50 676 58 678
rect 50 672 52 676
rect 56 672 58 676
rect 50 670 58 672
rect 64 676 72 678
rect 64 672 66 676
rect 70 672 72 676
rect 64 670 72 672
rect 74 676 82 678
rect 74 672 76 676
rect 80 672 82 676
rect 74 670 82 672
rect 160 676 168 678
rect 160 672 162 676
rect 166 672 168 676
rect 160 670 168 672
rect 170 676 178 678
rect 170 672 172 676
rect 176 672 178 676
rect 170 670 178 672
rect 184 676 192 678
rect 184 672 186 676
rect 190 672 192 676
rect 184 670 192 672
rect 194 676 202 678
rect 194 672 196 676
rect 200 672 202 676
rect 194 670 202 672
rect 248 676 256 678
rect 248 672 250 676
rect 254 672 256 676
rect 248 670 256 672
rect 258 676 266 678
rect 258 672 260 676
rect 264 672 266 676
rect 258 670 266 672
rect 274 676 282 678
rect 274 672 276 676
rect 280 672 282 676
rect 274 670 282 672
rect 284 676 292 678
rect 284 672 286 676
rect 290 672 292 676
rect 388 675 390 679
rect 394 675 396 679
rect 388 673 396 675
rect 398 679 406 681
rect 398 675 400 679
rect 404 675 406 679
rect 398 673 406 675
rect 408 679 416 681
rect 408 675 410 679
rect 414 675 416 679
rect 408 673 416 675
rect 418 679 426 681
rect 418 675 420 679
rect 424 675 426 679
rect 418 673 426 675
rect 434 676 442 678
rect 284 670 292 672
rect 434 672 436 676
rect 440 672 442 676
rect 434 670 442 672
rect 444 676 452 678
rect 444 672 446 676
rect 450 672 452 676
rect 444 670 452 672
rect 555 676 563 678
rect 555 672 557 676
rect 561 672 563 676
rect 555 670 563 672
rect 565 676 573 678
rect 565 672 567 676
rect 571 672 573 676
rect 565 670 573 672
rect 2 660 10 662
rect 2 656 4 660
rect 8 656 10 660
rect 2 654 10 656
rect 34 661 42 663
rect 34 657 36 661
rect 40 657 42 661
rect 34 655 42 657
rect 76 661 84 663
rect 76 657 78 661
rect 82 657 84 661
rect 76 655 84 657
rect 90 661 98 663
rect 90 657 92 661
rect 96 657 98 661
rect 90 655 98 657
rect 128 661 136 663
rect 128 657 130 661
rect 134 657 136 661
rect 128 655 136 657
rect 138 661 146 663
rect 138 657 140 661
rect 144 657 146 661
rect 138 655 146 657
rect 148 661 156 663
rect 148 657 150 661
rect 154 657 156 661
rect 148 655 156 657
rect 158 661 166 663
rect 158 657 160 661
rect 164 657 166 661
rect 158 655 166 657
rect 196 661 204 663
rect 196 657 198 661
rect 202 657 204 661
rect 196 655 204 657
rect 208 661 216 663
rect 208 657 210 661
rect 214 657 216 661
rect 208 655 216 657
rect 218 661 226 663
rect 218 657 220 661
rect 224 657 226 661
rect 218 655 226 657
rect 274 661 282 663
rect 274 657 276 661
rect 280 657 282 661
rect 274 655 282 657
rect 284 661 292 663
rect 284 657 286 661
rect 290 657 292 661
rect 284 655 292 657
rect 388 661 396 663
rect 388 657 390 661
rect 394 657 396 661
rect 388 655 396 657
rect 398 661 406 663
rect 398 657 400 661
rect 404 657 406 661
rect 398 655 406 657
rect 408 661 416 663
rect 408 657 410 661
rect 414 657 416 661
rect 408 655 416 657
rect 418 661 426 663
rect 418 657 420 661
rect 424 657 426 661
rect 418 655 426 657
rect 446 661 454 663
rect 446 657 448 661
rect 452 657 454 661
rect 446 655 454 657
rect 484 661 492 663
rect 484 657 486 661
rect 490 657 492 661
rect 484 655 492 657
rect 494 661 502 663
rect 494 657 496 661
rect 500 657 502 661
rect 494 655 502 657
rect 504 661 512 663
rect 504 657 506 661
rect 510 657 512 661
rect 504 655 512 657
rect 514 661 522 663
rect 514 657 516 661
rect 520 657 522 661
rect 514 655 522 657
rect 542 661 550 663
rect 542 657 544 661
rect 548 657 550 661
rect 542 655 550 657
rect 580 662 588 664
rect 580 658 582 662
rect 586 658 588 662
rect 580 656 588 658
rect 590 662 598 664
rect 590 658 592 662
rect 596 658 598 662
rect 590 656 598 658
rect 18 653 26 655
rect 2 650 10 652
rect 2 646 4 650
rect 8 646 10 650
rect 18 649 20 653
rect 24 649 26 653
rect 18 647 26 649
rect 50 653 58 655
rect 50 649 52 653
rect 56 649 58 653
rect 50 647 58 649
rect 104 653 112 655
rect 104 649 106 653
rect 110 649 112 653
rect 104 647 112 649
rect 114 653 122 655
rect 114 649 116 653
rect 120 649 122 653
rect 114 647 122 649
rect 172 653 180 655
rect 172 649 174 653
rect 178 649 180 653
rect 172 647 180 649
rect 182 653 190 655
rect 182 649 184 653
rect 188 649 190 653
rect 182 647 190 649
rect 248 653 256 655
rect 248 649 250 653
rect 254 649 256 653
rect 248 647 256 649
rect 258 653 266 655
rect 258 649 260 653
rect 264 649 266 653
rect 258 647 266 649
rect 460 653 468 655
rect 460 649 462 653
rect 466 649 468 653
rect 460 647 468 649
rect 470 653 478 655
rect 470 649 472 653
rect 476 649 478 653
rect 470 647 478 649
rect 556 653 564 655
rect 556 649 558 653
rect 562 649 564 653
rect 556 647 564 649
rect 566 653 574 655
rect 566 649 568 653
rect 572 649 574 653
rect 566 647 574 649
rect 590 652 598 654
rect 590 648 592 652
rect 596 648 598 652
rect 590 646 598 648
rect 2 644 10 646
rect 590 642 598 644
rect 2 640 10 642
rect 2 636 4 640
rect 8 636 10 640
rect 44 639 52 641
rect 94 639 102 641
rect 2 634 10 636
rect 14 634 22 636
rect 2 630 10 632
rect 2 626 4 630
rect 8 626 10 630
rect 14 630 16 634
rect 20 630 22 634
rect 44 635 46 639
rect 50 635 52 639
rect 44 633 52 635
rect 60 637 68 639
rect 60 633 62 637
rect 66 633 68 637
rect 94 635 96 639
rect 100 635 102 639
rect 94 633 102 635
rect 110 637 118 639
rect 110 633 112 637
rect 116 633 118 637
rect 142 637 150 639
rect 142 633 144 637
rect 148 633 150 637
rect 174 638 182 640
rect 222 639 230 641
rect 174 634 176 638
rect 180 634 182 638
rect 60 631 68 633
rect 110 631 118 633
rect 126 631 134 633
rect 142 631 150 633
rect 158 631 166 633
rect 174 632 182 634
rect 206 637 214 639
rect 206 633 208 637
rect 212 633 214 637
rect 222 635 224 639
rect 228 635 230 639
rect 222 633 230 635
rect 238 638 246 640
rect 238 634 240 638
rect 244 634 246 638
rect 14 628 22 630
rect 44 629 52 631
rect 94 629 102 631
rect 28 627 36 629
rect 2 624 10 626
rect 14 624 22 626
rect 2 620 10 622
rect 2 616 4 620
rect 8 616 10 620
rect 14 620 16 624
rect 20 620 22 624
rect 28 623 30 627
rect 34 623 36 627
rect 44 625 46 629
rect 50 625 52 629
rect 44 623 52 625
rect 60 627 68 629
rect 60 623 62 627
rect 66 623 68 627
rect 28 621 36 623
rect 60 621 68 623
rect 78 627 86 629
rect 78 623 80 627
rect 84 623 86 627
rect 94 625 96 629
rect 100 625 102 629
rect 94 623 102 625
rect 110 627 118 629
rect 110 623 112 627
rect 116 623 118 627
rect 126 627 128 631
rect 132 627 134 631
rect 126 625 134 627
rect 142 627 150 629
rect 142 623 144 627
rect 148 623 150 627
rect 158 627 160 631
rect 164 627 166 631
rect 190 631 198 633
rect 206 631 214 633
rect 238 632 246 634
rect 270 638 278 640
rect 270 634 272 638
rect 276 634 278 638
rect 270 632 278 634
rect 286 639 294 641
rect 286 635 288 639
rect 292 635 294 639
rect 590 638 592 642
rect 596 638 598 642
rect 590 636 598 638
rect 286 633 294 635
rect 386 631 394 633
rect 158 625 166 627
rect 174 628 182 630
rect 174 624 176 628
rect 180 624 182 628
rect 190 627 192 631
rect 196 627 198 631
rect 222 629 230 631
rect 190 625 198 627
rect 206 627 214 629
rect 78 621 86 623
rect 110 621 118 623
rect 126 621 134 623
rect 142 621 150 623
rect 158 621 166 623
rect 174 622 182 624
rect 206 623 208 627
rect 212 623 214 627
rect 222 625 224 629
rect 228 625 230 629
rect 222 623 230 625
rect 238 628 246 630
rect 286 629 294 631
rect 238 624 240 628
rect 244 624 246 628
rect 14 618 22 620
rect 44 619 52 621
rect 94 619 102 621
rect 28 617 36 619
rect 2 614 10 616
rect 14 614 22 616
rect 2 610 10 612
rect 2 606 4 610
rect 8 606 10 610
rect 14 610 16 614
rect 20 610 22 614
rect 28 613 30 617
rect 34 613 36 617
rect 44 615 46 619
rect 50 615 52 619
rect 44 613 52 615
rect 60 617 68 619
rect 60 613 62 617
rect 66 613 68 617
rect 28 611 36 613
rect 60 611 68 613
rect 78 617 86 619
rect 78 613 80 617
rect 84 613 86 617
rect 94 615 96 619
rect 100 615 102 619
rect 94 613 102 615
rect 110 617 118 619
rect 110 613 112 617
rect 116 613 118 617
rect 126 617 128 621
rect 132 617 134 621
rect 126 615 134 617
rect 142 617 150 619
rect 142 613 144 617
rect 148 613 150 617
rect 158 617 160 621
rect 164 617 166 621
rect 190 621 198 623
rect 206 621 214 623
rect 238 622 246 624
rect 270 627 278 629
rect 270 623 272 627
rect 276 623 278 627
rect 286 625 288 629
rect 292 625 294 629
rect 286 623 294 625
rect 302 627 310 629
rect 302 623 304 627
rect 308 623 310 627
rect 386 627 388 631
rect 392 627 394 631
rect 386 625 394 627
rect 402 631 410 633
rect 402 627 404 631
rect 408 627 410 631
rect 402 625 410 627
rect 418 631 426 633
rect 418 627 420 631
rect 424 627 426 631
rect 418 625 426 627
rect 434 631 442 633
rect 434 627 436 631
rect 440 627 442 631
rect 434 625 442 627
rect 450 631 458 633
rect 450 627 452 631
rect 456 627 458 631
rect 450 625 458 627
rect 466 631 474 633
rect 466 627 468 631
rect 472 627 474 631
rect 466 625 474 627
rect 482 631 490 633
rect 482 627 484 631
rect 488 627 490 631
rect 482 625 490 627
rect 498 631 506 633
rect 498 627 500 631
rect 504 627 506 631
rect 498 625 506 627
rect 514 631 522 633
rect 514 627 516 631
rect 520 627 522 631
rect 514 625 522 627
rect 530 631 538 633
rect 530 627 532 631
rect 536 627 538 631
rect 530 625 538 627
rect 546 631 554 633
rect 546 627 548 631
rect 552 627 554 631
rect 546 625 554 627
rect 562 631 570 633
rect 562 627 564 631
rect 568 627 570 631
rect 562 625 570 627
rect 578 631 586 633
rect 578 627 580 631
rect 584 627 586 631
rect 578 625 586 627
rect 590 632 598 634
rect 590 628 592 632
rect 596 628 598 632
rect 590 626 598 628
rect 254 621 262 623
rect 270 621 278 623
rect 302 621 310 623
rect 386 621 394 623
rect 158 615 166 617
rect 174 618 182 620
rect 174 614 176 618
rect 180 614 182 618
rect 190 617 192 621
rect 196 617 198 621
rect 222 619 230 621
rect 190 615 198 617
rect 206 617 214 619
rect 78 611 86 613
rect 110 611 118 613
rect 126 611 134 613
rect 142 611 150 613
rect 158 611 166 613
rect 174 612 182 614
rect 206 613 208 617
rect 212 613 214 617
rect 222 615 224 619
rect 228 615 230 619
rect 222 613 230 615
rect 238 618 246 620
rect 238 614 240 618
rect 244 614 246 618
rect 254 617 256 621
rect 260 617 262 621
rect 254 615 262 617
rect 286 619 294 621
rect 286 615 288 619
rect 292 615 294 619
rect 14 608 22 610
rect 44 609 52 611
rect 94 609 102 611
rect 28 607 36 609
rect 2 604 10 606
rect 14 604 22 606
rect 2 600 10 602
rect 2 596 4 600
rect 8 596 10 600
rect 14 600 16 604
rect 20 600 22 604
rect 28 603 30 607
rect 34 603 36 607
rect 44 605 46 609
rect 50 605 52 609
rect 44 603 52 605
rect 60 607 68 609
rect 60 603 62 607
rect 66 603 68 607
rect 28 601 36 603
rect 60 601 68 603
rect 78 607 86 609
rect 78 603 80 607
rect 84 603 86 607
rect 94 605 96 609
rect 100 605 102 609
rect 94 603 102 605
rect 110 607 118 609
rect 110 603 112 607
rect 116 603 118 607
rect 126 607 128 611
rect 132 607 134 611
rect 126 605 134 607
rect 142 607 150 609
rect 142 603 144 607
rect 148 603 150 607
rect 158 607 160 611
rect 164 607 166 611
rect 190 611 198 613
rect 206 611 214 613
rect 238 612 246 614
rect 254 611 262 613
rect 158 605 166 607
rect 174 608 182 610
rect 174 604 176 608
rect 180 604 182 608
rect 190 607 192 611
rect 196 607 198 611
rect 222 609 230 611
rect 190 605 198 607
rect 206 607 214 609
rect 78 601 86 603
rect 110 601 118 603
rect 126 601 134 603
rect 142 601 150 603
rect 158 601 166 603
rect 174 602 182 604
rect 206 603 208 607
rect 212 603 214 607
rect 222 605 224 609
rect 228 605 230 609
rect 222 603 230 605
rect 238 608 246 610
rect 238 604 240 608
rect 244 604 246 608
rect 254 607 256 611
rect 260 607 262 611
rect 254 605 262 607
rect 270 612 278 614
rect 286 613 294 615
rect 302 617 310 619
rect 302 613 304 617
rect 308 613 310 617
rect 386 617 388 621
rect 392 617 394 621
rect 386 615 394 617
rect 402 621 410 623
rect 402 617 404 621
rect 408 617 410 621
rect 402 615 410 617
rect 418 621 426 623
rect 418 617 420 621
rect 424 617 426 621
rect 418 615 426 617
rect 434 621 442 623
rect 434 617 436 621
rect 440 617 442 621
rect 434 615 442 617
rect 450 621 458 623
rect 450 617 452 621
rect 456 617 458 621
rect 450 615 458 617
rect 466 621 474 623
rect 466 617 468 621
rect 472 617 474 621
rect 466 615 474 617
rect 482 621 490 623
rect 482 617 484 621
rect 488 617 490 621
rect 482 615 490 617
rect 498 621 506 623
rect 498 617 500 621
rect 504 617 506 621
rect 498 615 506 617
rect 514 621 522 623
rect 514 617 516 621
rect 520 617 522 621
rect 514 615 522 617
rect 530 621 538 623
rect 530 617 532 621
rect 536 617 538 621
rect 530 615 538 617
rect 546 621 554 623
rect 546 617 548 621
rect 552 617 554 621
rect 546 615 554 617
rect 562 621 570 623
rect 562 617 564 621
rect 568 617 570 621
rect 562 615 570 617
rect 578 621 586 623
rect 578 617 580 621
rect 584 617 586 621
rect 578 615 586 617
rect 590 622 598 624
rect 590 618 592 622
rect 596 618 598 622
rect 590 616 598 618
rect 270 608 272 612
rect 276 608 278 612
rect 302 611 310 613
rect 386 611 394 613
rect 270 606 278 608
rect 286 609 294 611
rect 286 605 288 609
rect 292 605 294 609
rect 14 598 22 600
rect 44 599 52 601
rect 94 599 102 601
rect 28 597 36 599
rect 2 594 10 596
rect 14 594 22 596
rect 2 590 10 592
rect 2 586 4 590
rect 8 586 10 590
rect 14 590 16 594
rect 20 590 22 594
rect 28 593 30 597
rect 34 593 36 597
rect 44 595 46 599
rect 50 595 52 599
rect 44 593 52 595
rect 60 597 68 599
rect 60 593 62 597
rect 66 593 68 597
rect 28 591 36 593
rect 60 591 68 593
rect 78 597 86 599
rect 78 593 80 597
rect 84 593 86 597
rect 94 595 96 599
rect 100 595 102 599
rect 94 593 102 595
rect 110 597 118 599
rect 110 593 112 597
rect 116 593 118 597
rect 126 597 128 601
rect 132 597 134 601
rect 126 595 134 597
rect 142 597 150 599
rect 142 593 144 597
rect 148 593 150 597
rect 158 597 160 601
rect 164 597 166 601
rect 190 601 198 603
rect 206 601 214 603
rect 238 602 246 604
rect 254 601 262 603
rect 158 595 166 597
rect 174 598 182 600
rect 174 594 176 598
rect 180 594 182 598
rect 190 597 192 601
rect 196 597 198 601
rect 222 599 230 601
rect 190 595 198 597
rect 206 597 214 599
rect 78 591 86 593
rect 110 591 118 593
rect 126 591 134 593
rect 142 591 150 593
rect 158 591 166 593
rect 174 592 182 594
rect 206 593 208 597
rect 212 593 214 597
rect 222 595 224 599
rect 228 595 230 599
rect 222 593 230 595
rect 238 598 246 600
rect 238 594 240 598
rect 244 594 246 598
rect 254 597 256 601
rect 260 597 262 601
rect 254 595 262 597
rect 270 602 278 604
rect 286 603 294 605
rect 302 607 310 609
rect 302 603 304 607
rect 308 603 310 607
rect 386 607 388 611
rect 392 607 394 611
rect 386 605 394 607
rect 402 611 410 613
rect 402 607 404 611
rect 408 607 410 611
rect 402 605 410 607
rect 418 611 426 613
rect 418 607 420 611
rect 424 607 426 611
rect 418 605 426 607
rect 434 611 442 613
rect 434 607 436 611
rect 440 607 442 611
rect 434 605 442 607
rect 450 611 458 613
rect 450 607 452 611
rect 456 607 458 611
rect 450 605 458 607
rect 466 611 474 613
rect 466 607 468 611
rect 472 607 474 611
rect 466 605 474 607
rect 482 611 490 613
rect 482 607 484 611
rect 488 607 490 611
rect 482 605 490 607
rect 498 611 506 613
rect 498 607 500 611
rect 504 607 506 611
rect 498 605 506 607
rect 514 611 522 613
rect 514 607 516 611
rect 520 607 522 611
rect 514 605 522 607
rect 530 611 538 613
rect 530 607 532 611
rect 536 607 538 611
rect 530 605 538 607
rect 546 611 554 613
rect 546 607 548 611
rect 552 607 554 611
rect 546 605 554 607
rect 562 611 570 613
rect 562 607 564 611
rect 568 607 570 611
rect 562 605 570 607
rect 578 611 586 613
rect 578 607 580 611
rect 584 607 586 611
rect 578 605 586 607
rect 590 612 598 614
rect 590 608 592 612
rect 596 608 598 612
rect 590 606 598 608
rect 270 598 272 602
rect 276 598 278 602
rect 302 601 310 603
rect 386 601 394 603
rect 270 596 278 598
rect 286 599 294 601
rect 286 595 288 599
rect 292 595 294 599
rect 14 588 22 590
rect 44 589 52 591
rect 94 589 102 591
rect 28 587 36 589
rect 2 584 10 586
rect 14 584 22 586
rect 2 580 10 582
rect 2 576 4 580
rect 8 576 10 580
rect 14 580 16 584
rect 20 580 22 584
rect 28 583 30 587
rect 34 583 36 587
rect 44 585 46 589
rect 50 585 52 589
rect 44 583 52 585
rect 60 587 68 589
rect 60 583 62 587
rect 66 583 68 587
rect 28 581 36 583
rect 60 581 68 583
rect 78 587 86 589
rect 78 583 80 587
rect 84 583 86 587
rect 94 585 96 589
rect 100 585 102 589
rect 94 583 102 585
rect 110 587 118 589
rect 110 583 112 587
rect 116 583 118 587
rect 126 587 128 591
rect 132 587 134 591
rect 126 585 134 587
rect 142 587 150 589
rect 142 583 144 587
rect 148 583 150 587
rect 158 587 160 591
rect 164 587 166 591
rect 190 591 198 593
rect 206 591 214 593
rect 238 592 246 594
rect 254 591 262 593
rect 158 585 166 587
rect 174 588 182 590
rect 174 584 176 588
rect 180 584 182 588
rect 190 587 192 591
rect 196 587 198 591
rect 222 589 230 591
rect 190 585 198 587
rect 206 587 214 589
rect 78 581 86 583
rect 110 581 118 583
rect 126 581 134 583
rect 142 581 150 583
rect 158 581 166 583
rect 174 582 182 584
rect 206 583 208 587
rect 212 583 214 587
rect 222 585 224 589
rect 228 585 230 589
rect 222 583 230 585
rect 238 588 246 590
rect 238 584 240 588
rect 244 584 246 588
rect 254 587 256 591
rect 260 587 262 591
rect 254 585 262 587
rect 270 592 278 594
rect 286 593 294 595
rect 302 597 310 599
rect 302 593 304 597
rect 308 593 310 597
rect 386 597 388 601
rect 392 597 394 601
rect 386 595 394 597
rect 402 601 410 603
rect 402 597 404 601
rect 408 597 410 601
rect 402 595 410 597
rect 418 601 426 603
rect 418 597 420 601
rect 424 597 426 601
rect 418 595 426 597
rect 434 601 442 603
rect 434 597 436 601
rect 440 597 442 601
rect 434 595 442 597
rect 450 601 458 603
rect 450 597 452 601
rect 456 597 458 601
rect 450 595 458 597
rect 466 601 474 603
rect 466 597 468 601
rect 472 597 474 601
rect 466 595 474 597
rect 482 601 490 603
rect 482 597 484 601
rect 488 597 490 601
rect 482 595 490 597
rect 498 601 506 603
rect 498 597 500 601
rect 504 597 506 601
rect 498 595 506 597
rect 514 601 522 603
rect 514 597 516 601
rect 520 597 522 601
rect 514 595 522 597
rect 530 601 538 603
rect 530 597 532 601
rect 536 597 538 601
rect 530 595 538 597
rect 546 601 554 603
rect 546 597 548 601
rect 552 597 554 601
rect 546 595 554 597
rect 562 601 570 603
rect 562 597 564 601
rect 568 597 570 601
rect 562 595 570 597
rect 578 601 586 603
rect 578 597 580 601
rect 584 597 586 601
rect 578 595 586 597
rect 590 602 598 604
rect 590 598 592 602
rect 596 598 598 602
rect 590 596 598 598
rect 270 588 272 592
rect 276 588 278 592
rect 302 591 310 593
rect 386 591 394 593
rect 270 586 278 588
rect 286 589 294 591
rect 286 585 288 589
rect 292 585 294 589
rect 14 578 22 580
rect 44 579 52 581
rect 94 579 102 581
rect 28 577 36 579
rect 2 574 10 576
rect 14 574 22 576
rect 2 570 10 572
rect 2 566 4 570
rect 8 566 10 570
rect 14 570 16 574
rect 20 570 22 574
rect 28 573 30 577
rect 34 573 36 577
rect 44 575 46 579
rect 50 575 52 579
rect 44 573 52 575
rect 60 577 68 579
rect 60 573 62 577
rect 66 573 68 577
rect 28 571 36 573
rect 60 571 68 573
rect 78 577 86 579
rect 78 573 80 577
rect 84 573 86 577
rect 94 575 96 579
rect 100 575 102 579
rect 94 573 102 575
rect 110 577 118 579
rect 110 573 112 577
rect 116 573 118 577
rect 126 577 128 581
rect 132 577 134 581
rect 126 575 134 577
rect 142 577 150 579
rect 142 573 144 577
rect 148 573 150 577
rect 158 577 160 581
rect 164 577 166 581
rect 190 581 198 583
rect 206 581 214 583
rect 238 582 246 584
rect 254 581 262 583
rect 158 575 166 577
rect 174 578 182 580
rect 174 574 176 578
rect 180 574 182 578
rect 190 577 192 581
rect 196 577 198 581
rect 222 579 230 581
rect 190 575 198 577
rect 206 577 214 579
rect 78 571 86 573
rect 110 571 118 573
rect 126 571 134 573
rect 142 571 150 573
rect 158 571 166 573
rect 174 572 182 574
rect 206 573 208 577
rect 212 573 214 577
rect 222 575 224 579
rect 228 575 230 579
rect 222 573 230 575
rect 238 578 246 580
rect 238 574 240 578
rect 244 574 246 578
rect 254 577 256 581
rect 260 577 262 581
rect 254 575 262 577
rect 270 582 278 584
rect 286 583 294 585
rect 302 587 310 589
rect 302 583 304 587
rect 308 583 310 587
rect 386 587 388 591
rect 392 587 394 591
rect 386 585 394 587
rect 402 591 410 593
rect 402 587 404 591
rect 408 587 410 591
rect 402 585 410 587
rect 418 591 426 593
rect 418 587 420 591
rect 424 587 426 591
rect 418 585 426 587
rect 434 591 442 593
rect 434 587 436 591
rect 440 587 442 591
rect 434 585 442 587
rect 450 591 458 593
rect 450 587 452 591
rect 456 587 458 591
rect 450 585 458 587
rect 466 591 474 593
rect 466 587 468 591
rect 472 587 474 591
rect 466 585 474 587
rect 482 591 490 593
rect 482 587 484 591
rect 488 587 490 591
rect 482 585 490 587
rect 498 591 506 593
rect 498 587 500 591
rect 504 587 506 591
rect 498 585 506 587
rect 514 591 522 593
rect 514 587 516 591
rect 520 587 522 591
rect 514 585 522 587
rect 530 591 538 593
rect 530 587 532 591
rect 536 587 538 591
rect 530 585 538 587
rect 546 591 554 593
rect 546 587 548 591
rect 552 587 554 591
rect 546 585 554 587
rect 562 591 570 593
rect 562 587 564 591
rect 568 587 570 591
rect 562 585 570 587
rect 578 591 586 593
rect 578 587 580 591
rect 584 587 586 591
rect 578 585 586 587
rect 590 592 598 594
rect 590 588 592 592
rect 596 588 598 592
rect 590 586 598 588
rect 270 578 272 582
rect 276 578 278 582
rect 302 581 310 583
rect 386 581 394 583
rect 270 576 278 578
rect 286 579 294 581
rect 286 575 288 579
rect 292 575 294 579
rect 14 568 22 570
rect 44 569 52 571
rect 94 569 102 571
rect 28 567 36 569
rect 2 564 10 566
rect 14 564 22 566
rect 2 560 10 562
rect 2 556 4 560
rect 8 556 10 560
rect 14 560 16 564
rect 20 560 22 564
rect 28 563 30 567
rect 34 563 36 567
rect 44 565 46 569
rect 50 565 52 569
rect 44 563 52 565
rect 60 567 68 569
rect 60 563 62 567
rect 66 563 68 567
rect 28 561 36 563
rect 60 561 68 563
rect 78 567 86 569
rect 78 563 80 567
rect 84 563 86 567
rect 94 565 96 569
rect 100 565 102 569
rect 94 563 102 565
rect 110 567 118 569
rect 110 563 112 567
rect 116 563 118 567
rect 126 567 128 571
rect 132 567 134 571
rect 126 565 134 567
rect 142 567 150 569
rect 142 563 144 567
rect 148 563 150 567
rect 158 567 160 571
rect 164 567 166 571
rect 190 571 198 573
rect 206 571 214 573
rect 238 572 246 574
rect 254 571 262 573
rect 158 565 166 567
rect 174 568 182 570
rect 174 564 176 568
rect 180 564 182 568
rect 190 567 192 571
rect 196 567 198 571
rect 222 569 230 571
rect 190 565 198 567
rect 206 567 214 569
rect 78 561 86 563
rect 110 561 118 563
rect 126 561 134 563
rect 142 561 150 563
rect 158 561 166 563
rect 174 562 182 564
rect 206 563 208 567
rect 212 563 214 567
rect 222 565 224 569
rect 228 565 230 569
rect 222 563 230 565
rect 238 568 246 570
rect 238 564 240 568
rect 244 564 246 568
rect 254 567 256 571
rect 260 567 262 571
rect 254 565 262 567
rect 270 572 278 574
rect 286 573 294 575
rect 302 577 310 579
rect 302 573 304 577
rect 308 573 310 577
rect 386 577 388 581
rect 392 577 394 581
rect 386 575 394 577
rect 402 581 410 583
rect 402 577 404 581
rect 408 577 410 581
rect 402 575 410 577
rect 418 581 426 583
rect 418 577 420 581
rect 424 577 426 581
rect 418 575 426 577
rect 434 581 442 583
rect 434 577 436 581
rect 440 577 442 581
rect 434 575 442 577
rect 450 581 458 583
rect 450 577 452 581
rect 456 577 458 581
rect 450 575 458 577
rect 466 581 474 583
rect 466 577 468 581
rect 472 577 474 581
rect 466 575 474 577
rect 482 581 490 583
rect 482 577 484 581
rect 488 577 490 581
rect 482 575 490 577
rect 498 581 506 583
rect 498 577 500 581
rect 504 577 506 581
rect 498 575 506 577
rect 514 581 522 583
rect 514 577 516 581
rect 520 577 522 581
rect 514 575 522 577
rect 530 581 538 583
rect 530 577 532 581
rect 536 577 538 581
rect 530 575 538 577
rect 546 581 554 583
rect 546 577 548 581
rect 552 577 554 581
rect 546 575 554 577
rect 562 581 570 583
rect 562 577 564 581
rect 568 577 570 581
rect 562 575 570 577
rect 578 581 586 583
rect 578 577 580 581
rect 584 577 586 581
rect 578 575 586 577
rect 590 582 598 584
rect 590 578 592 582
rect 596 578 598 582
rect 590 576 598 578
rect 270 568 272 572
rect 276 568 278 572
rect 302 571 310 573
rect 386 571 394 573
rect 270 566 278 568
rect 286 569 294 571
rect 286 565 288 569
rect 292 565 294 569
rect 14 558 22 560
rect 44 559 52 561
rect 94 559 102 561
rect 28 557 36 559
rect 2 554 10 556
rect 14 554 22 556
rect 2 550 10 552
rect 2 546 4 550
rect 8 546 10 550
rect 14 550 16 554
rect 20 550 22 554
rect 28 553 30 557
rect 34 553 36 557
rect 44 555 46 559
rect 50 555 52 559
rect 44 553 52 555
rect 60 557 68 559
rect 60 553 62 557
rect 66 553 68 557
rect 28 551 36 553
rect 60 551 68 553
rect 78 557 86 559
rect 78 553 80 557
rect 84 553 86 557
rect 94 555 96 559
rect 100 555 102 559
rect 94 553 102 555
rect 110 557 118 559
rect 110 553 112 557
rect 116 553 118 557
rect 126 557 128 561
rect 132 557 134 561
rect 126 555 134 557
rect 142 557 150 559
rect 78 551 86 553
rect 110 551 118 553
rect 142 553 144 557
rect 148 553 150 557
rect 158 557 160 561
rect 164 557 166 561
rect 190 561 198 563
rect 206 561 214 563
rect 238 562 246 564
rect 254 561 262 563
rect 158 555 166 557
rect 174 558 182 560
rect 174 554 176 558
rect 180 554 182 558
rect 190 557 192 561
rect 196 557 198 561
rect 222 559 230 561
rect 190 555 198 557
rect 206 557 214 559
rect 142 551 150 553
rect 158 551 166 553
rect 174 552 182 554
rect 206 553 208 557
rect 212 553 214 557
rect 222 555 224 559
rect 228 555 230 559
rect 222 553 230 555
rect 238 558 246 560
rect 238 554 240 558
rect 244 554 246 558
rect 254 557 256 561
rect 260 557 262 561
rect 254 555 262 557
rect 270 562 278 564
rect 286 563 294 565
rect 302 567 310 569
rect 302 563 304 567
rect 308 563 310 567
rect 386 567 388 571
rect 392 567 394 571
rect 386 565 394 567
rect 402 571 410 573
rect 402 567 404 571
rect 408 567 410 571
rect 402 565 410 567
rect 418 571 426 573
rect 418 567 420 571
rect 424 567 426 571
rect 418 565 426 567
rect 434 571 442 573
rect 434 567 436 571
rect 440 567 442 571
rect 434 565 442 567
rect 450 571 458 573
rect 450 567 452 571
rect 456 567 458 571
rect 450 565 458 567
rect 466 571 474 573
rect 466 567 468 571
rect 472 567 474 571
rect 466 565 474 567
rect 482 571 490 573
rect 482 567 484 571
rect 488 567 490 571
rect 482 565 490 567
rect 498 571 506 573
rect 498 567 500 571
rect 504 567 506 571
rect 498 565 506 567
rect 514 571 522 573
rect 514 567 516 571
rect 520 567 522 571
rect 514 565 522 567
rect 530 571 538 573
rect 530 567 532 571
rect 536 567 538 571
rect 530 565 538 567
rect 546 571 554 573
rect 546 567 548 571
rect 552 567 554 571
rect 546 565 554 567
rect 562 571 570 573
rect 562 567 564 571
rect 568 567 570 571
rect 562 565 570 567
rect 578 571 586 573
rect 578 567 580 571
rect 584 567 586 571
rect 578 565 586 567
rect 590 572 598 574
rect 590 568 592 572
rect 596 568 598 572
rect 590 566 598 568
rect 270 558 272 562
rect 276 558 278 562
rect 302 561 310 563
rect 386 561 394 563
rect 270 556 278 558
rect 286 559 294 561
rect 286 555 288 559
rect 292 555 294 559
rect 14 548 22 550
rect 2 544 10 546
rect 28 547 36 549
rect 28 543 30 547
rect 34 543 36 547
rect 2 540 10 542
rect 28 541 36 543
rect 60 547 68 549
rect 60 543 62 547
rect 66 543 68 547
rect 60 541 68 543
rect 78 547 86 549
rect 78 543 80 547
rect 84 543 86 547
rect 78 541 86 543
rect 110 547 118 549
rect 110 543 112 547
rect 116 543 118 547
rect 110 541 118 543
rect 142 547 150 549
rect 142 543 144 547
rect 148 543 150 547
rect 158 547 160 551
rect 164 547 166 551
rect 190 551 198 553
rect 206 551 214 553
rect 238 552 246 554
rect 286 553 294 555
rect 302 557 310 559
rect 302 553 304 557
rect 308 553 310 557
rect 386 557 388 561
rect 392 557 394 561
rect 386 555 394 557
rect 402 561 410 563
rect 402 557 404 561
rect 408 557 410 561
rect 402 555 410 557
rect 418 561 426 563
rect 418 557 420 561
rect 424 557 426 561
rect 418 555 426 557
rect 434 561 442 563
rect 434 557 436 561
rect 440 557 442 561
rect 434 555 442 557
rect 450 561 458 563
rect 450 557 452 561
rect 456 557 458 561
rect 450 555 458 557
rect 466 561 474 563
rect 466 557 468 561
rect 472 557 474 561
rect 466 555 474 557
rect 482 561 490 563
rect 482 557 484 561
rect 488 557 490 561
rect 482 555 490 557
rect 498 561 506 563
rect 498 557 500 561
rect 504 557 506 561
rect 498 555 506 557
rect 514 561 522 563
rect 514 557 516 561
rect 520 557 522 561
rect 514 555 522 557
rect 530 561 538 563
rect 530 557 532 561
rect 536 557 538 561
rect 530 555 538 557
rect 546 561 554 563
rect 546 557 548 561
rect 552 557 554 561
rect 546 555 554 557
rect 562 561 570 563
rect 562 557 564 561
rect 568 557 570 561
rect 562 555 570 557
rect 578 561 586 563
rect 578 557 580 561
rect 584 557 586 561
rect 578 555 586 557
rect 590 562 598 564
rect 590 558 592 562
rect 596 558 598 562
rect 590 556 598 558
rect 254 551 262 553
rect 302 551 310 553
rect 386 551 394 553
rect 158 545 166 547
rect 174 548 182 550
rect 142 541 150 543
rect 174 544 176 548
rect 180 544 182 548
rect 190 547 192 551
rect 196 547 198 551
rect 190 545 198 547
rect 206 547 214 549
rect 174 542 182 544
rect 206 543 208 547
rect 212 543 214 547
rect 206 541 214 543
rect 238 548 246 550
rect 238 544 240 548
rect 244 544 246 548
rect 254 547 256 551
rect 260 547 262 551
rect 254 545 262 547
rect 286 549 294 551
rect 286 545 288 549
rect 292 545 294 549
rect 238 542 246 544
rect 286 543 294 545
rect 302 547 310 549
rect 302 543 304 547
rect 308 543 310 547
rect 386 547 388 551
rect 392 547 394 551
rect 386 545 394 547
rect 402 551 410 553
rect 402 547 404 551
rect 408 547 410 551
rect 402 545 410 547
rect 418 551 426 553
rect 418 547 420 551
rect 424 547 426 551
rect 418 545 426 547
rect 434 551 442 553
rect 434 547 436 551
rect 440 547 442 551
rect 434 545 442 547
rect 450 551 458 553
rect 450 547 452 551
rect 456 547 458 551
rect 450 545 458 547
rect 466 551 474 553
rect 466 547 468 551
rect 472 547 474 551
rect 466 545 474 547
rect 482 551 490 553
rect 482 547 484 551
rect 488 547 490 551
rect 482 545 490 547
rect 498 551 506 553
rect 498 547 500 551
rect 504 547 506 551
rect 498 545 506 547
rect 514 551 522 553
rect 514 547 516 551
rect 520 547 522 551
rect 514 545 522 547
rect 530 551 538 553
rect 530 547 532 551
rect 536 547 538 551
rect 530 545 538 547
rect 546 551 554 553
rect 546 547 548 551
rect 552 547 554 551
rect 546 545 554 547
rect 562 551 570 553
rect 562 547 564 551
rect 568 547 570 551
rect 562 545 570 547
rect 578 551 586 553
rect 578 547 580 551
rect 584 547 586 551
rect 578 545 586 547
rect 590 552 598 554
rect 590 548 592 552
rect 596 548 598 552
rect 590 546 598 548
rect 302 541 310 543
rect 590 542 598 544
rect 2 536 4 540
rect 8 536 10 540
rect 2 534 10 536
rect 580 539 588 541
rect 580 535 582 539
rect 586 535 588 539
rect 590 538 592 542
rect 596 538 598 542
rect 590 536 598 538
rect 22 533 30 535
rect 2 530 10 532
rect 2 526 4 530
rect 8 526 10 530
rect 22 529 24 533
rect 28 529 30 533
rect 22 527 30 529
rect 32 533 40 535
rect 32 529 34 533
rect 38 529 40 533
rect 32 527 40 529
rect 50 533 58 535
rect 50 529 52 533
rect 56 529 58 533
rect 50 527 58 529
rect 60 533 68 535
rect 60 529 62 533
rect 66 529 68 533
rect 60 527 68 529
rect 90 533 98 535
rect 90 529 92 533
rect 96 529 98 533
rect 90 527 98 529
rect 100 533 108 535
rect 580 533 588 535
rect 100 529 102 533
rect 106 529 108 533
rect 590 532 598 534
rect 580 529 588 531
rect 100 527 108 529
rect 386 527 394 529
rect 2 524 10 526
rect 118 524 126 526
rect 2 520 10 522
rect 2 516 4 520
rect 8 516 10 520
rect 118 520 120 524
rect 124 520 126 524
rect 118 518 126 520
rect 128 524 136 526
rect 128 520 130 524
rect 134 520 136 524
rect 128 518 136 520
rect 138 524 146 526
rect 138 520 140 524
rect 144 520 146 524
rect 138 518 146 520
rect 148 524 156 526
rect 148 520 150 524
rect 154 520 156 524
rect 148 518 156 520
rect 158 524 166 526
rect 158 520 160 524
rect 164 520 166 524
rect 158 518 166 520
rect 168 524 176 526
rect 168 520 170 524
rect 174 520 176 524
rect 168 518 176 520
rect 178 524 186 526
rect 178 520 180 524
rect 184 520 186 524
rect 178 518 186 520
rect 188 524 196 526
rect 188 520 190 524
rect 194 520 196 524
rect 188 518 196 520
rect 198 524 206 526
rect 198 520 200 524
rect 204 520 206 524
rect 198 518 206 520
rect 208 524 216 526
rect 208 520 210 524
rect 214 520 216 524
rect 208 518 216 520
rect 218 524 226 526
rect 218 520 220 524
rect 224 520 226 524
rect 386 523 388 527
rect 392 523 394 527
rect 386 521 394 523
rect 482 527 490 529
rect 482 523 484 527
rect 488 523 490 527
rect 580 525 582 529
rect 586 525 588 529
rect 590 528 592 532
rect 596 528 598 532
rect 590 526 598 528
rect 580 523 588 525
rect 482 521 490 523
rect 590 522 598 524
rect 218 518 226 520
rect 527 519 535 521
rect 480 517 488 519
rect 2 514 10 516
rect 34 514 42 516
rect 4 510 12 512
rect 4 506 6 510
rect 10 506 12 510
rect 34 510 36 514
rect 40 510 42 514
rect 34 508 42 510
rect 44 514 52 516
rect 44 510 46 514
rect 50 510 52 514
rect 44 508 52 510
rect 54 514 62 516
rect 54 510 56 514
rect 60 510 62 514
rect 54 508 62 510
rect 64 514 72 516
rect 218 514 226 516
rect 64 510 66 514
rect 70 510 72 514
rect 64 508 72 510
rect 108 512 116 514
rect 108 508 110 512
rect 114 508 116 512
rect 108 506 116 508
rect 118 512 126 514
rect 118 508 120 512
rect 124 508 126 512
rect 118 506 126 508
rect 128 512 136 514
rect 128 508 130 512
rect 134 508 136 512
rect 128 506 136 508
rect 138 512 146 514
rect 138 508 140 512
rect 144 508 146 512
rect 138 506 146 508
rect 148 512 156 514
rect 148 508 150 512
rect 154 508 156 512
rect 148 506 156 508
rect 158 512 166 514
rect 158 508 160 512
rect 164 508 166 512
rect 158 506 166 508
rect 168 512 176 514
rect 168 508 170 512
rect 174 508 176 512
rect 168 506 176 508
rect 178 512 186 514
rect 178 508 180 512
rect 184 508 186 512
rect 178 506 186 508
rect 188 512 196 514
rect 188 508 190 512
rect 194 508 196 512
rect 188 506 196 508
rect 198 512 206 514
rect 198 508 200 512
rect 204 508 206 512
rect 198 506 206 508
rect 208 512 216 514
rect 208 508 210 512
rect 214 508 216 512
rect 218 510 220 514
rect 224 510 226 514
rect 218 508 226 510
rect 389 514 397 516
rect 389 510 391 514
rect 395 510 397 514
rect 389 508 397 510
rect 399 514 407 516
rect 399 510 401 514
rect 405 510 407 514
rect 399 508 407 510
rect 409 514 417 516
rect 409 510 411 514
rect 415 510 417 514
rect 409 508 417 510
rect 419 514 427 516
rect 419 510 421 514
rect 425 510 427 514
rect 419 508 427 510
rect 429 514 437 516
rect 429 510 431 514
rect 435 510 437 514
rect 429 508 437 510
rect 439 514 447 516
rect 439 510 441 514
rect 445 510 447 514
rect 439 508 447 510
rect 449 514 457 516
rect 449 510 451 514
rect 455 510 457 514
rect 480 513 482 517
rect 486 513 488 517
rect 480 511 488 513
rect 490 517 498 519
rect 490 513 492 517
rect 496 513 498 517
rect 490 511 498 513
rect 500 517 508 519
rect 500 513 502 517
rect 506 513 508 517
rect 527 515 529 519
rect 533 515 535 519
rect 527 513 535 515
rect 540 519 548 521
rect 540 515 542 519
rect 546 515 548 519
rect 540 513 548 515
rect 550 519 558 521
rect 550 515 552 519
rect 556 515 558 519
rect 550 513 558 515
rect 560 519 568 521
rect 560 515 562 519
rect 566 515 568 519
rect 560 513 568 515
rect 570 519 578 521
rect 570 515 572 519
rect 576 515 578 519
rect 570 513 578 515
rect 580 519 588 521
rect 580 515 582 519
rect 586 515 588 519
rect 590 518 592 522
rect 596 518 598 522
rect 590 516 598 518
rect 580 513 588 515
rect 500 511 508 513
rect 449 508 457 510
rect 590 510 598 512
rect 208 506 216 508
rect 590 506 592 510
rect 596 506 598 510
rect 4 504 12 506
rect 590 504 598 506
rect 4 500 12 502
rect 4 496 6 500
rect 10 496 12 500
rect 4 494 12 496
rect 34 500 42 502
rect 34 496 36 500
rect 40 496 42 500
rect 34 494 42 496
rect 44 500 52 502
rect 44 496 46 500
rect 50 496 52 500
rect 44 494 52 496
rect 54 500 62 502
rect 54 496 56 500
rect 60 496 62 500
rect 54 494 62 496
rect 64 500 72 502
rect 64 496 66 500
rect 70 496 72 500
rect 64 494 72 496
rect 106 500 114 502
rect 106 496 108 500
rect 112 496 114 500
rect 106 494 114 496
rect 116 500 124 502
rect 116 496 118 500
rect 122 496 124 500
rect 116 494 124 496
rect 126 500 134 502
rect 126 496 128 500
rect 132 496 134 500
rect 126 494 134 496
rect 136 500 144 502
rect 136 496 138 500
rect 142 496 144 500
rect 136 494 144 496
rect 146 500 154 502
rect 146 496 148 500
rect 152 496 154 500
rect 146 494 154 496
rect 156 500 164 502
rect 156 496 158 500
rect 162 496 164 500
rect 156 494 164 496
rect 166 500 174 502
rect 166 496 168 500
rect 172 496 174 500
rect 166 494 174 496
rect 176 500 184 502
rect 176 496 178 500
rect 182 496 184 500
rect 176 494 184 496
rect 186 500 194 502
rect 186 496 188 500
rect 192 496 194 500
rect 186 494 194 496
rect 196 500 204 502
rect 196 496 198 500
rect 202 496 204 500
rect 196 494 204 496
rect 206 500 214 502
rect 206 496 208 500
rect 212 496 214 500
rect 206 494 214 496
rect 222 500 230 502
rect 222 496 224 500
rect 228 496 230 500
rect 222 494 230 496
rect 232 500 240 502
rect 232 496 234 500
rect 238 496 240 500
rect 232 494 240 496
rect 389 500 397 502
rect 389 496 391 500
rect 395 496 397 500
rect 389 494 397 496
rect 399 500 407 502
rect 399 496 401 500
rect 405 496 407 500
rect 399 494 407 496
rect 409 500 417 502
rect 409 496 411 500
rect 415 496 417 500
rect 409 494 417 496
rect 419 500 427 502
rect 419 496 421 500
rect 425 496 427 500
rect 419 494 427 496
rect 429 500 437 502
rect 429 496 431 500
rect 435 496 437 500
rect 429 494 437 496
rect 439 500 447 502
rect 439 496 441 500
rect 445 496 447 500
rect 439 494 447 496
rect 449 500 457 502
rect 449 496 451 500
rect 455 496 457 500
rect 449 494 457 496
rect 527 500 535 502
rect 527 496 529 500
rect 533 496 535 500
rect 527 494 535 496
rect 537 500 545 502
rect 537 496 539 500
rect 543 496 545 500
rect 537 494 545 496
rect 547 500 555 502
rect 547 496 549 500
rect 553 496 555 500
rect 547 494 555 496
rect 557 500 565 502
rect 557 496 559 500
rect 563 496 565 500
rect 557 494 565 496
rect 567 500 575 502
rect 567 496 569 500
rect 573 496 575 500
rect 567 494 575 496
rect 580 500 588 502
rect 580 496 582 500
rect 586 496 588 500
rect 580 494 588 496
rect 590 500 598 502
rect 590 496 592 500
rect 596 496 598 500
rect 590 494 598 496
rect 4 490 12 492
rect 4 486 6 490
rect 10 486 12 490
rect 580 490 588 492
rect 580 486 582 490
rect 586 486 588 490
rect 4 484 12 486
rect 106 484 114 486
rect 34 482 42 484
rect 4 480 12 482
rect 4 476 6 480
rect 10 476 12 480
rect 34 478 36 482
rect 40 478 42 482
rect 34 476 42 478
rect 44 482 52 484
rect 44 478 46 482
rect 50 478 52 482
rect 44 476 52 478
rect 54 482 62 484
rect 54 478 56 482
rect 60 478 62 482
rect 54 476 62 478
rect 64 482 72 484
rect 64 478 66 482
rect 70 478 72 482
rect 64 476 72 478
rect 78 482 86 484
rect 78 478 80 482
rect 84 478 86 482
rect 106 480 108 484
rect 112 480 114 484
rect 106 478 114 480
rect 116 484 124 486
rect 116 480 118 484
rect 122 480 124 484
rect 116 478 124 480
rect 126 484 134 486
rect 126 480 128 484
rect 132 480 134 484
rect 126 478 134 480
rect 136 484 144 486
rect 136 480 138 484
rect 142 480 144 484
rect 136 478 144 480
rect 146 484 154 486
rect 146 480 148 484
rect 152 480 154 484
rect 146 478 154 480
rect 156 484 164 486
rect 156 480 158 484
rect 162 480 164 484
rect 156 478 164 480
rect 166 484 174 486
rect 166 480 168 484
rect 172 480 174 484
rect 166 478 174 480
rect 176 484 184 486
rect 176 480 178 484
rect 182 480 184 484
rect 176 478 184 480
rect 186 484 194 486
rect 186 480 188 484
rect 192 480 194 484
rect 186 478 194 480
rect 196 484 204 486
rect 196 480 198 484
rect 202 480 204 484
rect 196 478 204 480
rect 206 484 214 486
rect 206 480 208 484
rect 212 480 214 484
rect 206 478 214 480
rect 216 484 224 486
rect 216 480 218 484
rect 222 480 224 484
rect 216 478 224 480
rect 226 484 234 486
rect 226 480 228 484
rect 232 480 234 484
rect 226 478 234 480
rect 364 484 372 486
rect 364 480 366 484
rect 370 480 372 484
rect 364 478 372 480
rect 374 484 382 486
rect 374 480 376 484
rect 380 480 382 484
rect 374 478 382 480
rect 384 484 392 486
rect 384 480 386 484
rect 390 480 392 484
rect 384 478 392 480
rect 394 484 402 486
rect 394 480 396 484
rect 400 480 402 484
rect 394 478 402 480
rect 404 484 412 486
rect 404 480 406 484
rect 410 480 412 484
rect 404 478 412 480
rect 414 484 422 486
rect 414 480 416 484
rect 420 480 422 484
rect 414 478 422 480
rect 424 484 432 486
rect 424 480 426 484
rect 430 480 432 484
rect 424 478 432 480
rect 434 484 442 486
rect 434 480 436 484
rect 440 480 442 484
rect 434 478 442 480
rect 444 484 452 486
rect 444 480 446 484
rect 450 480 452 484
rect 444 478 452 480
rect 454 484 462 486
rect 454 480 456 484
rect 460 480 462 484
rect 454 478 462 480
rect 464 484 472 486
rect 464 480 466 484
rect 470 480 472 484
rect 464 478 472 480
rect 474 484 482 486
rect 474 480 476 484
rect 480 480 482 484
rect 474 478 482 480
rect 484 484 492 486
rect 580 484 588 486
rect 590 490 598 492
rect 590 486 592 490
rect 596 486 598 490
rect 590 484 598 486
rect 484 480 486 484
rect 490 480 492 484
rect 484 478 492 480
rect 527 482 535 484
rect 527 478 529 482
rect 533 478 535 482
rect 78 476 86 478
rect 296 476 304 478
rect 527 476 535 478
rect 542 482 550 484
rect 542 478 544 482
rect 548 478 550 482
rect 542 476 550 478
rect 552 482 560 484
rect 552 478 554 482
rect 558 478 560 482
rect 552 476 560 478
rect 580 480 588 482
rect 580 476 582 480
rect 586 476 588 480
rect 4 474 12 476
rect 106 474 114 476
rect 34 472 42 474
rect 4 470 12 472
rect 4 466 6 470
rect 10 466 12 470
rect 34 468 36 472
rect 40 468 42 472
rect 34 466 42 468
rect 44 472 52 474
rect 44 468 46 472
rect 50 468 52 472
rect 44 466 52 468
rect 54 472 62 474
rect 54 468 56 472
rect 60 468 62 472
rect 54 466 62 468
rect 64 472 72 474
rect 64 468 66 472
rect 70 468 72 472
rect 64 466 72 468
rect 78 470 86 472
rect 78 466 80 470
rect 84 466 86 470
rect 106 470 108 474
rect 112 470 114 474
rect 106 468 114 470
rect 116 474 124 476
rect 116 470 118 474
rect 122 470 124 474
rect 116 468 124 470
rect 126 474 134 476
rect 126 470 128 474
rect 132 470 134 474
rect 126 468 134 470
rect 136 474 144 476
rect 136 470 138 474
rect 142 470 144 474
rect 136 468 144 470
rect 146 474 154 476
rect 146 470 148 474
rect 152 470 154 474
rect 146 468 154 470
rect 156 474 164 476
rect 156 470 158 474
rect 162 470 164 474
rect 156 468 164 470
rect 166 474 174 476
rect 166 470 168 474
rect 172 470 174 474
rect 166 468 174 470
rect 176 474 184 476
rect 176 470 178 474
rect 182 470 184 474
rect 176 468 184 470
rect 186 474 194 476
rect 186 470 188 474
rect 192 470 194 474
rect 186 468 194 470
rect 196 474 204 476
rect 196 470 198 474
rect 202 470 204 474
rect 196 468 204 470
rect 206 474 214 476
rect 206 470 208 474
rect 212 470 214 474
rect 206 468 214 470
rect 216 474 224 476
rect 216 470 218 474
rect 222 470 224 474
rect 216 468 224 470
rect 226 474 234 476
rect 226 470 228 474
rect 232 470 234 474
rect 296 472 298 476
rect 302 472 304 476
rect 296 470 304 472
rect 364 474 372 476
rect 364 470 366 474
rect 370 470 372 474
rect 226 468 234 470
rect 364 468 372 470
rect 374 474 382 476
rect 374 470 376 474
rect 380 470 382 474
rect 374 468 382 470
rect 384 474 392 476
rect 384 470 386 474
rect 390 470 392 474
rect 384 468 392 470
rect 394 474 402 476
rect 394 470 396 474
rect 400 470 402 474
rect 394 468 402 470
rect 404 474 412 476
rect 404 470 406 474
rect 410 470 412 474
rect 404 468 412 470
rect 414 474 422 476
rect 414 470 416 474
rect 420 470 422 474
rect 414 468 422 470
rect 424 474 432 476
rect 424 470 426 474
rect 430 470 432 474
rect 424 468 432 470
rect 434 474 442 476
rect 434 470 436 474
rect 440 470 442 474
rect 434 468 442 470
rect 444 474 452 476
rect 444 470 446 474
rect 450 470 452 474
rect 444 468 452 470
rect 454 474 462 476
rect 454 470 456 474
rect 460 470 462 474
rect 454 468 462 470
rect 464 474 472 476
rect 464 470 466 474
rect 470 470 472 474
rect 464 468 472 470
rect 474 474 482 476
rect 474 470 476 474
rect 480 470 482 474
rect 474 468 482 470
rect 484 474 492 476
rect 580 474 588 476
rect 590 480 598 482
rect 590 476 592 480
rect 596 476 598 480
rect 590 474 598 476
rect 484 470 486 474
rect 490 470 492 474
rect 542 472 550 474
rect 484 468 492 470
rect 527 470 535 472
rect 296 466 304 468
rect 527 466 529 470
rect 533 466 535 470
rect 542 468 544 472
rect 548 468 550 472
rect 542 466 550 468
rect 552 472 560 474
rect 552 468 554 472
rect 558 468 560 472
rect 552 466 560 468
rect 580 470 588 472
rect 580 466 582 470
rect 586 466 588 470
rect 4 464 12 466
rect 78 464 86 466
rect 108 464 116 466
rect 34 462 42 464
rect 4 460 12 462
rect 4 456 6 460
rect 10 456 12 460
rect 34 458 36 462
rect 40 458 42 462
rect 34 456 42 458
rect 44 462 52 464
rect 44 458 46 462
rect 50 458 52 462
rect 108 460 110 464
rect 114 460 116 464
rect 108 458 116 460
rect 118 464 126 466
rect 118 460 120 464
rect 124 460 126 464
rect 118 458 126 460
rect 128 464 136 466
rect 128 460 130 464
rect 134 460 136 464
rect 128 458 136 460
rect 138 464 146 466
rect 138 460 140 464
rect 144 460 146 464
rect 138 458 146 460
rect 148 464 156 466
rect 148 460 150 464
rect 154 460 156 464
rect 148 458 156 460
rect 158 464 166 466
rect 158 460 160 464
rect 164 460 166 464
rect 158 458 166 460
rect 168 464 176 466
rect 168 460 170 464
rect 174 460 176 464
rect 168 458 176 460
rect 178 464 186 466
rect 178 460 180 464
rect 184 460 186 464
rect 178 458 186 460
rect 188 464 196 466
rect 188 460 190 464
rect 194 460 196 464
rect 188 458 196 460
rect 198 464 206 466
rect 198 460 200 464
rect 204 460 206 464
rect 198 458 206 460
rect 208 464 216 466
rect 208 460 210 464
rect 214 460 216 464
rect 208 458 216 460
rect 218 464 226 466
rect 218 460 220 464
rect 224 460 226 464
rect 218 458 226 460
rect 228 464 236 466
rect 228 460 230 464
rect 234 460 236 464
rect 296 462 298 466
rect 302 462 304 466
rect 296 460 304 462
rect 364 464 372 466
rect 364 460 366 464
rect 370 460 372 464
rect 228 458 236 460
rect 364 458 372 460
rect 374 464 382 466
rect 374 460 376 464
rect 380 460 382 464
rect 374 458 382 460
rect 384 464 392 466
rect 384 460 386 464
rect 390 460 392 464
rect 384 458 392 460
rect 394 464 402 466
rect 394 460 396 464
rect 400 460 402 464
rect 394 458 402 460
rect 404 464 412 466
rect 404 460 406 464
rect 410 460 412 464
rect 404 458 412 460
rect 414 464 422 466
rect 414 460 416 464
rect 420 460 422 464
rect 414 458 422 460
rect 424 464 432 466
rect 424 460 426 464
rect 430 460 432 464
rect 424 458 432 460
rect 434 464 442 466
rect 434 460 436 464
rect 440 460 442 464
rect 434 458 442 460
rect 444 464 452 466
rect 444 460 446 464
rect 450 460 452 464
rect 444 458 452 460
rect 454 464 462 466
rect 454 460 456 464
rect 460 460 462 464
rect 454 458 462 460
rect 464 464 472 466
rect 464 460 466 464
rect 470 460 472 464
rect 464 458 472 460
rect 474 464 482 466
rect 474 460 476 464
rect 480 460 482 464
rect 474 458 482 460
rect 484 464 492 466
rect 527 464 535 466
rect 580 464 588 466
rect 590 470 598 472
rect 590 466 592 470
rect 596 466 598 470
rect 590 464 598 466
rect 484 460 486 464
rect 490 460 492 464
rect 484 458 492 460
rect 542 459 550 461
rect 44 456 52 458
rect 296 456 304 458
rect 4 454 12 456
rect 34 452 42 454
rect 4 450 12 452
rect 4 446 6 450
rect 10 446 12 450
rect 34 448 36 452
rect 40 448 42 452
rect 34 446 42 448
rect 44 452 52 454
rect 108 452 116 454
rect 44 448 46 452
rect 50 448 52 452
rect 44 446 52 448
rect 64 450 72 452
rect 64 446 66 450
rect 70 446 72 450
rect 108 448 110 452
rect 114 448 116 452
rect 108 446 116 448
rect 118 452 126 454
rect 118 448 120 452
rect 124 448 126 452
rect 118 446 126 448
rect 128 452 136 454
rect 128 448 130 452
rect 134 448 136 452
rect 128 446 136 448
rect 138 452 146 454
rect 138 448 140 452
rect 144 448 146 452
rect 138 446 146 448
rect 148 452 156 454
rect 148 448 150 452
rect 154 448 156 452
rect 148 446 156 448
rect 158 452 166 454
rect 158 448 160 452
rect 164 448 166 452
rect 158 446 166 448
rect 168 452 176 454
rect 168 448 170 452
rect 174 448 176 452
rect 168 446 176 448
rect 178 452 186 454
rect 178 448 180 452
rect 184 448 186 452
rect 178 446 186 448
rect 188 452 196 454
rect 188 448 190 452
rect 194 448 196 452
rect 188 446 196 448
rect 198 452 206 454
rect 198 448 200 452
rect 204 448 206 452
rect 198 446 206 448
rect 208 452 216 454
rect 208 448 210 452
rect 214 448 216 452
rect 208 446 216 448
rect 218 452 226 454
rect 218 448 220 452
rect 224 448 226 452
rect 218 446 226 448
rect 228 452 236 454
rect 228 448 230 452
rect 234 448 236 452
rect 296 452 298 456
rect 302 452 304 456
rect 542 455 544 459
rect 548 455 550 459
rect 296 450 304 452
rect 364 452 372 454
rect 364 448 366 452
rect 370 448 372 452
rect 228 446 236 448
rect 296 446 304 448
rect 364 446 372 448
rect 374 452 382 454
rect 374 448 376 452
rect 380 448 382 452
rect 374 446 382 448
rect 384 452 392 454
rect 384 448 386 452
rect 390 448 392 452
rect 384 446 392 448
rect 394 452 402 454
rect 394 448 396 452
rect 400 448 402 452
rect 394 446 402 448
rect 404 452 412 454
rect 404 448 406 452
rect 410 448 412 452
rect 404 446 412 448
rect 414 452 422 454
rect 414 448 416 452
rect 420 448 422 452
rect 414 446 422 448
rect 424 452 432 454
rect 424 448 426 452
rect 430 448 432 452
rect 424 446 432 448
rect 434 452 442 454
rect 434 448 436 452
rect 440 448 442 452
rect 434 446 442 448
rect 444 452 452 454
rect 444 448 446 452
rect 450 448 452 452
rect 444 446 452 448
rect 454 452 462 454
rect 454 448 456 452
rect 460 448 462 452
rect 454 446 462 448
rect 464 452 472 454
rect 464 448 466 452
rect 470 448 472 452
rect 464 446 472 448
rect 474 452 482 454
rect 474 448 476 452
rect 480 448 482 452
rect 474 446 482 448
rect 484 452 492 454
rect 542 453 550 455
rect 552 459 560 461
rect 580 460 588 462
rect 552 455 554 459
rect 558 455 560 459
rect 552 453 560 455
rect 564 457 572 459
rect 564 453 566 457
rect 570 453 572 457
rect 580 456 582 460
rect 586 456 588 460
rect 580 454 588 456
rect 590 460 598 462
rect 590 456 592 460
rect 596 456 598 460
rect 590 454 598 456
rect 484 448 486 452
rect 490 448 492 452
rect 564 451 572 453
rect 484 446 492 448
rect 542 449 550 451
rect 4 444 12 446
rect 64 444 72 446
rect 34 442 42 444
rect 4 440 12 442
rect 4 436 6 440
rect 10 436 12 440
rect 34 438 36 442
rect 40 438 42 442
rect 34 436 42 438
rect 44 442 52 444
rect 44 438 46 442
rect 50 438 52 442
rect 296 442 298 446
rect 302 442 304 446
rect 542 445 544 449
rect 548 445 550 449
rect 542 443 550 445
rect 552 449 560 451
rect 580 450 588 452
rect 552 445 554 449
rect 558 445 560 449
rect 552 443 560 445
rect 564 447 572 449
rect 564 443 566 447
rect 570 443 572 447
rect 580 446 582 450
rect 586 446 588 450
rect 580 444 588 446
rect 590 450 598 452
rect 590 446 592 450
rect 596 446 598 450
rect 590 444 598 446
rect 296 440 304 442
rect 564 441 572 443
rect 542 439 550 441
rect 44 436 52 438
rect 296 436 304 438
rect 4 434 12 436
rect 34 432 42 434
rect 4 430 12 432
rect 4 426 6 430
rect 10 426 12 430
rect 34 428 36 432
rect 40 428 42 432
rect 34 426 42 428
rect 44 432 52 434
rect 44 428 46 432
rect 50 428 52 432
rect 44 426 52 428
rect 64 432 72 434
rect 64 428 66 432
rect 70 428 72 432
rect 296 432 298 436
rect 302 432 304 436
rect 542 435 544 439
rect 548 435 550 439
rect 296 430 304 432
rect 528 432 536 434
rect 542 433 550 435
rect 552 439 560 441
rect 580 440 588 442
rect 552 435 554 439
rect 558 435 560 439
rect 552 433 560 435
rect 564 437 572 439
rect 564 433 566 437
rect 570 433 572 437
rect 580 436 582 440
rect 586 436 588 440
rect 580 434 588 436
rect 590 440 598 442
rect 590 436 592 440
rect 596 436 598 440
rect 590 434 598 436
rect 64 426 72 428
rect 108 427 116 429
rect 4 424 12 426
rect 34 422 42 424
rect 4 420 12 422
rect 4 416 6 420
rect 10 416 12 420
rect 34 418 36 422
rect 40 418 42 422
rect 34 416 42 418
rect 44 422 52 424
rect 44 418 46 422
rect 50 418 52 422
rect 44 416 52 418
rect 64 422 72 424
rect 64 418 66 422
rect 70 418 72 422
rect 108 423 110 427
rect 114 423 116 427
rect 108 421 116 423
rect 118 427 126 429
rect 118 423 120 427
rect 124 423 126 427
rect 118 421 126 423
rect 128 427 136 429
rect 128 423 130 427
rect 134 423 136 427
rect 128 421 136 423
rect 138 427 146 429
rect 138 423 140 427
rect 144 423 146 427
rect 138 421 146 423
rect 148 427 156 429
rect 148 423 150 427
rect 154 423 156 427
rect 148 421 156 423
rect 158 427 166 429
rect 158 423 160 427
rect 164 423 166 427
rect 158 421 166 423
rect 168 427 176 429
rect 168 423 170 427
rect 174 423 176 427
rect 168 421 176 423
rect 178 427 186 429
rect 178 423 180 427
rect 184 423 186 427
rect 178 421 186 423
rect 188 427 196 429
rect 188 423 190 427
rect 194 423 196 427
rect 188 421 196 423
rect 198 427 206 429
rect 198 423 200 427
rect 204 423 206 427
rect 198 421 206 423
rect 208 427 216 429
rect 208 423 210 427
rect 214 423 216 427
rect 208 421 216 423
rect 218 427 226 429
rect 218 423 220 427
rect 224 423 226 427
rect 218 421 226 423
rect 228 427 236 429
rect 228 423 230 427
rect 234 423 236 427
rect 228 421 236 423
rect 296 426 304 428
rect 296 422 298 426
rect 302 422 304 426
rect 296 420 304 422
rect 364 427 372 429
rect 364 423 366 427
rect 370 423 372 427
rect 364 421 372 423
rect 374 427 382 429
rect 374 423 376 427
rect 380 423 382 427
rect 374 421 382 423
rect 384 427 392 429
rect 384 423 386 427
rect 390 423 392 427
rect 384 421 392 423
rect 394 427 402 429
rect 394 423 396 427
rect 400 423 402 427
rect 394 421 402 423
rect 404 427 412 429
rect 404 423 406 427
rect 410 423 412 427
rect 404 421 412 423
rect 414 427 422 429
rect 414 423 416 427
rect 420 423 422 427
rect 414 421 422 423
rect 424 427 432 429
rect 424 423 426 427
rect 430 423 432 427
rect 424 421 432 423
rect 434 427 442 429
rect 434 423 436 427
rect 440 423 442 427
rect 434 421 442 423
rect 444 427 452 429
rect 444 423 446 427
rect 450 423 452 427
rect 444 421 452 423
rect 454 427 462 429
rect 454 423 456 427
rect 460 423 462 427
rect 454 421 462 423
rect 464 427 472 429
rect 464 423 466 427
rect 470 423 472 427
rect 464 421 472 423
rect 474 427 482 429
rect 474 423 476 427
rect 480 423 482 427
rect 474 421 482 423
rect 484 427 492 429
rect 484 423 486 427
rect 490 423 492 427
rect 528 428 530 432
rect 534 428 536 432
rect 564 431 572 433
rect 528 426 536 428
rect 542 429 550 431
rect 542 425 544 429
rect 548 425 550 429
rect 484 421 492 423
rect 528 422 536 424
rect 542 423 550 425
rect 552 429 560 431
rect 580 430 588 432
rect 552 425 554 429
rect 558 425 560 429
rect 552 423 560 425
rect 564 427 572 429
rect 564 423 566 427
rect 570 423 572 427
rect 580 426 582 430
rect 586 426 588 430
rect 580 424 588 426
rect 590 430 598 432
rect 590 426 592 430
rect 596 426 598 430
rect 590 424 598 426
rect 528 418 530 422
rect 534 418 536 422
rect 564 421 572 423
rect 64 416 72 418
rect 296 416 304 418
rect 528 416 536 418
rect 542 419 550 421
rect 4 414 12 416
rect 34 412 42 414
rect 4 410 12 412
rect 4 406 6 410
rect 10 406 12 410
rect 34 408 36 412
rect 40 408 42 412
rect 34 406 42 408
rect 44 412 52 414
rect 44 408 46 412
rect 50 408 52 412
rect 44 406 52 408
rect 64 412 72 414
rect 64 408 66 412
rect 70 408 72 412
rect 296 412 298 416
rect 302 412 304 416
rect 542 415 544 419
rect 548 415 550 419
rect 296 410 304 412
rect 528 412 536 414
rect 542 413 550 415
rect 552 419 560 421
rect 580 420 588 422
rect 552 415 554 419
rect 558 415 560 419
rect 552 413 560 415
rect 564 417 572 419
rect 564 413 566 417
rect 570 413 572 417
rect 580 416 582 420
rect 586 416 588 420
rect 580 414 588 416
rect 590 420 598 422
rect 590 416 592 420
rect 596 416 598 420
rect 590 414 598 416
rect 528 408 530 412
rect 534 408 536 412
rect 564 411 572 413
rect 64 406 72 408
rect 296 406 304 408
rect 528 406 536 408
rect 542 409 550 411
rect 4 404 12 406
rect 34 402 42 404
rect 4 400 12 402
rect 4 396 6 400
rect 10 396 12 400
rect 34 398 36 402
rect 40 398 42 402
rect 34 396 42 398
rect 44 402 52 404
rect 44 398 46 402
rect 50 398 52 402
rect 44 396 52 398
rect 64 402 72 404
rect 64 398 66 402
rect 70 398 72 402
rect 296 402 298 406
rect 302 402 304 406
rect 542 405 544 409
rect 548 405 550 409
rect 296 400 304 402
rect 528 402 536 404
rect 542 403 550 405
rect 552 409 560 411
rect 580 410 588 412
rect 552 405 554 409
rect 558 405 560 409
rect 552 403 560 405
rect 564 407 572 409
rect 564 403 566 407
rect 570 403 572 407
rect 580 406 582 410
rect 586 406 588 410
rect 580 404 588 406
rect 590 410 598 412
rect 590 406 592 410
rect 596 406 598 410
rect 590 404 598 406
rect 64 396 72 398
rect 112 398 120 400
rect 4 394 12 396
rect 112 394 114 398
rect 118 394 120 398
rect 34 392 42 394
rect 4 390 12 392
rect 4 386 6 390
rect 10 386 12 390
rect 34 388 36 392
rect 40 388 42 392
rect 34 386 42 388
rect 44 392 52 394
rect 44 388 46 392
rect 50 388 52 392
rect 44 386 52 388
rect 64 392 72 394
rect 112 392 120 394
rect 122 398 130 400
rect 122 394 124 398
rect 128 394 130 398
rect 122 392 130 394
rect 132 398 140 400
rect 132 394 134 398
rect 138 394 140 398
rect 132 392 140 394
rect 142 398 150 400
rect 142 394 144 398
rect 148 394 150 398
rect 142 392 150 394
rect 152 398 160 400
rect 152 394 154 398
rect 158 394 160 398
rect 152 392 160 394
rect 162 398 170 400
rect 162 394 164 398
rect 168 394 170 398
rect 162 392 170 394
rect 172 398 180 400
rect 172 394 174 398
rect 178 394 180 398
rect 172 392 180 394
rect 182 398 190 400
rect 182 394 184 398
rect 188 394 190 398
rect 182 392 190 394
rect 192 398 200 400
rect 192 394 194 398
rect 198 394 200 398
rect 192 392 200 394
rect 202 398 210 400
rect 202 394 204 398
rect 208 394 210 398
rect 202 392 210 394
rect 212 398 220 400
rect 212 394 214 398
rect 218 394 220 398
rect 212 392 220 394
rect 222 398 230 400
rect 222 394 224 398
rect 228 394 230 398
rect 222 392 230 394
rect 232 398 240 400
rect 360 398 368 400
rect 232 394 234 398
rect 238 394 240 398
rect 232 392 240 394
rect 296 396 304 398
rect 296 392 298 396
rect 302 392 304 396
rect 360 394 362 398
rect 366 394 368 398
rect 360 392 368 394
rect 370 398 378 400
rect 370 394 372 398
rect 376 394 378 398
rect 370 392 378 394
rect 380 398 388 400
rect 380 394 382 398
rect 386 394 388 398
rect 380 392 388 394
rect 390 398 398 400
rect 390 394 392 398
rect 396 394 398 398
rect 390 392 398 394
rect 400 398 408 400
rect 400 394 402 398
rect 406 394 408 398
rect 400 392 408 394
rect 410 398 418 400
rect 410 394 412 398
rect 416 394 418 398
rect 410 392 418 394
rect 420 398 428 400
rect 420 394 422 398
rect 426 394 428 398
rect 420 392 428 394
rect 430 398 438 400
rect 430 394 432 398
rect 436 394 438 398
rect 430 392 438 394
rect 440 398 448 400
rect 440 394 442 398
rect 446 394 448 398
rect 440 392 448 394
rect 450 398 458 400
rect 450 394 452 398
rect 456 394 458 398
rect 450 392 458 394
rect 460 398 468 400
rect 460 394 462 398
rect 466 394 468 398
rect 460 392 468 394
rect 470 398 478 400
rect 470 394 472 398
rect 476 394 478 398
rect 470 392 478 394
rect 480 398 488 400
rect 480 394 482 398
rect 486 394 488 398
rect 528 398 530 402
rect 534 398 536 402
rect 564 401 572 403
rect 528 396 536 398
rect 542 399 550 401
rect 542 395 544 399
rect 548 395 550 399
rect 480 392 488 394
rect 528 392 536 394
rect 542 393 550 395
rect 552 399 560 401
rect 580 400 588 402
rect 552 395 554 399
rect 558 395 560 399
rect 552 393 560 395
rect 564 397 572 399
rect 564 393 566 397
rect 570 393 572 397
rect 580 396 582 400
rect 586 396 588 400
rect 580 394 588 396
rect 590 400 598 402
rect 590 396 592 400
rect 596 396 598 400
rect 590 394 598 396
rect 64 388 66 392
rect 70 388 72 392
rect 296 390 304 392
rect 528 388 530 392
rect 534 388 536 392
rect 564 391 572 393
rect 64 386 72 388
rect 112 386 120 388
rect 4 384 12 386
rect 34 382 42 384
rect 4 380 12 382
rect 4 376 6 380
rect 10 376 12 380
rect 34 378 36 382
rect 40 378 42 382
rect 34 376 42 378
rect 44 382 52 384
rect 44 378 46 382
rect 50 378 52 382
rect 44 376 52 378
rect 64 382 72 384
rect 64 378 66 382
rect 70 378 72 382
rect 112 382 114 386
rect 118 382 120 386
rect 112 380 120 382
rect 122 386 130 388
rect 122 382 124 386
rect 128 382 130 386
rect 122 380 130 382
rect 132 386 140 388
rect 132 382 134 386
rect 138 382 140 386
rect 132 380 140 382
rect 142 386 150 388
rect 142 382 144 386
rect 148 382 150 386
rect 142 380 150 382
rect 152 386 160 388
rect 152 382 154 386
rect 158 382 160 386
rect 152 380 160 382
rect 162 386 170 388
rect 162 382 164 386
rect 168 382 170 386
rect 162 380 170 382
rect 172 386 180 388
rect 172 382 174 386
rect 178 382 180 386
rect 172 380 180 382
rect 182 386 190 388
rect 182 382 184 386
rect 188 382 190 386
rect 182 380 190 382
rect 192 386 200 388
rect 192 382 194 386
rect 198 382 200 386
rect 192 380 200 382
rect 202 386 210 388
rect 202 382 204 386
rect 208 382 210 386
rect 202 380 210 382
rect 212 386 220 388
rect 212 382 214 386
rect 218 382 220 386
rect 212 380 220 382
rect 222 386 230 388
rect 222 382 224 386
rect 228 382 230 386
rect 222 380 230 382
rect 232 386 240 388
rect 232 382 234 386
rect 238 382 240 386
rect 232 380 240 382
rect 296 386 304 388
rect 296 382 298 386
rect 302 382 304 386
rect 296 380 304 382
rect 360 386 368 388
rect 360 382 362 386
rect 366 382 368 386
rect 360 380 368 382
rect 370 386 378 388
rect 370 382 372 386
rect 376 382 378 386
rect 370 380 378 382
rect 380 386 388 388
rect 380 382 382 386
rect 386 382 388 386
rect 380 380 388 382
rect 390 386 398 388
rect 390 382 392 386
rect 396 382 398 386
rect 390 380 398 382
rect 400 386 408 388
rect 400 382 402 386
rect 406 382 408 386
rect 400 380 408 382
rect 410 386 418 388
rect 410 382 412 386
rect 416 382 418 386
rect 410 380 418 382
rect 420 386 428 388
rect 420 382 422 386
rect 426 382 428 386
rect 420 380 428 382
rect 430 386 438 388
rect 430 382 432 386
rect 436 382 438 386
rect 430 380 438 382
rect 440 386 448 388
rect 440 382 442 386
rect 446 382 448 386
rect 440 380 448 382
rect 450 386 458 388
rect 450 382 452 386
rect 456 382 458 386
rect 450 380 458 382
rect 460 386 468 388
rect 460 382 462 386
rect 466 382 468 386
rect 460 380 468 382
rect 470 386 478 388
rect 470 382 472 386
rect 476 382 478 386
rect 470 380 478 382
rect 480 386 488 388
rect 528 386 536 388
rect 542 389 550 391
rect 480 382 482 386
rect 486 382 488 386
rect 542 385 544 389
rect 548 385 550 389
rect 480 380 488 382
rect 528 382 536 384
rect 542 383 550 385
rect 552 389 560 391
rect 580 390 588 392
rect 552 385 554 389
rect 558 385 560 389
rect 552 383 560 385
rect 564 387 572 389
rect 564 383 566 387
rect 570 383 572 387
rect 580 386 582 390
rect 586 386 588 390
rect 580 384 588 386
rect 590 390 598 392
rect 590 386 592 390
rect 596 386 598 390
rect 590 384 598 386
rect 528 378 530 382
rect 534 378 536 382
rect 564 381 572 383
rect 64 376 72 378
rect 296 376 304 378
rect 528 376 536 378
rect 542 379 550 381
rect 4 374 12 376
rect 34 372 42 374
rect 4 370 12 372
rect 4 366 6 370
rect 10 366 12 370
rect 34 368 36 372
rect 40 368 42 372
rect 34 366 42 368
rect 44 372 52 374
rect 44 368 46 372
rect 50 368 52 372
rect 44 366 52 368
rect 64 372 72 374
rect 64 368 66 372
rect 70 368 72 372
rect 296 372 298 376
rect 302 372 304 376
rect 542 375 544 379
rect 548 375 550 379
rect 296 370 304 372
rect 528 372 536 374
rect 542 373 550 375
rect 552 379 560 381
rect 580 380 588 382
rect 552 375 554 379
rect 558 375 560 379
rect 552 373 560 375
rect 564 377 572 379
rect 564 373 566 377
rect 570 373 572 377
rect 580 376 582 380
rect 586 376 588 380
rect 580 374 588 376
rect 590 380 598 382
rect 590 376 592 380
rect 596 376 598 380
rect 590 374 598 376
rect 528 368 530 372
rect 534 368 536 372
rect 564 371 572 373
rect 64 366 72 368
rect 296 366 304 368
rect 528 366 536 368
rect 542 369 550 371
rect 4 364 12 366
rect 34 362 42 364
rect 4 360 12 362
rect 4 356 6 360
rect 10 356 12 360
rect 34 358 36 362
rect 40 358 42 362
rect 34 356 42 358
rect 44 362 52 364
rect 44 358 46 362
rect 50 358 52 362
rect 44 356 52 358
rect 64 362 72 364
rect 296 362 298 366
rect 302 362 304 366
rect 542 365 544 369
rect 548 365 550 369
rect 528 362 536 364
rect 542 363 550 365
rect 552 369 560 371
rect 580 370 588 372
rect 552 365 554 369
rect 558 365 560 369
rect 552 363 560 365
rect 564 367 572 369
rect 564 363 566 367
rect 570 363 572 367
rect 580 366 582 370
rect 586 366 588 370
rect 580 364 588 366
rect 590 370 598 372
rect 590 366 592 370
rect 596 366 598 370
rect 590 364 598 366
rect 64 358 66 362
rect 70 358 72 362
rect 64 356 72 358
rect 112 360 120 362
rect 112 356 114 360
rect 118 356 120 360
rect 4 354 12 356
rect 112 354 120 356
rect 122 360 130 362
rect 122 356 124 360
rect 128 356 130 360
rect 122 354 130 356
rect 132 360 140 362
rect 132 356 134 360
rect 138 356 140 360
rect 132 354 140 356
rect 142 360 150 362
rect 142 356 144 360
rect 148 356 150 360
rect 142 354 150 356
rect 152 360 160 362
rect 152 356 154 360
rect 158 356 160 360
rect 152 354 160 356
rect 162 360 170 362
rect 162 356 164 360
rect 168 356 170 360
rect 162 354 170 356
rect 172 360 180 362
rect 172 356 174 360
rect 178 356 180 360
rect 172 354 180 356
rect 182 360 190 362
rect 182 356 184 360
rect 188 356 190 360
rect 182 354 190 356
rect 192 360 200 362
rect 192 356 194 360
rect 198 356 200 360
rect 192 354 200 356
rect 202 360 210 362
rect 202 356 204 360
rect 208 356 210 360
rect 202 354 210 356
rect 212 360 220 362
rect 212 356 214 360
rect 218 356 220 360
rect 212 354 220 356
rect 222 360 230 362
rect 222 356 224 360
rect 228 356 230 360
rect 222 354 230 356
rect 232 360 240 362
rect 296 360 304 362
rect 364 360 372 362
rect 232 356 234 360
rect 238 356 240 360
rect 232 354 240 356
rect 296 356 304 358
rect 34 352 42 354
rect 4 350 12 352
rect 4 346 6 350
rect 10 346 12 350
rect 34 348 36 352
rect 40 348 42 352
rect 34 346 42 348
rect 44 352 52 354
rect 44 348 46 352
rect 50 348 52 352
rect 44 346 52 348
rect 64 352 72 354
rect 64 348 66 352
rect 70 348 72 352
rect 296 352 298 356
rect 302 352 304 356
rect 364 356 366 360
rect 370 356 372 360
rect 364 354 372 356
rect 374 360 382 362
rect 374 356 376 360
rect 380 356 382 360
rect 374 354 382 356
rect 384 360 392 362
rect 384 356 386 360
rect 390 356 392 360
rect 384 354 392 356
rect 394 360 402 362
rect 394 356 396 360
rect 400 356 402 360
rect 394 354 402 356
rect 404 360 412 362
rect 404 356 406 360
rect 410 356 412 360
rect 404 354 412 356
rect 414 360 422 362
rect 414 356 416 360
rect 420 356 422 360
rect 414 354 422 356
rect 424 360 432 362
rect 424 356 426 360
rect 430 356 432 360
rect 424 354 432 356
rect 434 360 442 362
rect 434 356 436 360
rect 440 356 442 360
rect 434 354 442 356
rect 444 360 452 362
rect 444 356 446 360
rect 450 356 452 360
rect 444 354 452 356
rect 454 360 462 362
rect 454 356 456 360
rect 460 356 462 360
rect 454 354 462 356
rect 464 360 472 362
rect 464 356 466 360
rect 470 356 472 360
rect 464 354 472 356
rect 474 360 482 362
rect 474 356 476 360
rect 480 356 482 360
rect 474 354 482 356
rect 484 360 492 362
rect 484 356 486 360
rect 490 356 492 360
rect 528 358 530 362
rect 534 358 536 362
rect 564 361 572 363
rect 528 356 536 358
rect 542 359 550 361
rect 484 354 492 356
rect 542 355 544 359
rect 548 355 550 359
rect 296 350 304 352
rect 528 352 536 354
rect 542 353 550 355
rect 552 359 560 361
rect 580 360 588 362
rect 552 355 554 359
rect 558 355 560 359
rect 552 353 560 355
rect 564 357 572 359
rect 564 353 566 357
rect 570 353 572 357
rect 580 356 582 360
rect 586 356 588 360
rect 580 354 588 356
rect 590 360 598 362
rect 590 356 592 360
rect 596 356 598 360
rect 590 354 598 356
rect 528 348 530 352
rect 534 348 536 352
rect 564 351 572 353
rect 64 346 72 348
rect 296 346 304 348
rect 528 346 536 348
rect 542 349 550 351
rect 4 344 12 346
rect 34 342 42 344
rect 4 340 12 342
rect 4 336 6 340
rect 10 336 12 340
rect 34 338 36 342
rect 40 338 42 342
rect 34 336 42 338
rect 44 342 52 344
rect 44 338 46 342
rect 50 338 52 342
rect 44 336 52 338
rect 64 342 72 344
rect 64 338 66 342
rect 70 338 72 342
rect 296 342 298 346
rect 302 342 304 346
rect 542 345 544 349
rect 548 345 550 349
rect 296 340 304 342
rect 528 342 536 344
rect 542 343 550 345
rect 552 349 560 351
rect 580 350 588 352
rect 552 345 554 349
rect 558 345 560 349
rect 552 343 560 345
rect 564 347 572 349
rect 564 343 566 347
rect 570 343 572 347
rect 580 346 582 350
rect 586 346 588 350
rect 580 344 588 346
rect 590 350 598 352
rect 590 346 592 350
rect 596 346 598 350
rect 590 344 598 346
rect 528 338 530 342
rect 534 338 536 342
rect 564 341 572 343
rect 64 336 72 338
rect 296 336 304 338
rect 528 336 536 338
rect 542 339 550 341
rect 4 334 12 336
rect 34 332 42 334
rect 4 330 12 332
rect 4 326 6 330
rect 10 326 12 330
rect 34 328 36 332
rect 40 328 42 332
rect 34 326 42 328
rect 44 332 52 334
rect 44 328 46 332
rect 50 328 52 332
rect 44 326 52 328
rect 64 332 72 334
rect 64 328 66 332
rect 70 328 72 332
rect 64 326 72 328
rect 110 332 118 334
rect 110 328 112 332
rect 116 328 118 332
rect 110 326 118 328
rect 120 332 128 334
rect 120 328 122 332
rect 126 328 128 332
rect 120 326 128 328
rect 130 332 138 334
rect 130 328 132 332
rect 136 328 138 332
rect 130 326 138 328
rect 140 332 148 334
rect 140 328 142 332
rect 146 328 148 332
rect 140 326 148 328
rect 150 332 158 334
rect 150 328 152 332
rect 156 328 158 332
rect 150 326 158 328
rect 160 332 168 334
rect 160 328 162 332
rect 166 328 168 332
rect 160 326 168 328
rect 170 332 178 334
rect 170 328 172 332
rect 176 328 178 332
rect 170 326 178 328
rect 180 332 188 334
rect 180 328 182 332
rect 186 328 188 332
rect 180 326 188 328
rect 190 332 198 334
rect 190 328 192 332
rect 196 328 198 332
rect 190 326 198 328
rect 200 332 208 334
rect 200 328 202 332
rect 206 328 208 332
rect 200 326 208 328
rect 210 332 218 334
rect 210 328 212 332
rect 216 328 218 332
rect 210 326 218 328
rect 220 332 228 334
rect 220 328 222 332
rect 226 328 228 332
rect 220 326 228 328
rect 230 332 238 334
rect 230 328 232 332
rect 236 328 238 332
rect 296 332 298 336
rect 302 332 304 336
rect 542 335 544 339
rect 548 335 550 339
rect 296 330 304 332
rect 363 333 371 335
rect 363 329 365 333
rect 369 329 371 333
rect 230 326 238 328
rect 296 326 304 328
rect 363 327 371 329
rect 373 333 381 335
rect 373 329 375 333
rect 379 329 381 333
rect 373 327 381 329
rect 383 333 391 335
rect 383 329 385 333
rect 389 329 391 333
rect 383 327 391 329
rect 393 333 401 335
rect 393 329 395 333
rect 399 329 401 333
rect 393 327 401 329
rect 403 333 411 335
rect 403 329 405 333
rect 409 329 411 333
rect 403 327 411 329
rect 413 333 421 335
rect 413 329 415 333
rect 419 329 421 333
rect 413 327 421 329
rect 423 333 431 335
rect 423 329 425 333
rect 429 329 431 333
rect 423 327 431 329
rect 433 333 441 335
rect 433 329 435 333
rect 439 329 441 333
rect 433 327 441 329
rect 443 333 451 335
rect 443 329 445 333
rect 449 329 451 333
rect 443 327 451 329
rect 453 333 461 335
rect 453 329 455 333
rect 459 329 461 333
rect 453 327 461 329
rect 463 333 471 335
rect 463 329 465 333
rect 469 329 471 333
rect 463 327 471 329
rect 473 333 481 335
rect 473 329 475 333
rect 479 329 481 333
rect 473 327 481 329
rect 483 333 491 335
rect 483 329 485 333
rect 489 329 491 333
rect 483 327 491 329
rect 528 332 536 334
rect 542 333 550 335
rect 552 339 560 341
rect 580 340 588 342
rect 552 335 554 339
rect 558 335 560 339
rect 552 333 560 335
rect 564 337 572 339
rect 564 333 566 337
rect 570 333 572 337
rect 580 336 582 340
rect 586 336 588 340
rect 580 334 588 336
rect 590 340 598 342
rect 590 336 592 340
rect 596 336 598 340
rect 590 334 598 336
rect 528 328 530 332
rect 534 328 536 332
rect 564 331 572 333
rect 528 326 536 328
rect 542 329 550 331
rect 4 324 12 326
rect 34 322 42 324
rect 4 320 12 322
rect 4 316 6 320
rect 10 316 12 320
rect 34 318 36 322
rect 40 318 42 322
rect 34 316 42 318
rect 44 322 52 324
rect 44 318 46 322
rect 50 318 52 322
rect 44 316 52 318
rect 64 322 72 324
rect 296 322 298 326
rect 302 322 304 326
rect 542 325 544 329
rect 548 325 550 329
rect 64 318 66 322
rect 70 318 72 322
rect 64 316 72 318
rect 110 320 118 322
rect 110 316 112 320
rect 116 316 118 320
rect 4 314 12 316
rect 110 314 118 316
rect 120 320 128 322
rect 120 316 122 320
rect 126 316 128 320
rect 120 314 128 316
rect 130 320 138 322
rect 130 316 132 320
rect 136 316 138 320
rect 130 314 138 316
rect 140 320 148 322
rect 140 316 142 320
rect 146 316 148 320
rect 140 314 148 316
rect 150 320 158 322
rect 150 316 152 320
rect 156 316 158 320
rect 150 314 158 316
rect 160 320 168 322
rect 160 316 162 320
rect 166 316 168 320
rect 160 314 168 316
rect 170 320 178 322
rect 170 316 172 320
rect 176 316 178 320
rect 170 314 178 316
rect 180 320 188 322
rect 180 316 182 320
rect 186 316 188 320
rect 180 314 188 316
rect 190 320 198 322
rect 190 316 192 320
rect 196 316 198 320
rect 190 314 198 316
rect 200 320 208 322
rect 200 316 202 320
rect 206 316 208 320
rect 200 314 208 316
rect 210 320 218 322
rect 210 316 212 320
rect 216 316 218 320
rect 210 314 218 316
rect 220 320 228 322
rect 220 316 222 320
rect 226 316 228 320
rect 220 314 228 316
rect 230 320 238 322
rect 296 320 304 322
rect 363 321 371 323
rect 230 316 232 320
rect 236 316 238 320
rect 230 314 238 316
rect 296 316 304 318
rect 34 312 42 314
rect 4 310 12 312
rect 4 306 6 310
rect 10 306 12 310
rect 34 308 36 312
rect 40 308 42 312
rect 34 306 42 308
rect 44 312 52 314
rect 44 308 46 312
rect 50 308 52 312
rect 44 306 52 308
rect 64 312 72 314
rect 64 308 66 312
rect 70 308 72 312
rect 296 312 298 316
rect 302 312 304 316
rect 363 317 365 321
rect 369 317 371 321
rect 363 315 371 317
rect 373 321 381 323
rect 373 317 375 321
rect 379 317 381 321
rect 373 315 381 317
rect 383 321 391 323
rect 383 317 385 321
rect 389 317 391 321
rect 383 315 391 317
rect 393 321 401 323
rect 393 317 395 321
rect 399 317 401 321
rect 393 315 401 317
rect 403 321 411 323
rect 403 317 405 321
rect 409 317 411 321
rect 403 315 411 317
rect 413 321 421 323
rect 413 317 415 321
rect 419 317 421 321
rect 413 315 421 317
rect 423 321 431 323
rect 423 317 425 321
rect 429 317 431 321
rect 423 315 431 317
rect 433 321 441 323
rect 433 317 435 321
rect 439 317 441 321
rect 433 315 441 317
rect 443 321 451 323
rect 443 317 445 321
rect 449 317 451 321
rect 443 315 451 317
rect 453 321 461 323
rect 453 317 455 321
rect 459 317 461 321
rect 453 315 461 317
rect 463 321 471 323
rect 463 317 465 321
rect 469 317 471 321
rect 463 315 471 317
rect 473 321 481 323
rect 473 317 475 321
rect 479 317 481 321
rect 473 315 481 317
rect 483 321 491 323
rect 483 317 485 321
rect 489 317 491 321
rect 483 315 491 317
rect 528 322 536 324
rect 542 323 550 325
rect 552 329 560 331
rect 580 330 588 332
rect 552 325 554 329
rect 558 325 560 329
rect 552 323 560 325
rect 564 327 572 329
rect 564 323 566 327
rect 570 323 572 327
rect 580 326 582 330
rect 586 326 588 330
rect 580 324 588 326
rect 590 330 598 332
rect 590 326 592 330
rect 596 326 598 330
rect 590 324 598 326
rect 528 318 530 322
rect 534 318 536 322
rect 564 321 572 323
rect 528 316 536 318
rect 542 319 550 321
rect 542 315 544 319
rect 548 315 550 319
rect 296 310 304 312
rect 528 312 536 314
rect 542 313 550 315
rect 552 319 560 321
rect 580 320 588 322
rect 552 315 554 319
rect 558 315 560 319
rect 552 313 560 315
rect 564 317 572 319
rect 564 313 566 317
rect 570 313 572 317
rect 580 316 582 320
rect 586 316 588 320
rect 580 314 588 316
rect 590 320 598 322
rect 590 316 592 320
rect 596 316 598 320
rect 590 314 598 316
rect 528 308 530 312
rect 534 308 536 312
rect 564 311 572 313
rect 64 306 72 308
rect 296 306 304 308
rect 528 306 536 308
rect 542 309 550 311
rect 4 304 12 306
rect 34 302 42 304
rect 4 300 12 302
rect 4 296 6 300
rect 10 296 12 300
rect 34 298 36 302
rect 40 298 42 302
rect 34 296 42 298
rect 44 302 52 304
rect 44 298 46 302
rect 50 298 52 302
rect 44 296 52 298
rect 64 302 72 304
rect 64 298 66 302
rect 70 298 72 302
rect 296 302 298 306
rect 302 302 304 306
rect 542 305 544 309
rect 548 305 550 309
rect 296 300 304 302
rect 528 302 536 304
rect 542 303 550 305
rect 552 309 560 311
rect 580 310 588 312
rect 552 305 554 309
rect 558 305 560 309
rect 552 303 560 305
rect 564 307 572 309
rect 564 303 566 307
rect 570 303 572 307
rect 580 306 582 310
rect 586 306 588 310
rect 580 304 588 306
rect 590 310 598 312
rect 590 306 592 310
rect 596 306 598 310
rect 590 304 598 306
rect 64 296 72 298
rect 528 298 530 302
rect 534 298 536 302
rect 564 301 572 303
rect 528 296 536 298
rect 542 299 550 301
rect 4 294 12 296
rect 110 294 118 296
rect 34 292 42 294
rect 4 290 12 292
rect 4 286 6 290
rect 10 286 12 290
rect 34 288 36 292
rect 40 288 42 292
rect 34 286 42 288
rect 44 292 52 294
rect 44 288 46 292
rect 50 288 52 292
rect 44 286 52 288
rect 64 292 72 294
rect 64 288 66 292
rect 70 288 72 292
rect 110 290 112 294
rect 116 290 118 294
rect 110 288 118 290
rect 120 294 128 296
rect 120 290 122 294
rect 126 290 128 294
rect 120 288 128 290
rect 130 294 138 296
rect 130 290 132 294
rect 136 290 138 294
rect 130 288 138 290
rect 140 294 148 296
rect 140 290 142 294
rect 146 290 148 294
rect 140 288 148 290
rect 150 294 158 296
rect 150 290 152 294
rect 156 290 158 294
rect 150 288 158 290
rect 160 294 168 296
rect 160 290 162 294
rect 166 290 168 294
rect 160 288 168 290
rect 170 294 178 296
rect 170 290 172 294
rect 176 290 178 294
rect 170 288 178 290
rect 180 294 188 296
rect 180 290 182 294
rect 186 290 188 294
rect 180 288 188 290
rect 190 294 198 296
rect 190 290 192 294
rect 196 290 198 294
rect 190 288 198 290
rect 200 294 208 296
rect 200 290 202 294
rect 206 290 208 294
rect 200 288 208 290
rect 210 294 218 296
rect 210 290 212 294
rect 216 290 218 294
rect 210 288 218 290
rect 220 294 228 296
rect 220 290 222 294
rect 226 290 228 294
rect 220 288 228 290
rect 230 294 238 296
rect 230 290 232 294
rect 236 290 238 294
rect 230 288 238 290
rect 363 294 371 296
rect 363 290 365 294
rect 369 290 371 294
rect 363 288 371 290
rect 373 294 381 296
rect 373 290 375 294
rect 379 290 381 294
rect 373 288 381 290
rect 383 294 391 296
rect 383 290 385 294
rect 389 290 391 294
rect 383 288 391 290
rect 393 294 401 296
rect 393 290 395 294
rect 399 290 401 294
rect 393 288 401 290
rect 403 294 411 296
rect 403 290 405 294
rect 409 290 411 294
rect 403 288 411 290
rect 413 294 421 296
rect 413 290 415 294
rect 419 290 421 294
rect 413 288 421 290
rect 423 294 431 296
rect 423 290 425 294
rect 429 290 431 294
rect 423 288 431 290
rect 433 294 441 296
rect 433 290 435 294
rect 439 290 441 294
rect 433 288 441 290
rect 443 294 451 296
rect 443 290 445 294
rect 449 290 451 294
rect 443 288 451 290
rect 453 294 461 296
rect 453 290 455 294
rect 459 290 461 294
rect 453 288 461 290
rect 463 294 471 296
rect 463 290 465 294
rect 469 290 471 294
rect 463 288 471 290
rect 473 294 481 296
rect 473 290 475 294
rect 479 290 481 294
rect 473 288 481 290
rect 483 294 491 296
rect 542 295 544 299
rect 548 295 550 299
rect 483 290 485 294
rect 489 290 491 294
rect 483 288 491 290
rect 528 292 536 294
rect 542 293 550 295
rect 552 299 560 301
rect 580 300 588 302
rect 552 295 554 299
rect 558 295 560 299
rect 552 293 560 295
rect 564 297 572 299
rect 564 293 566 297
rect 570 293 572 297
rect 580 296 582 300
rect 586 296 588 300
rect 580 294 588 296
rect 590 300 598 302
rect 590 296 592 300
rect 596 296 598 300
rect 590 294 598 296
rect 528 288 530 292
rect 534 288 536 292
rect 564 291 572 293
rect 64 286 72 288
rect 296 286 304 288
rect 528 286 536 288
rect 542 289 550 291
rect 4 284 12 286
rect 34 282 42 284
rect 4 280 12 282
rect 4 276 6 280
rect 10 276 12 280
rect 34 278 36 282
rect 40 278 42 282
rect 34 276 42 278
rect 44 282 52 284
rect 44 278 46 282
rect 50 278 52 282
rect 44 276 52 278
rect 64 282 72 284
rect 64 278 66 282
rect 70 278 72 282
rect 296 282 298 286
rect 302 282 304 286
rect 542 285 544 289
rect 548 285 550 289
rect 296 280 304 282
rect 528 282 536 284
rect 542 283 550 285
rect 552 289 560 291
rect 580 290 588 292
rect 552 285 554 289
rect 558 285 560 289
rect 552 283 560 285
rect 564 287 572 289
rect 564 283 566 287
rect 570 283 572 287
rect 580 286 582 290
rect 586 286 588 290
rect 580 284 588 286
rect 590 290 598 292
rect 590 286 592 290
rect 596 286 598 290
rect 590 284 598 286
rect 528 278 530 282
rect 534 278 536 282
rect 564 281 572 283
rect 64 276 72 278
rect 296 276 304 278
rect 528 276 536 278
rect 542 279 550 281
rect 4 274 12 276
rect 34 272 42 274
rect 4 270 12 272
rect 4 266 6 270
rect 10 266 12 270
rect 34 268 36 272
rect 40 268 42 272
rect 34 266 42 268
rect 44 272 52 274
rect 44 268 46 272
rect 50 268 52 272
rect 44 266 52 268
rect 64 272 72 274
rect 64 268 66 272
rect 70 268 72 272
rect 296 272 298 276
rect 302 272 304 276
rect 542 275 544 279
rect 548 275 550 279
rect 296 270 304 272
rect 528 272 536 274
rect 542 273 550 275
rect 552 279 560 281
rect 580 280 588 282
rect 552 275 554 279
rect 558 275 560 279
rect 552 273 560 275
rect 564 277 572 279
rect 564 273 566 277
rect 570 273 572 277
rect 580 276 582 280
rect 586 276 588 280
rect 580 274 588 276
rect 590 280 598 282
rect 590 276 592 280
rect 596 276 598 280
rect 590 274 598 276
rect 528 268 530 272
rect 534 268 536 272
rect 564 271 572 273
rect 64 266 72 268
rect 112 266 120 268
rect 4 264 12 266
rect 34 262 42 264
rect 4 260 12 262
rect 4 256 6 260
rect 10 256 12 260
rect 34 258 36 262
rect 40 258 42 262
rect 34 256 42 258
rect 44 262 52 264
rect 44 258 46 262
rect 50 258 52 262
rect 44 256 52 258
rect 64 262 72 264
rect 64 258 66 262
rect 70 258 72 262
rect 112 262 114 266
rect 118 262 120 266
rect 112 260 120 262
rect 122 266 130 268
rect 122 262 124 266
rect 128 262 130 266
rect 122 260 130 262
rect 132 266 140 268
rect 132 262 134 266
rect 138 262 140 266
rect 132 260 140 262
rect 142 266 150 268
rect 142 262 144 266
rect 148 262 150 266
rect 142 260 150 262
rect 152 266 160 268
rect 152 262 154 266
rect 158 262 160 266
rect 152 260 160 262
rect 162 266 170 268
rect 162 262 164 266
rect 168 262 170 266
rect 162 260 170 262
rect 172 266 180 268
rect 172 262 174 266
rect 178 262 180 266
rect 172 260 180 262
rect 182 266 190 268
rect 182 262 184 266
rect 188 262 190 266
rect 182 260 190 262
rect 192 266 200 268
rect 192 262 194 266
rect 198 262 200 266
rect 192 260 200 262
rect 202 266 210 268
rect 202 262 204 266
rect 208 262 210 266
rect 202 260 210 262
rect 212 266 220 268
rect 212 262 214 266
rect 218 262 220 266
rect 212 260 220 262
rect 222 266 230 268
rect 222 262 224 266
rect 228 262 230 266
rect 222 260 230 262
rect 232 266 240 268
rect 232 262 234 266
rect 238 262 240 266
rect 232 260 240 262
rect 296 266 304 268
rect 296 262 298 266
rect 302 262 304 266
rect 296 260 304 262
rect 360 266 368 268
rect 360 262 362 266
rect 366 262 368 266
rect 360 260 368 262
rect 370 266 378 268
rect 370 262 372 266
rect 376 262 378 266
rect 370 260 378 262
rect 380 266 388 268
rect 380 262 382 266
rect 386 262 388 266
rect 380 260 388 262
rect 390 266 398 268
rect 390 262 392 266
rect 396 262 398 266
rect 390 260 398 262
rect 400 266 408 268
rect 400 262 402 266
rect 406 262 408 266
rect 400 260 408 262
rect 410 266 418 268
rect 410 262 412 266
rect 416 262 418 266
rect 410 260 418 262
rect 420 266 428 268
rect 420 262 422 266
rect 426 262 428 266
rect 420 260 428 262
rect 430 266 438 268
rect 430 262 432 266
rect 436 262 438 266
rect 430 260 438 262
rect 440 266 448 268
rect 440 262 442 266
rect 446 262 448 266
rect 440 260 448 262
rect 450 266 458 268
rect 450 262 452 266
rect 456 262 458 266
rect 450 260 458 262
rect 460 266 468 268
rect 460 262 462 266
rect 466 262 468 266
rect 460 260 468 262
rect 470 266 478 268
rect 470 262 472 266
rect 476 262 478 266
rect 470 260 478 262
rect 480 266 488 268
rect 528 266 536 268
rect 542 269 550 271
rect 480 262 482 266
rect 486 262 488 266
rect 542 265 544 269
rect 548 265 550 269
rect 480 260 488 262
rect 528 262 536 264
rect 542 263 550 265
rect 552 269 560 271
rect 580 270 588 272
rect 552 265 554 269
rect 558 265 560 269
rect 552 263 560 265
rect 564 267 572 269
rect 564 263 566 267
rect 570 263 572 267
rect 580 266 582 270
rect 586 266 588 270
rect 580 264 588 266
rect 590 270 598 272
rect 590 266 592 270
rect 596 266 598 270
rect 590 264 598 266
rect 528 258 530 262
rect 534 258 536 262
rect 564 261 572 263
rect 64 256 72 258
rect 112 256 120 258
rect 4 254 12 256
rect 34 252 42 254
rect 4 250 12 252
rect 4 246 6 250
rect 10 246 12 250
rect 34 248 36 252
rect 40 248 42 252
rect 34 246 42 248
rect 44 252 52 254
rect 44 248 46 252
rect 50 248 52 252
rect 44 246 52 248
rect 64 252 72 254
rect 64 248 66 252
rect 70 248 72 252
rect 112 252 114 256
rect 118 252 120 256
rect 112 250 120 252
rect 122 256 130 258
rect 122 252 124 256
rect 128 252 130 256
rect 122 250 130 252
rect 132 256 140 258
rect 132 252 134 256
rect 138 252 140 256
rect 132 250 140 252
rect 142 256 150 258
rect 142 252 144 256
rect 148 252 150 256
rect 142 250 150 252
rect 152 256 160 258
rect 152 252 154 256
rect 158 252 160 256
rect 152 250 160 252
rect 162 256 170 258
rect 162 252 164 256
rect 168 252 170 256
rect 162 250 170 252
rect 172 256 180 258
rect 172 252 174 256
rect 178 252 180 256
rect 172 250 180 252
rect 182 256 190 258
rect 182 252 184 256
rect 188 252 190 256
rect 182 250 190 252
rect 192 256 200 258
rect 192 252 194 256
rect 198 252 200 256
rect 192 250 200 252
rect 202 256 210 258
rect 202 252 204 256
rect 208 252 210 256
rect 202 250 210 252
rect 212 256 220 258
rect 212 252 214 256
rect 218 252 220 256
rect 212 250 220 252
rect 222 256 230 258
rect 222 252 224 256
rect 228 252 230 256
rect 222 250 230 252
rect 232 256 240 258
rect 232 252 234 256
rect 238 252 240 256
rect 232 250 240 252
rect 296 256 304 258
rect 296 252 298 256
rect 302 252 304 256
rect 296 250 304 252
rect 360 256 368 258
rect 360 252 362 256
rect 366 252 368 256
rect 360 250 368 252
rect 370 256 378 258
rect 370 252 372 256
rect 376 252 378 256
rect 370 250 378 252
rect 380 256 388 258
rect 380 252 382 256
rect 386 252 388 256
rect 380 250 388 252
rect 390 256 398 258
rect 390 252 392 256
rect 396 252 398 256
rect 390 250 398 252
rect 400 256 408 258
rect 400 252 402 256
rect 406 252 408 256
rect 400 250 408 252
rect 410 256 418 258
rect 410 252 412 256
rect 416 252 418 256
rect 410 250 418 252
rect 420 256 428 258
rect 420 252 422 256
rect 426 252 428 256
rect 420 250 428 252
rect 430 256 438 258
rect 430 252 432 256
rect 436 252 438 256
rect 430 250 438 252
rect 440 256 448 258
rect 440 252 442 256
rect 446 252 448 256
rect 440 250 448 252
rect 450 256 458 258
rect 450 252 452 256
rect 456 252 458 256
rect 450 250 458 252
rect 460 256 468 258
rect 460 252 462 256
rect 466 252 468 256
rect 460 250 468 252
rect 470 256 478 258
rect 470 252 472 256
rect 476 252 478 256
rect 470 250 478 252
rect 480 256 488 258
rect 528 256 536 258
rect 542 259 550 261
rect 480 252 482 256
rect 486 252 488 256
rect 542 255 544 259
rect 548 255 550 259
rect 480 250 488 252
rect 528 252 536 254
rect 542 253 550 255
rect 552 259 560 261
rect 580 260 588 262
rect 552 255 554 259
rect 558 255 560 259
rect 552 253 560 255
rect 564 257 572 259
rect 564 253 566 257
rect 570 253 572 257
rect 580 256 582 260
rect 586 256 588 260
rect 580 254 588 256
rect 590 260 598 262
rect 590 256 592 260
rect 596 256 598 260
rect 590 254 598 256
rect 528 248 530 252
rect 534 248 536 252
rect 564 251 572 253
rect 64 246 72 248
rect 296 246 304 248
rect 528 246 536 248
rect 542 249 550 251
rect 4 244 12 246
rect 34 242 42 244
rect 4 240 12 242
rect 4 236 6 240
rect 10 236 12 240
rect 34 238 36 242
rect 40 238 42 242
rect 34 236 42 238
rect 44 242 52 244
rect 44 238 46 242
rect 50 238 52 242
rect 44 236 52 238
rect 64 242 72 244
rect 64 238 66 242
rect 70 238 72 242
rect 296 242 298 246
rect 302 242 304 246
rect 542 245 544 249
rect 548 245 550 249
rect 296 240 304 242
rect 528 242 536 244
rect 542 243 550 245
rect 552 249 560 251
rect 580 250 588 252
rect 552 245 554 249
rect 558 245 560 249
rect 552 243 560 245
rect 564 247 572 249
rect 564 243 566 247
rect 570 243 572 247
rect 580 246 582 250
rect 586 246 588 250
rect 580 244 588 246
rect 590 250 598 252
rect 590 246 592 250
rect 596 246 598 250
rect 590 244 598 246
rect 528 238 530 242
rect 534 238 536 242
rect 564 241 572 243
rect 64 236 72 238
rect 296 236 304 238
rect 528 236 536 238
rect 542 239 550 241
rect 4 234 12 236
rect 34 232 42 234
rect 4 230 12 232
rect 4 226 6 230
rect 10 226 12 230
rect 34 228 36 232
rect 40 228 42 232
rect 34 226 42 228
rect 44 232 52 234
rect 44 228 46 232
rect 50 228 52 232
rect 44 226 52 228
rect 64 232 72 234
rect 296 232 298 236
rect 302 232 304 236
rect 542 235 544 239
rect 548 235 550 239
rect 64 228 66 232
rect 70 228 72 232
rect 64 226 72 228
rect 110 230 118 232
rect 110 226 112 230
rect 116 226 118 230
rect 4 224 12 226
rect 110 224 118 226
rect 120 230 128 232
rect 120 226 122 230
rect 126 226 128 230
rect 120 224 128 226
rect 130 230 138 232
rect 130 226 132 230
rect 136 226 138 230
rect 130 224 138 226
rect 140 230 148 232
rect 140 226 142 230
rect 146 226 148 230
rect 140 224 148 226
rect 150 230 158 232
rect 150 226 152 230
rect 156 226 158 230
rect 150 224 158 226
rect 160 230 168 232
rect 160 226 162 230
rect 166 226 168 230
rect 160 224 168 226
rect 170 230 178 232
rect 170 226 172 230
rect 176 226 178 230
rect 170 224 178 226
rect 180 230 188 232
rect 180 226 182 230
rect 186 226 188 230
rect 180 224 188 226
rect 190 230 198 232
rect 190 226 192 230
rect 196 226 198 230
rect 190 224 198 226
rect 200 230 208 232
rect 200 226 202 230
rect 206 226 208 230
rect 200 224 208 226
rect 210 230 218 232
rect 210 226 212 230
rect 216 226 218 230
rect 210 224 218 226
rect 220 230 228 232
rect 220 226 222 230
rect 226 226 228 230
rect 220 224 228 226
rect 230 230 238 232
rect 296 230 304 232
rect 528 232 536 234
rect 542 233 550 235
rect 552 239 560 241
rect 580 240 588 242
rect 552 235 554 239
rect 558 235 560 239
rect 552 233 560 235
rect 564 237 572 239
rect 564 233 566 237
rect 570 233 572 237
rect 580 236 582 240
rect 586 236 588 240
rect 580 234 588 236
rect 590 240 598 242
rect 590 236 592 240
rect 596 236 598 240
rect 590 234 598 236
rect 230 226 232 230
rect 236 226 238 230
rect 364 229 372 231
rect 230 224 238 226
rect 296 226 304 228
rect 34 222 42 224
rect 4 220 12 222
rect 4 216 6 220
rect 10 216 12 220
rect 34 218 36 222
rect 40 218 42 222
rect 34 216 42 218
rect 44 222 52 224
rect 44 218 46 222
rect 50 218 52 222
rect 44 216 52 218
rect 64 222 72 224
rect 64 218 66 222
rect 70 218 72 222
rect 296 222 298 226
rect 302 222 304 226
rect 364 225 366 229
rect 370 225 372 229
rect 364 223 372 225
rect 374 229 382 231
rect 374 225 376 229
rect 380 225 382 229
rect 374 223 382 225
rect 384 229 392 231
rect 384 225 386 229
rect 390 225 392 229
rect 384 223 392 225
rect 394 229 402 231
rect 394 225 396 229
rect 400 225 402 229
rect 394 223 402 225
rect 404 229 412 231
rect 404 225 406 229
rect 410 225 412 229
rect 404 223 412 225
rect 414 229 422 231
rect 414 225 416 229
rect 420 225 422 229
rect 414 223 422 225
rect 424 229 432 231
rect 424 225 426 229
rect 430 225 432 229
rect 424 223 432 225
rect 434 229 442 231
rect 434 225 436 229
rect 440 225 442 229
rect 434 223 442 225
rect 444 229 452 231
rect 444 225 446 229
rect 450 225 452 229
rect 444 223 452 225
rect 454 229 462 231
rect 454 225 456 229
rect 460 225 462 229
rect 454 223 462 225
rect 464 229 472 231
rect 464 225 466 229
rect 470 225 472 229
rect 464 223 472 225
rect 474 229 482 231
rect 474 225 476 229
rect 480 225 482 229
rect 474 223 482 225
rect 484 229 492 231
rect 484 225 486 229
rect 490 225 492 229
rect 528 228 530 232
rect 534 228 536 232
rect 564 231 572 233
rect 528 226 536 228
rect 542 229 550 231
rect 484 223 492 225
rect 542 225 544 229
rect 548 225 550 229
rect 296 220 304 222
rect 528 222 536 224
rect 542 223 550 225
rect 552 229 560 231
rect 580 230 588 232
rect 552 225 554 229
rect 558 225 560 229
rect 552 223 560 225
rect 564 227 572 229
rect 564 223 566 227
rect 570 223 572 227
rect 580 226 582 230
rect 586 226 588 230
rect 580 224 588 226
rect 590 230 598 232
rect 590 226 592 230
rect 596 226 598 230
rect 590 224 598 226
rect 528 218 530 222
rect 534 218 536 222
rect 564 221 572 223
rect 64 216 72 218
rect 296 216 304 218
rect 528 216 536 218
rect 542 219 550 221
rect 4 214 12 216
rect 34 212 42 214
rect 4 210 12 212
rect 4 206 6 210
rect 10 206 12 210
rect 34 208 36 212
rect 40 208 42 212
rect 34 206 42 208
rect 44 212 52 214
rect 44 208 46 212
rect 50 208 52 212
rect 44 206 52 208
rect 64 212 72 214
rect 64 208 66 212
rect 70 208 72 212
rect 296 212 298 216
rect 302 212 304 216
rect 542 215 544 219
rect 548 215 550 219
rect 296 210 304 212
rect 528 212 536 214
rect 542 213 550 215
rect 552 219 560 221
rect 580 220 588 222
rect 552 215 554 219
rect 558 215 560 219
rect 552 213 560 215
rect 564 217 572 219
rect 564 213 566 217
rect 570 213 572 217
rect 580 216 582 220
rect 586 216 588 220
rect 580 214 588 216
rect 590 220 598 222
rect 590 216 592 220
rect 596 216 598 220
rect 590 214 598 216
rect 528 208 530 212
rect 534 208 536 212
rect 564 211 572 213
rect 64 206 72 208
rect 296 206 304 208
rect 528 206 536 208
rect 542 209 550 211
rect 4 204 12 206
rect 34 202 42 204
rect 4 200 12 202
rect 4 196 6 200
rect 10 196 12 200
rect 34 198 36 202
rect 40 198 42 202
rect 34 196 42 198
rect 44 202 52 204
rect 44 198 46 202
rect 50 198 52 202
rect 44 196 52 198
rect 64 202 72 204
rect 64 198 66 202
rect 70 198 72 202
rect 64 196 72 198
rect 109 202 117 204
rect 109 198 111 202
rect 115 198 117 202
rect 109 196 117 198
rect 119 202 127 204
rect 119 198 121 202
rect 125 198 127 202
rect 119 196 127 198
rect 129 202 137 204
rect 129 198 131 202
rect 135 198 137 202
rect 129 196 137 198
rect 139 202 147 204
rect 139 198 141 202
rect 145 198 147 202
rect 139 196 147 198
rect 149 202 157 204
rect 149 198 151 202
rect 155 198 157 202
rect 149 196 157 198
rect 159 202 167 204
rect 159 198 161 202
rect 165 198 167 202
rect 159 196 167 198
rect 169 202 177 204
rect 169 198 171 202
rect 175 198 177 202
rect 169 196 177 198
rect 179 202 187 204
rect 179 198 181 202
rect 185 198 187 202
rect 179 196 187 198
rect 189 202 197 204
rect 189 198 191 202
rect 195 198 197 202
rect 189 196 197 198
rect 199 202 207 204
rect 199 198 201 202
rect 205 198 207 202
rect 199 196 207 198
rect 209 202 217 204
rect 209 198 211 202
rect 215 198 217 202
rect 209 196 217 198
rect 219 202 227 204
rect 219 198 221 202
rect 225 198 227 202
rect 219 196 227 198
rect 229 202 237 204
rect 229 198 231 202
rect 235 198 237 202
rect 296 202 298 206
rect 302 202 304 206
rect 542 205 544 209
rect 548 205 550 209
rect 296 200 304 202
rect 364 202 372 204
rect 364 198 366 202
rect 370 198 372 202
rect 229 196 237 198
rect 296 196 304 198
rect 364 196 372 198
rect 374 202 382 204
rect 374 198 376 202
rect 380 198 382 202
rect 374 196 382 198
rect 384 202 392 204
rect 384 198 386 202
rect 390 198 392 202
rect 384 196 392 198
rect 394 202 402 204
rect 394 198 396 202
rect 400 198 402 202
rect 394 196 402 198
rect 404 202 412 204
rect 404 198 406 202
rect 410 198 412 202
rect 404 196 412 198
rect 414 202 422 204
rect 414 198 416 202
rect 420 198 422 202
rect 414 196 422 198
rect 424 202 432 204
rect 424 198 426 202
rect 430 198 432 202
rect 424 196 432 198
rect 434 202 442 204
rect 434 198 436 202
rect 440 198 442 202
rect 434 196 442 198
rect 444 202 452 204
rect 444 198 446 202
rect 450 198 452 202
rect 444 196 452 198
rect 454 202 462 204
rect 454 198 456 202
rect 460 198 462 202
rect 454 196 462 198
rect 464 202 472 204
rect 464 198 466 202
rect 470 198 472 202
rect 464 196 472 198
rect 474 202 482 204
rect 474 198 476 202
rect 480 198 482 202
rect 474 196 482 198
rect 484 202 492 204
rect 484 198 486 202
rect 490 198 492 202
rect 484 196 492 198
rect 528 202 536 204
rect 542 203 550 205
rect 552 209 560 211
rect 580 210 588 212
rect 552 205 554 209
rect 558 205 560 209
rect 552 203 560 205
rect 564 207 572 209
rect 564 203 566 207
rect 570 203 572 207
rect 580 206 582 210
rect 586 206 588 210
rect 580 204 588 206
rect 590 210 598 212
rect 590 206 592 210
rect 596 206 598 210
rect 590 204 598 206
rect 528 198 530 202
rect 534 198 536 202
rect 564 201 572 203
rect 528 196 536 198
rect 542 199 550 201
rect 4 194 12 196
rect 34 192 42 194
rect 4 190 12 192
rect 4 186 6 190
rect 10 186 12 190
rect 34 188 36 192
rect 40 188 42 192
rect 34 186 42 188
rect 44 192 52 194
rect 44 188 46 192
rect 50 188 52 192
rect 44 186 52 188
rect 64 192 72 194
rect 296 192 298 196
rect 302 192 304 196
rect 542 195 544 199
rect 548 195 550 199
rect 528 192 536 194
rect 542 193 550 195
rect 552 199 560 201
rect 580 200 588 202
rect 552 195 554 199
rect 558 195 560 199
rect 552 193 560 195
rect 564 197 572 199
rect 564 193 566 197
rect 570 193 572 197
rect 580 196 582 200
rect 586 196 588 200
rect 580 194 588 196
rect 590 200 598 202
rect 590 196 592 200
rect 596 196 598 200
rect 590 194 598 196
rect 64 188 66 192
rect 70 188 72 192
rect 64 186 72 188
rect 109 190 117 192
rect 109 186 111 190
rect 115 186 117 190
rect 4 184 12 186
rect 109 184 117 186
rect 119 190 127 192
rect 119 186 121 190
rect 125 186 127 190
rect 119 184 127 186
rect 129 190 137 192
rect 129 186 131 190
rect 135 186 137 190
rect 129 184 137 186
rect 139 190 147 192
rect 139 186 141 190
rect 145 186 147 190
rect 139 184 147 186
rect 149 190 157 192
rect 149 186 151 190
rect 155 186 157 190
rect 149 184 157 186
rect 159 190 167 192
rect 159 186 161 190
rect 165 186 167 190
rect 159 184 167 186
rect 169 190 177 192
rect 169 186 171 190
rect 175 186 177 190
rect 169 184 177 186
rect 179 190 187 192
rect 179 186 181 190
rect 185 186 187 190
rect 179 184 187 186
rect 189 190 197 192
rect 189 186 191 190
rect 195 186 197 190
rect 189 184 197 186
rect 199 190 207 192
rect 199 186 201 190
rect 205 186 207 190
rect 199 184 207 186
rect 209 190 217 192
rect 209 186 211 190
rect 215 186 217 190
rect 209 184 217 186
rect 219 190 227 192
rect 219 186 221 190
rect 225 186 227 190
rect 219 184 227 186
rect 229 190 237 192
rect 296 190 304 192
rect 364 190 372 192
rect 229 186 231 190
rect 235 186 237 190
rect 229 184 237 186
rect 296 186 304 188
rect 34 182 42 184
rect 4 180 12 182
rect 4 176 6 180
rect 10 176 12 180
rect 34 178 36 182
rect 40 178 42 182
rect 34 176 42 178
rect 44 182 52 184
rect 44 178 46 182
rect 50 178 52 182
rect 44 176 52 178
rect 64 182 72 184
rect 64 178 66 182
rect 70 178 72 182
rect 296 182 298 186
rect 302 182 304 186
rect 364 186 366 190
rect 370 186 372 190
rect 364 184 372 186
rect 374 190 382 192
rect 374 186 376 190
rect 380 186 382 190
rect 374 184 382 186
rect 384 190 392 192
rect 384 186 386 190
rect 390 186 392 190
rect 384 184 392 186
rect 394 190 402 192
rect 394 186 396 190
rect 400 186 402 190
rect 394 184 402 186
rect 404 190 412 192
rect 404 186 406 190
rect 410 186 412 190
rect 404 184 412 186
rect 414 190 422 192
rect 414 186 416 190
rect 420 186 422 190
rect 414 184 422 186
rect 424 190 432 192
rect 424 186 426 190
rect 430 186 432 190
rect 424 184 432 186
rect 434 190 442 192
rect 434 186 436 190
rect 440 186 442 190
rect 434 184 442 186
rect 444 190 452 192
rect 444 186 446 190
rect 450 186 452 190
rect 444 184 452 186
rect 454 190 462 192
rect 454 186 456 190
rect 460 186 462 190
rect 454 184 462 186
rect 464 190 472 192
rect 464 186 466 190
rect 470 186 472 190
rect 464 184 472 186
rect 474 190 482 192
rect 474 186 476 190
rect 480 186 482 190
rect 474 184 482 186
rect 484 190 492 192
rect 484 186 486 190
rect 490 186 492 190
rect 528 188 530 192
rect 534 188 536 192
rect 564 191 572 193
rect 528 186 536 188
rect 542 189 550 191
rect 484 184 492 186
rect 542 185 544 189
rect 548 185 550 189
rect 296 180 304 182
rect 528 182 536 184
rect 542 183 550 185
rect 552 189 560 191
rect 580 190 588 192
rect 552 185 554 189
rect 558 185 560 189
rect 552 183 560 185
rect 564 187 572 189
rect 564 183 566 187
rect 570 183 572 187
rect 580 186 582 190
rect 586 186 588 190
rect 580 184 588 186
rect 590 190 598 192
rect 590 186 592 190
rect 596 186 598 190
rect 590 184 598 186
rect 528 178 530 182
rect 534 178 536 182
rect 564 181 572 183
rect 64 176 72 178
rect 296 176 304 178
rect 528 176 536 178
rect 542 179 550 181
rect 4 174 12 176
rect 34 172 42 174
rect 4 170 12 172
rect 4 166 6 170
rect 10 166 12 170
rect 34 168 36 172
rect 40 168 42 172
rect 34 166 42 168
rect 44 172 52 174
rect 44 168 46 172
rect 50 168 52 172
rect 44 166 52 168
rect 64 172 72 174
rect 64 168 66 172
rect 70 168 72 172
rect 296 172 298 176
rect 302 172 304 176
rect 542 175 544 179
rect 548 175 550 179
rect 296 170 304 172
rect 528 172 536 174
rect 542 173 550 175
rect 552 179 560 181
rect 580 180 588 182
rect 552 175 554 179
rect 558 175 560 179
rect 552 173 560 175
rect 564 177 572 179
rect 564 173 566 177
rect 570 173 572 177
rect 580 176 582 180
rect 586 176 588 180
rect 580 174 588 176
rect 590 180 598 182
rect 590 176 592 180
rect 596 176 598 180
rect 590 174 598 176
rect 528 168 530 172
rect 534 168 536 172
rect 564 171 572 173
rect 64 166 72 168
rect 110 166 118 168
rect 4 164 12 166
rect 34 162 42 164
rect 4 160 12 162
rect 4 156 6 160
rect 10 156 12 160
rect 34 158 36 162
rect 40 158 42 162
rect 34 156 42 158
rect 44 162 52 164
rect 44 158 46 162
rect 50 158 52 162
rect 44 156 52 158
rect 64 162 72 164
rect 64 158 66 162
rect 70 158 72 162
rect 110 162 112 166
rect 116 162 118 166
rect 110 160 118 162
rect 120 166 128 168
rect 120 162 122 166
rect 126 162 128 166
rect 120 160 128 162
rect 130 166 138 168
rect 130 162 132 166
rect 136 162 138 166
rect 130 160 138 162
rect 140 166 148 168
rect 140 162 142 166
rect 146 162 148 166
rect 140 160 148 162
rect 150 166 158 168
rect 150 162 152 166
rect 156 162 158 166
rect 150 160 158 162
rect 160 166 168 168
rect 160 162 162 166
rect 166 162 168 166
rect 160 160 168 162
rect 170 166 178 168
rect 170 162 172 166
rect 176 162 178 166
rect 170 160 178 162
rect 180 166 188 168
rect 180 162 182 166
rect 186 162 188 166
rect 180 160 188 162
rect 190 166 198 168
rect 190 162 192 166
rect 196 162 198 166
rect 190 160 198 162
rect 200 166 208 168
rect 200 162 202 166
rect 206 162 208 166
rect 200 160 208 162
rect 210 166 218 168
rect 210 162 212 166
rect 216 162 218 166
rect 210 160 218 162
rect 220 166 228 168
rect 220 162 222 166
rect 226 162 228 166
rect 220 160 228 162
rect 230 166 238 168
rect 230 162 232 166
rect 236 162 238 166
rect 230 160 238 162
rect 364 166 372 168
rect 364 162 366 166
rect 370 162 372 166
rect 364 160 372 162
rect 374 166 382 168
rect 374 162 376 166
rect 380 162 382 166
rect 374 160 382 162
rect 384 166 392 168
rect 384 162 386 166
rect 390 162 392 166
rect 384 160 392 162
rect 394 166 402 168
rect 394 162 396 166
rect 400 162 402 166
rect 394 160 402 162
rect 404 166 412 168
rect 404 162 406 166
rect 410 162 412 166
rect 404 160 412 162
rect 414 166 422 168
rect 414 162 416 166
rect 420 162 422 166
rect 414 160 422 162
rect 424 166 432 168
rect 424 162 426 166
rect 430 162 432 166
rect 424 160 432 162
rect 434 166 442 168
rect 434 162 436 166
rect 440 162 442 166
rect 434 160 442 162
rect 444 166 452 168
rect 444 162 446 166
rect 450 162 452 166
rect 444 160 452 162
rect 454 166 462 168
rect 454 162 456 166
rect 460 162 462 166
rect 454 160 462 162
rect 464 166 472 168
rect 464 162 466 166
rect 470 162 472 166
rect 464 160 472 162
rect 474 166 482 168
rect 474 162 476 166
rect 480 162 482 166
rect 474 160 482 162
rect 484 166 492 168
rect 528 166 536 168
rect 542 169 550 171
rect 484 162 486 166
rect 490 162 492 166
rect 542 165 544 169
rect 548 165 550 169
rect 484 160 492 162
rect 528 162 536 164
rect 542 163 550 165
rect 552 169 560 171
rect 580 170 588 172
rect 552 165 554 169
rect 558 165 560 169
rect 552 163 560 165
rect 564 167 572 169
rect 564 163 566 167
rect 570 163 572 167
rect 580 166 582 170
rect 586 166 588 170
rect 580 164 588 166
rect 590 170 598 172
rect 590 166 592 170
rect 596 166 598 170
rect 590 164 598 166
rect 528 158 530 162
rect 534 158 536 162
rect 564 161 572 163
rect 64 156 72 158
rect 296 156 304 158
rect 528 156 536 158
rect 542 159 550 161
rect 4 154 12 156
rect 34 152 42 154
rect 4 150 12 152
rect 4 146 6 150
rect 10 146 12 150
rect 34 148 36 152
rect 40 148 42 152
rect 34 146 42 148
rect 44 152 52 154
rect 44 148 46 152
rect 50 148 52 152
rect 44 146 52 148
rect 64 152 72 154
rect 64 148 66 152
rect 70 148 72 152
rect 296 152 298 156
rect 302 152 304 156
rect 542 155 544 159
rect 548 155 550 159
rect 296 150 304 152
rect 528 152 536 154
rect 542 153 550 155
rect 552 159 560 161
rect 580 160 588 162
rect 552 155 554 159
rect 558 155 560 159
rect 552 153 560 155
rect 564 157 572 159
rect 564 153 566 157
rect 570 153 572 157
rect 580 156 582 160
rect 586 156 588 160
rect 580 154 588 156
rect 590 160 598 162
rect 590 156 592 160
rect 596 156 598 160
rect 590 154 598 156
rect 528 148 530 152
rect 534 148 536 152
rect 564 151 572 153
rect 64 146 72 148
rect 296 146 304 148
rect 528 146 536 148
rect 542 149 550 151
rect 4 144 12 146
rect 34 142 42 144
rect 4 140 12 142
rect 4 136 6 140
rect 10 136 12 140
rect 34 138 36 142
rect 40 138 42 142
rect 34 136 42 138
rect 44 142 52 144
rect 44 138 46 142
rect 50 138 52 142
rect 44 136 52 138
rect 64 142 72 144
rect 64 138 66 142
rect 70 138 72 142
rect 296 142 298 146
rect 302 142 304 146
rect 542 145 544 149
rect 548 145 550 149
rect 296 140 304 142
rect 528 142 536 144
rect 542 143 550 145
rect 552 149 560 151
rect 580 150 588 152
rect 552 145 554 149
rect 558 145 560 149
rect 552 143 560 145
rect 564 147 572 149
rect 564 143 566 147
rect 570 143 572 147
rect 580 146 582 150
rect 586 146 588 150
rect 580 144 588 146
rect 590 150 598 152
rect 590 146 592 150
rect 596 146 598 150
rect 590 144 598 146
rect 528 138 530 142
rect 534 138 536 142
rect 564 141 572 143
rect 64 136 72 138
rect 112 136 120 138
rect 4 134 12 136
rect 34 132 42 134
rect 4 130 12 132
rect 4 126 6 130
rect 10 126 12 130
rect 34 128 36 132
rect 40 128 42 132
rect 34 126 42 128
rect 44 132 52 134
rect 44 128 46 132
rect 50 128 52 132
rect 44 126 52 128
rect 64 132 72 134
rect 64 128 66 132
rect 70 128 72 132
rect 112 132 114 136
rect 118 132 120 136
rect 112 130 120 132
rect 122 136 130 138
rect 122 132 124 136
rect 128 132 130 136
rect 122 130 130 132
rect 132 136 140 138
rect 132 132 134 136
rect 138 132 140 136
rect 132 130 140 132
rect 142 136 150 138
rect 142 132 144 136
rect 148 132 150 136
rect 142 130 150 132
rect 152 136 160 138
rect 152 132 154 136
rect 158 132 160 136
rect 152 130 160 132
rect 162 136 170 138
rect 162 132 164 136
rect 168 132 170 136
rect 162 130 170 132
rect 172 136 180 138
rect 172 132 174 136
rect 178 132 180 136
rect 172 130 180 132
rect 182 136 190 138
rect 182 132 184 136
rect 188 132 190 136
rect 182 130 190 132
rect 192 136 200 138
rect 192 132 194 136
rect 198 132 200 136
rect 192 130 200 132
rect 202 136 210 138
rect 202 132 204 136
rect 208 132 210 136
rect 202 130 210 132
rect 212 136 220 138
rect 212 132 214 136
rect 218 132 220 136
rect 212 130 220 132
rect 222 136 230 138
rect 222 132 224 136
rect 228 132 230 136
rect 222 130 230 132
rect 232 136 240 138
rect 232 132 234 136
rect 238 132 240 136
rect 232 130 240 132
rect 296 136 304 138
rect 296 132 298 136
rect 302 132 304 136
rect 296 130 304 132
rect 360 136 368 138
rect 360 132 362 136
rect 366 132 368 136
rect 360 130 368 132
rect 370 136 378 138
rect 370 132 372 136
rect 376 132 378 136
rect 370 130 378 132
rect 380 136 388 138
rect 380 132 382 136
rect 386 132 388 136
rect 380 130 388 132
rect 390 136 398 138
rect 390 132 392 136
rect 396 132 398 136
rect 390 130 398 132
rect 400 136 408 138
rect 400 132 402 136
rect 406 132 408 136
rect 400 130 408 132
rect 410 136 418 138
rect 410 132 412 136
rect 416 132 418 136
rect 410 130 418 132
rect 420 136 428 138
rect 420 132 422 136
rect 426 132 428 136
rect 420 130 428 132
rect 430 136 438 138
rect 430 132 432 136
rect 436 132 438 136
rect 430 130 438 132
rect 440 136 448 138
rect 440 132 442 136
rect 446 132 448 136
rect 440 130 448 132
rect 450 136 458 138
rect 450 132 452 136
rect 456 132 458 136
rect 450 130 458 132
rect 460 136 468 138
rect 460 132 462 136
rect 466 132 468 136
rect 460 130 468 132
rect 470 136 478 138
rect 470 132 472 136
rect 476 132 478 136
rect 470 130 478 132
rect 480 136 488 138
rect 528 136 536 138
rect 542 139 550 141
rect 480 132 482 136
rect 486 132 488 136
rect 542 135 544 139
rect 548 135 550 139
rect 480 130 488 132
rect 528 132 536 134
rect 542 133 550 135
rect 552 139 560 141
rect 580 140 588 142
rect 552 135 554 139
rect 558 135 560 139
rect 552 133 560 135
rect 564 137 572 139
rect 564 133 566 137
rect 570 133 572 137
rect 580 136 582 140
rect 586 136 588 140
rect 580 134 588 136
rect 590 140 598 142
rect 590 136 592 140
rect 596 136 598 140
rect 590 134 598 136
rect 528 128 530 132
rect 534 128 536 132
rect 564 131 572 133
rect 64 126 72 128
rect 112 126 120 128
rect 4 124 12 126
rect 34 122 42 124
rect 4 120 12 122
rect 4 116 6 120
rect 10 116 12 120
rect 34 118 36 122
rect 40 118 42 122
rect 34 116 42 118
rect 44 122 52 124
rect 44 118 46 122
rect 50 118 52 122
rect 44 116 52 118
rect 64 122 72 124
rect 64 118 66 122
rect 70 118 72 122
rect 112 122 114 126
rect 118 122 120 126
rect 112 120 120 122
rect 122 126 130 128
rect 122 122 124 126
rect 128 122 130 126
rect 122 120 130 122
rect 132 126 140 128
rect 132 122 134 126
rect 138 122 140 126
rect 132 120 140 122
rect 142 126 150 128
rect 142 122 144 126
rect 148 122 150 126
rect 142 120 150 122
rect 152 126 160 128
rect 152 122 154 126
rect 158 122 160 126
rect 152 120 160 122
rect 162 126 170 128
rect 162 122 164 126
rect 168 122 170 126
rect 162 120 170 122
rect 172 126 180 128
rect 172 122 174 126
rect 178 122 180 126
rect 172 120 180 122
rect 182 126 190 128
rect 182 122 184 126
rect 188 122 190 126
rect 182 120 190 122
rect 192 126 200 128
rect 192 122 194 126
rect 198 122 200 126
rect 192 120 200 122
rect 202 126 210 128
rect 202 122 204 126
rect 208 122 210 126
rect 202 120 210 122
rect 212 126 220 128
rect 212 122 214 126
rect 218 122 220 126
rect 212 120 220 122
rect 222 126 230 128
rect 222 122 224 126
rect 228 122 230 126
rect 222 120 230 122
rect 232 126 240 128
rect 232 122 234 126
rect 238 122 240 126
rect 232 120 240 122
rect 296 126 304 128
rect 296 122 298 126
rect 302 122 304 126
rect 296 120 304 122
rect 360 126 368 128
rect 360 122 362 126
rect 366 122 368 126
rect 360 120 368 122
rect 370 126 378 128
rect 370 122 372 126
rect 376 122 378 126
rect 370 120 378 122
rect 380 126 388 128
rect 380 122 382 126
rect 386 122 388 126
rect 380 120 388 122
rect 390 126 398 128
rect 390 122 392 126
rect 396 122 398 126
rect 390 120 398 122
rect 400 126 408 128
rect 400 122 402 126
rect 406 122 408 126
rect 400 120 408 122
rect 410 126 418 128
rect 410 122 412 126
rect 416 122 418 126
rect 410 120 418 122
rect 420 126 428 128
rect 420 122 422 126
rect 426 122 428 126
rect 420 120 428 122
rect 430 126 438 128
rect 430 122 432 126
rect 436 122 438 126
rect 430 120 438 122
rect 440 126 448 128
rect 440 122 442 126
rect 446 122 448 126
rect 440 120 448 122
rect 450 126 458 128
rect 450 122 452 126
rect 456 122 458 126
rect 450 120 458 122
rect 460 126 468 128
rect 460 122 462 126
rect 466 122 468 126
rect 460 120 468 122
rect 470 126 478 128
rect 470 122 472 126
rect 476 122 478 126
rect 470 120 478 122
rect 480 126 488 128
rect 528 126 536 128
rect 542 129 550 131
rect 480 122 482 126
rect 486 122 488 126
rect 542 125 544 129
rect 548 125 550 129
rect 480 120 488 122
rect 528 122 536 124
rect 542 123 550 125
rect 552 129 560 131
rect 580 130 588 132
rect 552 125 554 129
rect 558 125 560 129
rect 552 123 560 125
rect 564 127 572 129
rect 564 123 566 127
rect 570 123 572 127
rect 580 126 582 130
rect 586 126 588 130
rect 580 124 588 126
rect 590 130 598 132
rect 590 126 592 130
rect 596 126 598 130
rect 590 124 598 126
rect 528 118 530 122
rect 534 118 536 122
rect 564 121 572 123
rect 64 116 72 118
rect 296 116 304 118
rect 528 116 536 118
rect 542 119 550 121
rect 4 114 12 116
rect 34 112 42 114
rect 4 110 12 112
rect 4 106 6 110
rect 10 106 12 110
rect 34 108 36 112
rect 40 108 42 112
rect 34 106 42 108
rect 44 112 52 114
rect 44 108 46 112
rect 50 108 52 112
rect 44 106 52 108
rect 64 112 72 114
rect 64 108 66 112
rect 70 108 72 112
rect 296 112 298 116
rect 302 112 304 116
rect 542 115 544 119
rect 548 115 550 119
rect 296 110 304 112
rect 528 112 536 114
rect 542 113 550 115
rect 552 119 560 121
rect 580 120 588 122
rect 552 115 554 119
rect 558 115 560 119
rect 552 113 560 115
rect 564 117 572 119
rect 564 113 566 117
rect 570 113 572 117
rect 580 116 582 120
rect 586 116 588 120
rect 580 114 588 116
rect 590 120 598 122
rect 590 116 592 120
rect 596 116 598 120
rect 590 114 598 116
rect 64 106 72 108
rect 528 108 530 112
rect 534 108 536 112
rect 564 111 572 113
rect 528 106 536 108
rect 542 109 550 111
rect 4 104 12 106
rect 542 105 544 109
rect 548 105 550 109
rect 34 102 42 104
rect 4 100 12 102
rect 4 96 6 100
rect 10 96 12 100
rect 34 98 36 102
rect 40 98 42 102
rect 34 96 42 98
rect 44 102 52 104
rect 44 98 46 102
rect 50 98 52 102
rect 44 96 52 98
rect 64 102 72 104
rect 64 98 66 102
rect 70 98 72 102
rect 64 96 72 98
rect 108 100 116 102
rect 108 96 110 100
rect 114 96 116 100
rect 4 94 12 96
rect 108 94 116 96
rect 118 100 126 102
rect 118 96 120 100
rect 124 96 126 100
rect 118 94 126 96
rect 128 100 136 102
rect 128 96 130 100
rect 134 96 136 100
rect 128 94 136 96
rect 138 100 146 102
rect 138 96 140 100
rect 144 96 146 100
rect 138 94 146 96
rect 148 100 156 102
rect 148 96 150 100
rect 154 96 156 100
rect 148 94 156 96
rect 158 100 166 102
rect 158 96 160 100
rect 164 96 166 100
rect 158 94 166 96
rect 168 100 176 102
rect 168 96 170 100
rect 174 96 176 100
rect 168 94 176 96
rect 178 100 186 102
rect 178 96 180 100
rect 184 96 186 100
rect 178 94 186 96
rect 188 100 196 102
rect 188 96 190 100
rect 194 96 196 100
rect 188 94 196 96
rect 198 100 206 102
rect 198 96 200 100
rect 204 96 206 100
rect 198 94 206 96
rect 208 100 216 102
rect 208 96 210 100
rect 214 96 216 100
rect 208 94 216 96
rect 218 100 226 102
rect 218 96 220 100
rect 224 96 226 100
rect 218 94 226 96
rect 228 100 236 102
rect 228 96 230 100
rect 234 96 236 100
rect 228 94 236 96
rect 364 101 372 103
rect 364 97 366 101
rect 370 97 372 101
rect 364 95 372 97
rect 374 101 382 103
rect 374 97 376 101
rect 380 97 382 101
rect 374 95 382 97
rect 384 101 392 103
rect 384 97 386 101
rect 390 97 392 101
rect 384 95 392 97
rect 394 101 402 103
rect 394 97 396 101
rect 400 97 402 101
rect 394 95 402 97
rect 404 101 412 103
rect 404 97 406 101
rect 410 97 412 101
rect 404 95 412 97
rect 414 101 422 103
rect 414 97 416 101
rect 420 97 422 101
rect 414 95 422 97
rect 424 101 432 103
rect 424 97 426 101
rect 430 97 432 101
rect 424 95 432 97
rect 434 101 442 103
rect 434 97 436 101
rect 440 97 442 101
rect 434 95 442 97
rect 444 101 452 103
rect 444 97 446 101
rect 450 97 452 101
rect 444 95 452 97
rect 454 101 462 103
rect 454 97 456 101
rect 460 97 462 101
rect 454 95 462 97
rect 464 101 472 103
rect 464 97 466 101
rect 470 97 472 101
rect 464 95 472 97
rect 474 101 482 103
rect 474 97 476 101
rect 480 97 482 101
rect 474 95 482 97
rect 484 101 492 103
rect 484 97 486 101
rect 490 97 492 101
rect 484 95 492 97
rect 528 102 536 104
rect 542 103 550 105
rect 552 109 560 111
rect 580 110 588 112
rect 552 105 554 109
rect 558 105 560 109
rect 552 103 560 105
rect 564 107 572 109
rect 564 103 566 107
rect 570 103 572 107
rect 580 106 582 110
rect 586 106 588 110
rect 580 104 588 106
rect 590 110 598 112
rect 590 106 592 110
rect 596 106 598 110
rect 590 104 598 106
rect 528 98 530 102
rect 534 98 536 102
rect 564 101 572 103
rect 528 96 536 98
rect 542 99 550 101
rect 542 95 544 99
rect 548 95 550 99
rect 34 92 42 94
rect 4 90 12 92
rect 4 86 6 90
rect 10 86 12 90
rect 34 88 36 92
rect 40 88 42 92
rect 34 86 42 88
rect 44 92 52 94
rect 44 88 46 92
rect 50 88 52 92
rect 44 86 52 88
rect 64 92 72 94
rect 64 88 66 92
rect 70 88 72 92
rect 64 86 72 88
rect 528 92 536 94
rect 542 93 550 95
rect 552 99 560 101
rect 580 100 588 102
rect 552 95 554 99
rect 558 95 560 99
rect 552 93 560 95
rect 564 97 572 99
rect 564 93 566 97
rect 570 93 572 97
rect 580 96 582 100
rect 586 96 588 100
rect 580 94 588 96
rect 590 100 598 102
rect 590 96 592 100
rect 596 96 598 100
rect 590 94 598 96
rect 528 88 530 92
rect 534 88 536 92
rect 564 91 572 93
rect 528 86 536 88
rect 542 89 550 91
rect 4 84 12 86
rect 542 85 544 89
rect 548 85 550 89
rect 34 82 42 84
rect 4 80 12 82
rect 4 76 6 80
rect 10 76 12 80
rect 34 78 36 82
rect 40 78 42 82
rect 34 76 42 78
rect 44 82 52 84
rect 542 83 550 85
rect 552 89 560 91
rect 580 90 588 92
rect 552 85 554 89
rect 558 85 560 89
rect 552 83 560 85
rect 564 87 572 89
rect 564 83 566 87
rect 570 83 572 87
rect 580 86 582 90
rect 586 86 588 90
rect 580 84 588 86
rect 590 90 598 92
rect 590 86 592 90
rect 596 86 598 90
rect 590 84 598 86
rect 44 78 46 82
rect 50 78 52 82
rect 564 81 572 83
rect 44 76 52 78
rect 542 79 550 81
rect 4 74 12 76
rect 542 75 544 79
rect 548 75 550 79
rect 34 72 42 74
rect 4 70 12 72
rect 4 66 6 70
rect 10 66 12 70
rect 34 68 36 72
rect 40 68 42 72
rect 34 66 42 68
rect 44 72 52 74
rect 78 73 86 75
rect 44 68 46 72
rect 50 68 52 72
rect 44 66 52 68
rect 64 70 72 72
rect 64 66 66 70
rect 70 66 72 70
rect 78 69 80 73
rect 84 69 86 73
rect 78 67 86 69
rect 107 72 115 74
rect 107 68 109 72
rect 113 68 115 72
rect 107 66 115 68
rect 118 72 126 74
rect 118 68 120 72
rect 124 68 126 72
rect 118 66 126 68
rect 128 72 136 74
rect 128 68 130 72
rect 134 68 136 72
rect 128 66 136 68
rect 138 72 146 74
rect 138 68 140 72
rect 144 68 146 72
rect 138 66 146 68
rect 148 72 156 74
rect 148 68 150 72
rect 154 68 156 72
rect 148 66 156 68
rect 158 72 166 74
rect 158 68 160 72
rect 164 68 166 72
rect 158 66 166 68
rect 168 72 176 74
rect 168 68 170 72
rect 174 68 176 72
rect 168 66 176 68
rect 178 72 186 74
rect 178 68 180 72
rect 184 68 186 72
rect 178 66 186 68
rect 188 72 196 74
rect 188 68 190 72
rect 194 68 196 72
rect 188 66 196 68
rect 198 72 206 74
rect 198 68 200 72
rect 204 68 206 72
rect 198 66 206 68
rect 208 72 216 74
rect 208 68 210 72
rect 214 68 216 72
rect 208 66 216 68
rect 218 72 226 74
rect 218 68 220 72
rect 224 68 226 72
rect 218 66 226 68
rect 228 72 236 74
rect 228 68 230 72
rect 234 68 236 72
rect 228 66 236 68
rect 364 72 372 74
rect 364 68 366 72
rect 370 68 372 72
rect 364 66 372 68
rect 374 72 382 74
rect 374 68 376 72
rect 380 68 382 72
rect 374 66 382 68
rect 384 72 392 74
rect 384 68 386 72
rect 390 68 392 72
rect 384 66 392 68
rect 394 72 402 74
rect 394 68 396 72
rect 400 68 402 72
rect 394 66 402 68
rect 404 72 412 74
rect 404 68 406 72
rect 410 68 412 72
rect 404 66 412 68
rect 414 72 422 74
rect 414 68 416 72
rect 420 68 422 72
rect 414 66 422 68
rect 424 72 432 74
rect 424 68 426 72
rect 430 68 432 72
rect 424 66 432 68
rect 434 72 442 74
rect 434 68 436 72
rect 440 68 442 72
rect 434 66 442 68
rect 444 72 452 74
rect 444 68 446 72
rect 450 68 452 72
rect 444 66 452 68
rect 454 72 462 74
rect 454 68 456 72
rect 460 68 462 72
rect 454 66 462 68
rect 464 72 472 74
rect 464 68 466 72
rect 470 68 472 72
rect 464 66 472 68
rect 474 72 482 74
rect 474 68 476 72
rect 480 68 482 72
rect 474 66 482 68
rect 484 72 492 74
rect 542 73 550 75
rect 552 79 560 81
rect 580 80 588 82
rect 552 75 554 79
rect 558 75 560 79
rect 552 73 560 75
rect 564 77 572 79
rect 564 73 566 77
rect 570 73 572 77
rect 580 76 582 80
rect 586 76 588 80
rect 580 74 588 76
rect 590 80 598 82
rect 590 76 592 80
rect 596 76 598 80
rect 590 74 598 76
rect 484 68 486 72
rect 490 68 492 72
rect 484 66 492 68
rect 528 71 536 73
rect 564 71 572 73
rect 528 67 530 71
rect 534 67 536 71
rect 4 64 12 66
rect 64 64 72 66
rect 528 65 536 67
rect 542 69 550 71
rect 542 65 544 69
rect 548 65 550 69
rect 78 62 86 64
rect 4 60 12 62
rect 4 56 6 60
rect 10 56 12 60
rect 78 58 80 62
rect 84 58 86 62
rect 4 54 12 56
rect 34 56 42 58
rect 34 52 36 56
rect 40 52 42 56
rect 4 50 12 52
rect 34 50 42 52
rect 48 56 56 58
rect 48 52 50 56
rect 54 52 56 56
rect 48 50 56 52
rect 58 56 66 58
rect 58 52 60 56
rect 64 52 66 56
rect 58 50 66 52
rect 68 56 76 58
rect 78 56 86 58
rect 107 62 115 64
rect 474 62 482 64
rect 107 58 109 62
rect 113 58 115 62
rect 107 56 115 58
rect 118 60 126 62
rect 118 56 120 60
rect 124 56 126 60
rect 68 52 70 56
rect 74 52 76 56
rect 118 54 126 56
rect 128 60 136 62
rect 128 56 130 60
rect 134 56 136 60
rect 128 54 136 56
rect 138 60 146 62
rect 138 56 140 60
rect 144 56 146 60
rect 138 54 146 56
rect 148 60 156 62
rect 148 56 150 60
rect 154 56 156 60
rect 148 54 156 56
rect 158 60 166 62
rect 158 56 160 60
rect 164 56 166 60
rect 158 54 166 56
rect 168 60 176 62
rect 168 56 170 60
rect 174 56 176 60
rect 168 54 176 56
rect 178 60 186 62
rect 178 56 180 60
rect 184 56 186 60
rect 178 54 186 56
rect 188 60 196 62
rect 188 56 190 60
rect 194 56 196 60
rect 188 54 196 56
rect 198 60 206 62
rect 198 56 200 60
rect 204 56 206 60
rect 198 54 206 56
rect 208 60 216 62
rect 208 56 210 60
rect 214 56 216 60
rect 208 54 216 56
rect 218 60 226 62
rect 218 56 220 60
rect 224 56 226 60
rect 218 54 226 56
rect 228 60 236 62
rect 228 56 230 60
rect 234 56 236 60
rect 228 54 236 56
rect 364 60 372 62
rect 364 56 366 60
rect 370 56 372 60
rect 364 54 372 56
rect 374 60 382 62
rect 374 56 376 60
rect 380 56 382 60
rect 374 54 382 56
rect 384 60 392 62
rect 384 56 386 60
rect 390 56 392 60
rect 384 54 392 56
rect 394 60 402 62
rect 394 56 396 60
rect 400 56 402 60
rect 394 54 402 56
rect 404 60 412 62
rect 404 56 406 60
rect 410 56 412 60
rect 404 54 412 56
rect 414 60 422 62
rect 414 56 416 60
rect 420 56 422 60
rect 414 54 422 56
rect 424 60 432 62
rect 424 56 426 60
rect 430 56 432 60
rect 424 54 432 56
rect 434 60 442 62
rect 434 56 436 60
rect 440 56 442 60
rect 434 54 442 56
rect 444 60 452 62
rect 444 56 446 60
rect 450 56 452 60
rect 444 54 452 56
rect 454 60 462 62
rect 454 56 456 60
rect 460 56 462 60
rect 454 54 462 56
rect 464 60 472 62
rect 464 56 466 60
rect 470 56 472 60
rect 474 58 476 62
rect 480 58 482 62
rect 474 56 482 58
rect 484 62 492 64
rect 542 63 550 65
rect 552 69 560 71
rect 580 70 588 72
rect 552 65 554 69
rect 558 65 560 69
rect 552 63 560 65
rect 564 67 572 69
rect 564 63 566 67
rect 570 63 572 67
rect 580 66 582 70
rect 586 66 588 70
rect 580 64 588 66
rect 590 70 598 72
rect 590 66 592 70
rect 596 66 598 70
rect 590 64 598 66
rect 484 58 486 62
rect 490 58 492 62
rect 564 61 572 63
rect 580 60 588 62
rect 484 56 492 58
rect 526 56 534 58
rect 464 54 472 56
rect 68 50 76 52
rect 78 52 86 54
rect 4 46 6 50
rect 10 46 12 50
rect 78 48 80 52
rect 84 48 86 52
rect 4 44 12 46
rect 34 46 42 48
rect 34 42 36 46
rect 40 42 42 46
rect 4 40 12 42
rect 34 40 42 42
rect 48 46 56 48
rect 48 42 50 46
rect 54 42 56 46
rect 48 40 56 42
rect 58 46 66 48
rect 58 42 60 46
rect 64 42 66 46
rect 58 40 66 42
rect 68 46 76 48
rect 78 46 86 48
rect 107 52 115 54
rect 474 52 482 54
rect 107 48 109 52
rect 113 48 115 52
rect 107 46 115 48
rect 118 50 126 52
rect 118 46 120 50
rect 124 46 126 50
rect 68 42 70 46
rect 74 42 76 46
rect 118 44 126 46
rect 128 50 136 52
rect 128 46 130 50
rect 134 46 136 50
rect 128 44 136 46
rect 138 50 146 52
rect 138 46 140 50
rect 144 46 146 50
rect 138 44 146 46
rect 148 50 156 52
rect 148 46 150 50
rect 154 46 156 50
rect 148 44 156 46
rect 158 50 166 52
rect 158 46 160 50
rect 164 46 166 50
rect 158 44 166 46
rect 168 50 176 52
rect 168 46 170 50
rect 174 46 176 50
rect 168 44 176 46
rect 178 50 186 52
rect 178 46 180 50
rect 184 46 186 50
rect 178 44 186 46
rect 188 50 196 52
rect 188 46 190 50
rect 194 46 196 50
rect 188 44 196 46
rect 198 50 206 52
rect 198 46 200 50
rect 204 46 206 50
rect 198 44 206 46
rect 208 50 216 52
rect 208 46 210 50
rect 214 46 216 50
rect 208 44 216 46
rect 218 50 226 52
rect 218 46 220 50
rect 224 46 226 50
rect 218 44 226 46
rect 228 50 236 52
rect 228 46 230 50
rect 234 46 236 50
rect 228 44 236 46
rect 364 50 372 52
rect 364 46 366 50
rect 370 46 372 50
rect 364 44 372 46
rect 374 50 382 52
rect 374 46 376 50
rect 380 46 382 50
rect 374 44 382 46
rect 384 50 392 52
rect 384 46 386 50
rect 390 46 392 50
rect 384 44 392 46
rect 394 50 402 52
rect 394 46 396 50
rect 400 46 402 50
rect 394 44 402 46
rect 404 50 412 52
rect 404 46 406 50
rect 410 46 412 50
rect 404 44 412 46
rect 414 50 422 52
rect 414 46 416 50
rect 420 46 422 50
rect 414 44 422 46
rect 424 50 432 52
rect 424 46 426 50
rect 430 46 432 50
rect 424 44 432 46
rect 434 50 442 52
rect 434 46 436 50
rect 440 46 442 50
rect 434 44 442 46
rect 444 50 452 52
rect 444 46 446 50
rect 450 46 452 50
rect 444 44 452 46
rect 454 50 462 52
rect 454 46 456 50
rect 460 46 462 50
rect 454 44 462 46
rect 464 50 472 52
rect 464 46 466 50
rect 470 46 472 50
rect 474 48 476 52
rect 480 48 482 52
rect 474 46 482 48
rect 484 52 492 54
rect 484 48 486 52
rect 490 48 492 52
rect 526 52 528 56
rect 532 52 534 56
rect 526 50 534 52
rect 536 56 544 58
rect 536 52 538 56
rect 542 52 544 56
rect 536 50 544 52
rect 552 56 560 58
rect 552 52 554 56
rect 558 52 560 56
rect 552 50 560 52
rect 564 57 572 59
rect 564 53 566 57
rect 570 53 572 57
rect 580 56 582 60
rect 586 56 588 60
rect 580 54 588 56
rect 590 60 598 62
rect 590 56 592 60
rect 596 56 598 60
rect 590 54 598 56
rect 564 51 572 53
rect 580 50 588 52
rect 484 46 492 48
rect 536 46 544 48
rect 464 44 472 46
rect 68 40 76 42
rect 78 42 86 44
rect 4 36 6 40
rect 10 36 12 40
rect 78 38 80 42
rect 84 38 86 42
rect 4 34 12 36
rect 48 36 56 38
rect 48 32 50 36
rect 54 32 56 36
rect 4 30 12 32
rect 48 30 56 32
rect 58 36 66 38
rect 58 32 60 36
rect 64 32 66 36
rect 58 30 66 32
rect 68 36 76 38
rect 78 36 86 38
rect 107 42 115 44
rect 474 42 482 44
rect 107 38 109 42
rect 113 38 115 42
rect 107 36 115 38
rect 118 40 126 42
rect 118 36 120 40
rect 124 36 126 40
rect 68 32 70 36
rect 74 32 76 36
rect 118 34 126 36
rect 128 40 136 42
rect 128 36 130 40
rect 134 36 136 40
rect 128 34 136 36
rect 138 40 146 42
rect 138 36 140 40
rect 144 36 146 40
rect 138 34 146 36
rect 148 40 156 42
rect 148 36 150 40
rect 154 36 156 40
rect 148 34 156 36
rect 158 40 166 42
rect 158 36 160 40
rect 164 36 166 40
rect 158 34 166 36
rect 168 40 176 42
rect 168 36 170 40
rect 174 36 176 40
rect 168 34 176 36
rect 178 40 186 42
rect 178 36 180 40
rect 184 36 186 40
rect 178 34 186 36
rect 188 40 196 42
rect 188 36 190 40
rect 194 36 196 40
rect 188 34 196 36
rect 198 40 206 42
rect 198 36 200 40
rect 204 36 206 40
rect 198 34 206 36
rect 208 40 216 42
rect 208 36 210 40
rect 214 36 216 40
rect 208 34 216 36
rect 218 40 226 42
rect 218 36 220 40
rect 224 36 226 40
rect 218 34 226 36
rect 228 40 236 42
rect 228 36 230 40
rect 234 36 236 40
rect 364 40 372 42
rect 228 34 236 36
rect 256 36 264 38
rect 68 30 76 32
rect 256 32 258 36
rect 262 32 264 36
rect 256 30 264 32
rect 266 36 274 38
rect 266 32 268 36
rect 272 32 274 36
rect 266 30 274 32
rect 276 36 284 38
rect 276 32 278 36
rect 282 32 284 36
rect 276 30 284 32
rect 286 36 294 38
rect 286 32 288 36
rect 292 32 294 36
rect 286 30 294 32
rect 296 36 304 38
rect 296 32 298 36
rect 302 32 304 36
rect 296 30 304 32
rect 306 36 314 38
rect 306 32 308 36
rect 312 32 314 36
rect 306 30 314 32
rect 316 36 324 38
rect 316 32 318 36
rect 322 32 324 36
rect 316 30 324 32
rect 326 36 334 38
rect 326 32 328 36
rect 332 32 334 36
rect 326 30 334 32
rect 336 36 344 38
rect 336 32 338 36
rect 342 32 344 36
rect 364 36 366 40
rect 370 36 372 40
rect 364 34 372 36
rect 374 40 382 42
rect 374 36 376 40
rect 380 36 382 40
rect 374 34 382 36
rect 384 40 392 42
rect 384 36 386 40
rect 390 36 392 40
rect 384 34 392 36
rect 394 40 402 42
rect 394 36 396 40
rect 400 36 402 40
rect 394 34 402 36
rect 404 40 412 42
rect 404 36 406 40
rect 410 36 412 40
rect 404 34 412 36
rect 414 40 422 42
rect 414 36 416 40
rect 420 36 422 40
rect 414 34 422 36
rect 424 40 432 42
rect 424 36 426 40
rect 430 36 432 40
rect 424 34 432 36
rect 434 40 442 42
rect 434 36 436 40
rect 440 36 442 40
rect 434 34 442 36
rect 444 40 452 42
rect 444 36 446 40
rect 450 36 452 40
rect 444 34 452 36
rect 454 40 462 42
rect 454 36 456 40
rect 460 36 462 40
rect 454 34 462 36
rect 464 40 472 42
rect 464 36 466 40
rect 470 36 472 40
rect 474 38 476 42
rect 480 38 482 42
rect 474 36 482 38
rect 484 42 492 44
rect 484 38 486 42
rect 490 38 492 42
rect 536 42 538 46
rect 542 42 544 46
rect 536 40 544 42
rect 552 46 560 48
rect 552 42 554 46
rect 558 42 560 46
rect 552 40 560 42
rect 564 47 572 49
rect 564 43 566 47
rect 570 43 572 47
rect 580 46 582 50
rect 586 46 588 50
rect 580 44 588 46
rect 590 50 598 52
rect 590 46 592 50
rect 596 46 598 50
rect 590 44 598 46
rect 564 41 572 43
rect 580 40 588 42
rect 484 36 492 38
rect 526 38 534 40
rect 464 34 472 36
rect 526 34 528 38
rect 532 34 534 38
rect 526 32 534 34
rect 552 36 560 38
rect 552 32 554 36
rect 558 32 560 36
rect 336 30 344 32
rect 552 30 560 32
rect 564 37 572 39
rect 564 33 566 37
rect 570 33 572 37
rect 580 36 582 40
rect 586 36 588 40
rect 580 34 588 36
rect 590 40 598 42
rect 590 36 592 40
rect 596 36 598 40
rect 590 34 598 36
rect 564 31 572 33
rect 580 30 588 32
rect 4 26 6 30
rect 10 26 12 30
rect 580 26 582 30
rect 586 26 588 30
rect 4 24 12 26
rect 22 24 30 26
rect 4 20 12 22
rect 4 16 6 20
rect 10 16 12 20
rect 22 20 24 24
rect 28 20 30 24
rect 22 18 30 20
rect 32 24 40 26
rect 32 20 34 24
rect 38 20 40 24
rect 32 18 40 20
rect 88 24 96 26
rect 88 20 90 24
rect 94 20 96 24
rect 88 18 96 20
rect 98 24 106 26
rect 98 20 100 24
rect 104 20 106 24
rect 98 18 106 20
rect 488 24 496 26
rect 488 20 490 24
rect 494 20 496 24
rect 488 18 496 20
rect 498 24 506 26
rect 498 20 500 24
rect 504 20 506 24
rect 498 18 506 20
rect 514 24 522 26
rect 514 20 516 24
rect 520 20 522 24
rect 514 18 522 20
rect 524 24 532 26
rect 580 24 588 26
rect 590 30 598 32
rect 590 26 592 30
rect 596 26 598 30
rect 590 24 598 26
rect 524 20 526 24
rect 530 20 532 24
rect 524 18 532 20
rect 580 20 588 22
rect 4 14 12 16
rect 580 16 582 20
rect 586 16 588 20
rect 580 14 588 16
rect 590 20 598 22
rect 590 16 592 20
rect 596 16 598 20
rect 590 14 598 16
rect 4 10 12 12
rect 56 10 64 12
rect 4 6 6 10
rect 10 6 12 10
rect 4 4 12 6
rect 14 8 22 10
rect 14 4 16 8
rect 20 4 22 8
rect 14 2 22 4
rect 24 8 32 10
rect 24 4 26 8
rect 30 4 32 8
rect 24 2 32 4
rect 34 8 42 10
rect 34 4 36 8
rect 40 4 42 8
rect 34 2 42 4
rect 46 8 54 10
rect 46 4 48 8
rect 52 4 54 8
rect 56 6 58 10
rect 62 6 64 10
rect 56 4 64 6
rect 66 10 74 12
rect 116 10 124 12
rect 66 6 68 10
rect 72 6 74 10
rect 66 4 74 6
rect 76 8 84 10
rect 76 4 78 8
rect 82 4 84 8
rect 46 2 54 4
rect 76 2 84 4
rect 86 8 94 10
rect 86 4 88 8
rect 92 4 94 8
rect 86 2 94 4
rect 96 8 104 10
rect 96 4 98 8
rect 102 4 104 8
rect 96 2 104 4
rect 106 8 114 10
rect 106 4 108 8
rect 112 4 114 8
rect 116 6 118 10
rect 122 6 124 10
rect 116 4 124 6
rect 126 10 134 12
rect 126 6 128 10
rect 132 6 134 10
rect 126 4 134 6
rect 136 10 144 12
rect 136 6 138 10
rect 142 6 144 10
rect 136 4 144 6
rect 146 10 154 12
rect 146 6 148 10
rect 152 6 154 10
rect 146 4 154 6
rect 156 10 164 12
rect 156 6 158 10
rect 162 6 164 10
rect 156 4 164 6
rect 166 10 174 12
rect 166 6 168 10
rect 172 6 174 10
rect 166 4 174 6
rect 176 10 184 12
rect 176 6 178 10
rect 182 6 184 10
rect 176 4 184 6
rect 186 10 194 12
rect 186 6 188 10
rect 192 6 194 10
rect 186 4 194 6
rect 196 10 204 12
rect 196 6 198 10
rect 202 6 204 10
rect 196 4 204 6
rect 206 10 214 12
rect 206 6 208 10
rect 212 6 214 10
rect 206 4 214 6
rect 216 10 224 12
rect 216 6 218 10
rect 222 6 224 10
rect 216 4 224 6
rect 226 10 234 12
rect 226 6 228 10
rect 232 6 234 10
rect 226 4 234 6
rect 236 10 244 12
rect 236 6 238 10
rect 242 6 244 10
rect 236 4 244 6
rect 246 10 254 12
rect 246 6 248 10
rect 252 6 254 10
rect 246 4 254 6
rect 256 10 264 12
rect 256 6 258 10
rect 262 6 264 10
rect 256 4 264 6
rect 266 10 274 12
rect 266 6 268 10
rect 272 6 274 10
rect 266 4 274 6
rect 276 10 284 12
rect 276 6 278 10
rect 282 6 284 10
rect 276 4 284 6
rect 286 10 294 12
rect 286 6 288 10
rect 292 6 294 10
rect 286 4 294 6
rect 296 10 304 12
rect 296 6 298 10
rect 302 6 304 10
rect 296 4 304 6
rect 306 10 314 12
rect 306 6 308 10
rect 312 6 314 10
rect 306 4 314 6
rect 316 10 324 12
rect 316 6 318 10
rect 322 6 324 10
rect 316 4 324 6
rect 326 10 334 12
rect 326 6 328 10
rect 332 6 334 10
rect 326 4 334 6
rect 338 10 346 12
rect 338 6 340 10
rect 344 6 346 10
rect 338 4 346 6
rect 348 10 356 12
rect 348 6 350 10
rect 354 6 356 10
rect 348 4 356 6
rect 358 10 366 12
rect 358 6 360 10
rect 364 6 366 10
rect 358 4 366 6
rect 368 10 376 12
rect 368 6 370 10
rect 374 6 376 10
rect 368 4 376 6
rect 378 10 386 12
rect 378 6 380 10
rect 384 6 386 10
rect 378 4 386 6
rect 388 10 396 12
rect 388 6 390 10
rect 394 6 396 10
rect 388 4 396 6
rect 398 10 406 12
rect 398 6 400 10
rect 404 6 406 10
rect 398 4 406 6
rect 408 10 416 12
rect 408 6 410 10
rect 414 6 416 10
rect 408 4 416 6
rect 418 10 426 12
rect 418 6 420 10
rect 424 6 426 10
rect 418 4 426 6
rect 428 10 436 12
rect 428 6 430 10
rect 434 6 436 10
rect 428 4 436 6
rect 438 10 446 12
rect 438 6 440 10
rect 444 6 446 10
rect 438 4 446 6
rect 448 10 456 12
rect 448 6 450 10
rect 454 6 456 10
rect 448 4 456 6
rect 458 10 466 12
rect 458 6 460 10
rect 464 6 466 10
rect 458 4 466 6
rect 468 10 476 12
rect 538 10 546 12
rect 468 6 470 10
rect 474 6 476 10
rect 468 4 476 6
rect 478 8 486 10
rect 478 4 480 8
rect 484 4 486 8
rect 106 2 114 4
rect 478 2 486 4
rect 488 8 496 10
rect 488 4 490 8
rect 494 4 496 8
rect 488 2 496 4
rect 498 8 506 10
rect 498 4 500 8
rect 504 4 506 8
rect 498 2 506 4
rect 508 8 516 10
rect 508 4 510 8
rect 514 4 516 8
rect 508 2 516 4
rect 518 8 526 10
rect 518 4 520 8
rect 524 4 526 8
rect 518 2 526 4
rect 528 8 536 10
rect 528 4 530 8
rect 534 4 536 8
rect 538 6 540 10
rect 544 6 546 10
rect 538 4 546 6
rect 548 10 556 12
rect 548 6 550 10
rect 554 6 556 10
rect 548 4 556 6
rect 558 10 566 12
rect 558 6 560 10
rect 564 6 566 10
rect 558 4 566 6
rect 568 10 576 12
rect 568 6 570 10
rect 574 6 576 10
rect 568 4 576 6
rect 578 10 586 12
rect 578 6 580 10
rect 584 6 586 10
rect 578 4 586 6
rect 590 10 598 12
rect 590 6 592 10
rect 596 6 598 10
rect 590 4 598 6
rect 528 2 536 4
<< genericcontact >>
rect 4 1328 8 1332
rect 16 1328 20 1332
rect 26 1328 30 1332
rect 36 1328 40 1332
rect 46 1328 50 1332
rect 56 1328 60 1332
rect 66 1328 70 1332
rect 76 1328 80 1332
rect 86 1328 90 1332
rect 96 1328 100 1332
rect 106 1328 110 1332
rect 116 1328 120 1332
rect 126 1328 130 1332
rect 136 1328 140 1332
rect 146 1328 150 1332
rect 156 1328 160 1332
rect 166 1328 170 1332
rect 176 1328 180 1332
rect 186 1328 190 1332
rect 196 1328 200 1332
rect 206 1328 210 1332
rect 216 1328 220 1332
rect 226 1328 230 1332
rect 370 1328 374 1332
rect 380 1328 384 1332
rect 390 1328 394 1332
rect 400 1328 404 1332
rect 410 1328 414 1332
rect 420 1328 424 1332
rect 430 1328 434 1332
rect 440 1328 444 1332
rect 450 1328 454 1332
rect 460 1328 464 1332
rect 470 1328 474 1332
rect 480 1328 484 1332
rect 490 1328 494 1332
rect 500 1328 504 1332
rect 510 1328 514 1332
rect 520 1328 524 1332
rect 530 1328 534 1332
rect 540 1328 544 1332
rect 550 1328 554 1332
rect 560 1328 564 1332
rect 570 1328 574 1332
rect 582 1326 586 1330
rect 592 1326 596 1330
rect 4 1318 8 1322
rect 16 1318 20 1322
rect 26 1318 30 1322
rect 36 1318 40 1322
rect 46 1318 50 1322
rect 56 1318 60 1322
rect 66 1318 70 1322
rect 76 1318 80 1322
rect 86 1318 90 1322
rect 96 1318 100 1322
rect 106 1318 110 1322
rect 116 1318 120 1322
rect 126 1318 130 1322
rect 136 1318 140 1322
rect 146 1318 150 1322
rect 156 1318 160 1322
rect 166 1318 170 1322
rect 176 1318 180 1322
rect 186 1318 190 1322
rect 196 1318 200 1322
rect 206 1318 210 1322
rect 216 1318 220 1322
rect 226 1318 230 1322
rect 370 1318 374 1322
rect 380 1318 384 1322
rect 390 1318 394 1322
rect 400 1318 404 1322
rect 410 1318 414 1322
rect 420 1318 424 1322
rect 430 1318 434 1322
rect 440 1318 444 1322
rect 450 1318 454 1322
rect 460 1318 464 1322
rect 470 1318 474 1322
rect 480 1318 484 1322
rect 490 1318 494 1322
rect 500 1318 504 1322
rect 510 1318 514 1322
rect 520 1318 524 1322
rect 530 1318 534 1322
rect 540 1318 544 1322
rect 550 1318 554 1322
rect 560 1318 564 1322
rect 570 1318 574 1322
rect 582 1316 586 1320
rect 592 1316 596 1320
rect 4 1308 8 1312
rect 14 1308 18 1312
rect 582 1306 586 1310
rect 592 1306 596 1310
rect 4 1298 8 1302
rect 14 1298 18 1302
rect 582 1296 586 1300
rect 592 1296 596 1300
rect 4 1288 8 1292
rect 14 1288 18 1292
rect 298 1288 302 1292
rect 92 1284 96 1288
rect 102 1284 106 1288
rect 114 1284 118 1288
rect 134 1284 138 1288
rect 144 1284 148 1288
rect 164 1284 168 1288
rect 174 1284 178 1288
rect 194 1284 198 1288
rect 204 1284 208 1288
rect 224 1284 228 1288
rect 368 1284 372 1288
rect 388 1284 392 1288
rect 398 1284 402 1288
rect 418 1284 422 1288
rect 428 1284 432 1288
rect 448 1284 452 1288
rect 458 1284 462 1288
rect 478 1284 482 1288
rect 490 1284 494 1288
rect 500 1284 504 1288
rect 582 1286 586 1290
rect 592 1286 596 1290
rect 4 1278 8 1282
rect 14 1278 18 1282
rect 42 1274 46 1278
rect 52 1274 56 1278
rect 92 1274 96 1278
rect 102 1274 106 1278
rect 114 1274 118 1278
rect 134 1274 138 1278
rect 144 1274 148 1278
rect 164 1274 168 1278
rect 174 1274 178 1278
rect 194 1274 198 1278
rect 204 1274 208 1278
rect 224 1274 228 1278
rect 368 1274 372 1278
rect 388 1274 392 1278
rect 398 1274 402 1278
rect 418 1274 422 1278
rect 428 1274 432 1278
rect 448 1274 452 1278
rect 458 1274 462 1278
rect 478 1274 482 1278
rect 490 1274 494 1278
rect 500 1274 504 1278
rect 544 1274 548 1278
rect 554 1274 558 1278
rect 582 1276 586 1280
rect 592 1276 596 1280
rect 4 1268 8 1272
rect 14 1268 18 1272
rect 298 1268 302 1272
rect 42 1264 46 1268
rect 52 1264 56 1268
rect 92 1264 96 1268
rect 102 1264 106 1268
rect 114 1264 118 1268
rect 134 1264 138 1268
rect 144 1264 148 1268
rect 164 1264 168 1268
rect 174 1264 178 1268
rect 194 1264 198 1268
rect 204 1264 208 1268
rect 224 1264 228 1268
rect 368 1264 372 1268
rect 388 1264 392 1268
rect 398 1264 402 1268
rect 418 1264 422 1268
rect 428 1264 432 1268
rect 448 1264 452 1268
rect 458 1264 462 1268
rect 478 1264 482 1268
rect 490 1264 494 1268
rect 500 1264 504 1268
rect 544 1264 548 1268
rect 554 1264 558 1268
rect 582 1266 586 1270
rect 592 1266 596 1270
rect 4 1258 8 1262
rect 14 1258 18 1262
rect 298 1258 302 1262
rect 42 1254 46 1258
rect 52 1254 56 1258
rect 544 1254 548 1258
rect 554 1254 558 1258
rect 582 1256 586 1260
rect 592 1256 596 1260
rect 4 1248 8 1252
rect 14 1248 18 1252
rect 298 1248 302 1252
rect 582 1246 586 1250
rect 592 1246 596 1250
rect 4 1238 8 1242
rect 14 1238 18 1242
rect 42 1234 46 1238
rect 52 1234 56 1238
rect 544 1234 548 1238
rect 554 1234 558 1238
rect 582 1236 586 1240
rect 592 1236 596 1240
rect 4 1228 8 1232
rect 14 1228 18 1232
rect 298 1228 302 1232
rect 42 1224 46 1228
rect 52 1224 56 1228
rect 66 1222 70 1226
rect 544 1224 548 1228
rect 554 1224 558 1228
rect 582 1226 586 1230
rect 592 1226 596 1230
rect 4 1218 8 1222
rect 14 1218 18 1222
rect 298 1218 302 1222
rect 530 1219 534 1223
rect 42 1214 46 1218
rect 52 1214 56 1218
rect 66 1212 70 1216
rect 544 1214 548 1218
rect 554 1214 558 1218
rect 582 1216 586 1220
rect 592 1216 596 1220
rect 4 1208 8 1212
rect 14 1208 18 1212
rect 114 1210 118 1214
rect 124 1210 128 1214
rect 134 1210 138 1214
rect 144 1210 148 1214
rect 154 1210 158 1214
rect 164 1210 168 1214
rect 174 1210 178 1214
rect 184 1210 188 1214
rect 194 1210 198 1214
rect 204 1210 208 1214
rect 214 1210 218 1214
rect 224 1210 228 1214
rect 234 1210 238 1214
rect 298 1208 302 1212
rect 362 1210 366 1214
rect 372 1210 376 1214
rect 382 1210 386 1214
rect 392 1210 396 1214
rect 402 1210 406 1214
rect 412 1210 416 1214
rect 422 1210 426 1214
rect 432 1210 436 1214
rect 442 1210 446 1214
rect 452 1210 456 1214
rect 462 1210 466 1214
rect 472 1210 476 1214
rect 482 1210 486 1214
rect 530 1209 534 1213
rect 582 1206 586 1210
rect 592 1206 596 1210
rect 66 1202 70 1206
rect 4 1198 8 1202
rect 14 1198 18 1202
rect 114 1200 118 1204
rect 124 1200 128 1204
rect 134 1200 138 1204
rect 144 1200 148 1204
rect 154 1200 158 1204
rect 164 1200 168 1204
rect 174 1200 178 1204
rect 184 1200 188 1204
rect 194 1200 198 1204
rect 204 1200 208 1204
rect 214 1200 218 1204
rect 224 1200 228 1204
rect 234 1200 238 1204
rect 362 1200 366 1204
rect 372 1200 376 1204
rect 382 1200 386 1204
rect 392 1200 396 1204
rect 402 1200 406 1204
rect 412 1200 416 1204
rect 422 1200 426 1204
rect 432 1200 436 1204
rect 442 1200 446 1204
rect 452 1200 456 1204
rect 462 1200 466 1204
rect 472 1200 476 1204
rect 482 1200 486 1204
rect 530 1199 534 1203
rect 42 1194 46 1198
rect 52 1194 56 1198
rect 66 1192 70 1196
rect 544 1194 548 1198
rect 554 1194 558 1198
rect 582 1196 586 1200
rect 592 1196 596 1200
rect 4 1188 8 1192
rect 14 1188 18 1192
rect 298 1188 302 1192
rect 530 1189 534 1193
rect 42 1184 46 1188
rect 52 1184 56 1188
rect 544 1184 548 1188
rect 554 1184 558 1188
rect 582 1186 586 1190
rect 592 1186 596 1190
rect 4 1178 8 1182
rect 14 1178 18 1182
rect 298 1178 302 1182
rect 42 1174 46 1178
rect 52 1174 56 1178
rect 544 1174 548 1178
rect 554 1174 558 1178
rect 582 1176 586 1180
rect 592 1176 596 1180
rect 4 1168 8 1172
rect 14 1168 18 1172
rect 298 1168 302 1172
rect 582 1166 586 1170
rect 592 1166 596 1170
rect 4 1158 8 1162
rect 14 1158 18 1162
rect 42 1154 46 1158
rect 52 1154 56 1158
rect 544 1154 548 1158
rect 554 1154 558 1158
rect 582 1156 586 1160
rect 592 1156 596 1160
rect 4 1148 8 1152
rect 14 1148 18 1152
rect 42 1144 46 1148
rect 52 1144 56 1148
rect 125 1146 129 1150
rect 135 1146 139 1150
rect 155 1146 159 1150
rect 165 1146 169 1150
rect 185 1146 189 1150
rect 195 1146 199 1150
rect 215 1146 219 1150
rect 225 1146 229 1150
rect 298 1148 302 1152
rect 370 1146 374 1150
rect 380 1146 384 1150
rect 400 1146 404 1150
rect 410 1146 414 1150
rect 430 1146 434 1150
rect 440 1146 444 1150
rect 460 1146 464 1150
rect 470 1146 474 1150
rect 544 1144 548 1148
rect 554 1144 558 1148
rect 582 1146 586 1150
rect 592 1146 596 1150
rect 4 1138 8 1142
rect 14 1138 18 1142
rect 298 1138 302 1142
rect 42 1134 46 1138
rect 52 1134 56 1138
rect 125 1134 129 1138
rect 135 1134 139 1138
rect 155 1134 159 1138
rect 165 1134 169 1138
rect 185 1134 189 1138
rect 195 1134 199 1138
rect 215 1134 219 1138
rect 225 1134 229 1138
rect 370 1134 374 1138
rect 380 1134 384 1138
rect 400 1134 404 1138
rect 410 1134 414 1138
rect 430 1134 434 1138
rect 440 1134 444 1138
rect 460 1134 464 1138
rect 470 1134 474 1138
rect 544 1134 548 1138
rect 554 1134 558 1138
rect 582 1136 586 1140
rect 592 1136 596 1140
rect 4 1128 8 1132
rect 14 1128 18 1132
rect 298 1128 302 1132
rect 582 1126 586 1130
rect 592 1126 596 1130
rect 4 1118 8 1122
rect 14 1118 18 1122
rect 42 1114 46 1118
rect 52 1114 56 1118
rect 544 1114 548 1118
rect 554 1114 558 1118
rect 582 1116 586 1120
rect 592 1116 596 1120
rect 4 1108 8 1112
rect 14 1108 18 1112
rect 298 1108 302 1112
rect 42 1104 46 1108
rect 52 1104 56 1108
rect 544 1104 548 1108
rect 554 1104 558 1108
rect 582 1106 586 1110
rect 592 1106 596 1110
rect 4 1098 8 1102
rect 14 1098 18 1102
rect 298 1098 302 1102
rect 42 1094 46 1098
rect 52 1094 56 1098
rect 66 1092 70 1096
rect 530 1092 534 1096
rect 544 1094 548 1098
rect 554 1094 558 1098
rect 582 1096 586 1100
rect 592 1096 596 1100
rect 4 1088 8 1092
rect 14 1088 18 1092
rect 298 1088 302 1092
rect 582 1086 586 1090
rect 592 1086 596 1090
rect 66 1082 70 1086
rect 4 1078 8 1082
rect 14 1078 18 1082
rect 114 1081 118 1085
rect 124 1081 128 1085
rect 134 1081 138 1085
rect 144 1081 148 1085
rect 154 1081 158 1085
rect 164 1081 168 1085
rect 174 1081 178 1085
rect 184 1081 188 1085
rect 194 1081 198 1085
rect 204 1081 208 1085
rect 214 1081 218 1085
rect 224 1081 228 1085
rect 234 1081 238 1085
rect 362 1081 366 1085
rect 372 1081 376 1085
rect 382 1081 386 1085
rect 392 1081 396 1085
rect 402 1081 406 1085
rect 412 1081 416 1085
rect 422 1081 426 1085
rect 432 1081 436 1085
rect 442 1081 446 1085
rect 452 1081 456 1085
rect 462 1081 466 1085
rect 472 1081 476 1085
rect 482 1081 486 1085
rect 530 1082 534 1086
rect 42 1074 46 1078
rect 52 1074 56 1078
rect 66 1072 70 1076
rect 4 1068 8 1072
rect 14 1068 18 1072
rect 114 1071 118 1075
rect 124 1071 128 1075
rect 134 1071 138 1075
rect 144 1071 148 1075
rect 154 1071 158 1075
rect 164 1071 168 1075
rect 174 1071 178 1075
rect 184 1071 188 1075
rect 194 1071 198 1075
rect 204 1071 208 1075
rect 214 1071 218 1075
rect 224 1071 228 1075
rect 234 1071 238 1075
rect 298 1068 302 1072
rect 362 1071 366 1075
rect 372 1071 376 1075
rect 382 1071 386 1075
rect 392 1071 396 1075
rect 402 1071 406 1075
rect 412 1071 416 1075
rect 422 1071 426 1075
rect 432 1071 436 1075
rect 442 1071 446 1075
rect 452 1071 456 1075
rect 462 1071 466 1075
rect 472 1071 476 1075
rect 482 1071 486 1075
rect 530 1072 534 1076
rect 544 1074 548 1078
rect 554 1074 558 1078
rect 582 1076 586 1080
rect 592 1076 596 1080
rect 42 1064 46 1068
rect 52 1064 56 1068
rect 66 1062 70 1066
rect 530 1062 534 1066
rect 544 1064 548 1068
rect 554 1064 558 1068
rect 582 1066 586 1070
rect 592 1066 596 1070
rect 4 1058 8 1062
rect 14 1058 18 1062
rect 298 1058 302 1062
rect 42 1054 46 1058
rect 52 1054 56 1058
rect 544 1054 548 1058
rect 554 1054 558 1058
rect 582 1056 586 1060
rect 592 1056 596 1060
rect 4 1048 8 1052
rect 14 1048 18 1052
rect 298 1048 302 1052
rect 582 1046 586 1050
rect 592 1046 596 1050
rect 4 1038 8 1042
rect 14 1038 18 1042
rect 42 1034 46 1038
rect 52 1034 56 1038
rect 544 1034 548 1038
rect 554 1034 558 1038
rect 582 1036 586 1040
rect 592 1036 596 1040
rect 4 1028 8 1032
rect 14 1028 18 1032
rect 298 1028 302 1032
rect 42 1024 46 1028
rect 52 1024 56 1028
rect 544 1024 548 1028
rect 554 1024 558 1028
rect 582 1026 586 1030
rect 592 1026 596 1030
rect 4 1018 8 1022
rect 14 1018 18 1022
rect 124 1018 128 1022
rect 134 1018 138 1022
rect 154 1018 158 1022
rect 164 1018 168 1022
rect 184 1018 188 1022
rect 194 1018 198 1022
rect 214 1018 218 1022
rect 224 1018 228 1022
rect 298 1018 302 1022
rect 369 1018 373 1022
rect 379 1018 383 1022
rect 399 1018 403 1022
rect 409 1018 413 1022
rect 429 1018 433 1022
rect 439 1018 443 1022
rect 459 1018 463 1022
rect 469 1018 473 1022
rect 42 1014 46 1018
rect 52 1014 56 1018
rect 544 1014 548 1018
rect 554 1014 558 1018
rect 582 1016 586 1020
rect 592 1016 596 1020
rect 4 1008 8 1012
rect 14 1008 18 1012
rect 124 1006 128 1010
rect 134 1006 138 1010
rect 154 1006 158 1010
rect 164 1006 168 1010
rect 184 1006 188 1010
rect 194 1006 198 1010
rect 214 1006 218 1010
rect 224 1006 228 1010
rect 298 1008 302 1012
rect 369 1006 373 1010
rect 379 1006 383 1010
rect 399 1006 403 1010
rect 409 1006 413 1010
rect 429 1006 433 1010
rect 439 1006 443 1010
rect 459 1006 463 1010
rect 469 1006 473 1010
rect 582 1006 586 1010
rect 592 1006 596 1010
rect 4 998 8 1002
rect 14 998 18 1002
rect 42 994 46 998
rect 52 994 56 998
rect 544 994 548 998
rect 554 994 558 998
rect 582 996 586 1000
rect 592 996 596 1000
rect 4 988 8 992
rect 14 988 18 992
rect 298 988 302 992
rect 42 984 46 988
rect 52 984 56 988
rect 544 984 548 988
rect 554 984 558 988
rect 582 986 586 990
rect 592 986 596 990
rect 4 978 8 982
rect 14 978 18 982
rect 298 978 302 982
rect 42 974 46 978
rect 52 974 56 978
rect 544 974 548 978
rect 554 974 558 978
rect 582 976 586 980
rect 592 976 596 980
rect 4 968 8 972
rect 14 968 18 972
rect 298 968 302 972
rect 582 966 586 970
rect 592 966 596 970
rect 530 962 534 966
rect 4 958 8 962
rect 14 958 18 962
rect 42 954 46 958
rect 52 954 56 958
rect 66 956 70 960
rect 114 952 118 956
rect 124 952 128 956
rect 134 952 138 956
rect 144 952 148 956
rect 154 952 158 956
rect 164 952 168 956
rect 174 952 178 956
rect 184 952 188 956
rect 194 952 198 956
rect 204 952 208 956
rect 214 952 218 956
rect 224 952 228 956
rect 234 952 238 956
rect 362 952 366 956
rect 372 952 376 956
rect 382 952 386 956
rect 392 952 396 956
rect 402 952 406 956
rect 412 952 416 956
rect 422 952 426 956
rect 432 952 436 956
rect 442 952 446 956
rect 452 952 456 956
rect 462 952 466 956
rect 472 952 476 956
rect 482 952 486 956
rect 530 952 534 956
rect 544 954 548 958
rect 554 954 558 958
rect 582 956 586 960
rect 592 956 596 960
rect 4 948 8 952
rect 14 948 18 952
rect 42 944 46 948
rect 52 944 56 948
rect 66 946 70 950
rect 298 948 302 952
rect 114 942 118 946
rect 124 942 128 946
rect 134 942 138 946
rect 144 942 148 946
rect 154 942 158 946
rect 164 942 168 946
rect 174 942 178 946
rect 184 942 188 946
rect 194 942 198 946
rect 204 942 208 946
rect 214 942 218 946
rect 224 942 228 946
rect 234 942 238 946
rect 362 942 366 946
rect 372 942 376 946
rect 382 942 386 946
rect 392 942 396 946
rect 402 942 406 946
rect 412 942 416 946
rect 422 942 426 946
rect 432 942 436 946
rect 442 942 446 946
rect 452 942 456 946
rect 462 942 466 946
rect 472 942 476 946
rect 482 942 486 946
rect 530 942 534 946
rect 544 944 548 948
rect 554 944 558 948
rect 582 946 586 950
rect 592 946 596 950
rect 4 938 8 942
rect 14 938 18 942
rect 42 934 46 938
rect 52 934 56 938
rect 66 936 70 940
rect 298 938 302 942
rect 530 932 534 936
rect 544 934 548 938
rect 554 934 558 938
rect 582 936 586 940
rect 592 936 596 940
rect 4 928 8 932
rect 14 928 18 932
rect 66 926 70 930
rect 298 928 302 932
rect 582 926 586 930
rect 592 926 596 930
rect 530 922 534 926
rect 4 918 8 922
rect 14 918 18 922
rect 42 914 46 918
rect 52 914 56 918
rect 66 916 70 920
rect 530 912 534 916
rect 544 914 548 918
rect 554 914 558 918
rect 582 916 586 920
rect 592 916 596 920
rect 4 908 8 912
rect 14 908 18 912
rect 42 904 46 908
rect 52 904 56 908
rect 66 906 70 910
rect 298 908 302 912
rect 544 904 548 908
rect 554 904 558 908
rect 582 906 586 910
rect 592 906 596 910
rect 4 898 8 902
rect 14 898 18 902
rect 298 898 302 902
rect 42 894 46 898
rect 52 894 56 898
rect 544 894 548 898
rect 554 894 558 898
rect 582 896 586 900
rect 592 896 596 900
rect 4 888 8 892
rect 14 888 18 892
rect 125 888 129 892
rect 135 888 139 892
rect 155 888 159 892
rect 165 888 169 892
rect 185 888 189 892
rect 195 888 199 892
rect 215 888 219 892
rect 225 888 229 892
rect 298 888 302 892
rect 371 888 375 892
rect 381 888 385 892
rect 401 888 405 892
rect 411 888 415 892
rect 431 888 435 892
rect 441 888 445 892
rect 461 888 465 892
rect 471 888 475 892
rect 582 886 586 890
rect 592 886 596 890
rect 4 878 8 882
rect 14 878 18 882
rect 42 874 46 878
rect 52 874 56 878
rect 105 876 109 880
rect 125 876 129 880
rect 135 876 139 880
rect 155 876 159 880
rect 165 876 169 880
rect 185 876 189 880
rect 195 876 199 880
rect 215 876 219 880
rect 225 876 229 880
rect 371 876 375 880
rect 381 876 385 880
rect 401 876 405 880
rect 411 876 415 880
rect 431 876 435 880
rect 441 876 445 880
rect 461 876 465 880
rect 471 876 475 880
rect 491 876 495 880
rect 544 874 548 878
rect 554 874 558 878
rect 582 876 586 880
rect 592 876 596 880
rect 4 868 8 872
rect 14 868 18 872
rect 298 868 302 872
rect 42 864 46 868
rect 52 864 56 868
rect 95 864 99 868
rect 105 864 109 868
rect 115 864 119 868
rect 125 864 129 868
rect 135 864 139 868
rect 145 864 149 868
rect 155 864 159 868
rect 165 864 169 868
rect 175 864 179 868
rect 185 864 189 868
rect 195 864 199 868
rect 205 864 209 868
rect 215 864 219 868
rect 225 864 229 868
rect 371 864 375 868
rect 381 864 385 868
rect 391 864 395 868
rect 401 864 405 868
rect 411 864 415 868
rect 421 864 425 868
rect 431 864 435 868
rect 441 864 445 868
rect 451 864 455 868
rect 461 864 465 868
rect 471 864 475 868
rect 481 864 485 868
rect 491 864 495 868
rect 501 864 505 868
rect 544 864 548 868
rect 554 864 558 868
rect 582 866 586 870
rect 592 866 596 870
rect 4 858 8 862
rect 14 858 18 862
rect 582 856 586 860
rect 592 856 596 860
rect 4 848 8 852
rect 14 848 18 852
rect 582 846 586 850
rect 592 846 596 850
rect 4 838 8 842
rect 14 838 18 842
rect 32 833 36 837
rect 42 833 46 837
rect 52 833 56 837
rect 80 833 84 837
rect 90 833 94 837
rect 100 833 104 837
rect 110 833 114 837
rect 120 833 124 837
rect 130 833 134 837
rect 140 833 144 837
rect 150 833 154 837
rect 160 833 164 837
rect 170 833 174 837
rect 180 833 184 837
rect 190 833 194 837
rect 200 833 204 837
rect 210 833 214 837
rect 220 833 224 837
rect 298 833 302 837
rect 370 833 374 837
rect 380 833 384 837
rect 390 833 394 837
rect 400 833 404 837
rect 410 833 414 837
rect 420 833 424 837
rect 430 833 434 837
rect 440 833 444 837
rect 450 833 454 837
rect 460 833 464 837
rect 470 833 474 837
rect 480 833 484 837
rect 490 833 494 837
rect 500 833 504 837
rect 510 833 514 837
rect 520 833 524 837
rect 530 833 534 837
rect 540 833 544 837
rect 550 833 554 837
rect 560 833 564 837
rect 570 833 574 837
rect 582 836 586 840
rect 592 836 596 840
rect 4 828 8 832
rect 14 828 18 832
rect 32 823 36 827
rect 42 823 46 827
rect 52 823 56 827
rect 80 823 84 827
rect 90 823 94 827
rect 100 823 104 827
rect 110 823 114 827
rect 120 823 124 827
rect 130 823 134 827
rect 140 823 144 827
rect 150 823 154 827
rect 160 823 164 827
rect 170 823 174 827
rect 180 823 184 827
rect 190 823 194 827
rect 200 823 204 827
rect 210 823 214 827
rect 220 823 224 827
rect 298 823 302 827
rect 370 823 374 827
rect 380 823 384 827
rect 390 823 394 827
rect 400 823 404 827
rect 410 823 414 827
rect 420 823 424 827
rect 430 823 434 827
rect 440 823 444 827
rect 450 823 454 827
rect 460 823 464 827
rect 470 823 474 827
rect 480 823 484 827
rect 490 823 494 827
rect 500 823 504 827
rect 510 823 514 827
rect 520 823 524 827
rect 530 823 534 827
rect 540 823 544 827
rect 550 823 554 827
rect 560 823 564 827
rect 570 823 574 827
rect 582 826 586 830
rect 592 826 596 830
rect 4 808 8 812
rect 592 807 596 811
rect 225 803 229 807
rect 235 803 239 807
rect 245 803 249 807
rect 553 803 557 807
rect 563 803 567 807
rect 573 803 577 807
rect 4 798 8 802
rect 225 793 229 797
rect 235 793 239 797
rect 245 793 249 797
rect 389 793 393 797
rect 399 793 403 797
rect 409 793 413 797
rect 553 793 557 797
rect 563 793 567 797
rect 573 793 577 797
rect 4 788 8 792
rect 592 787 596 791
rect 389 783 393 787
rect 399 783 403 787
rect 409 783 413 787
rect 4 778 8 782
rect 52 772 56 776
rect 62 772 66 776
rect 4 768 8 772
rect 592 767 596 771
rect 4 758 8 762
rect 30 754 34 758
rect 46 754 50 758
rect 62 752 66 756
rect 80 753 84 757
rect 4 748 8 752
rect 96 750 100 754
rect 112 753 116 757
rect 128 750 132 754
rect 144 753 148 757
rect 160 750 164 754
rect 176 753 180 757
rect 208 754 212 758
rect 288 757 292 761
rect 304 758 308 762
rect 192 750 196 754
rect 224 750 228 754
rect 240 752 244 756
rect 256 750 260 754
rect 272 752 276 756
rect 388 754 392 758
rect 404 754 408 758
rect 436 754 440 758
rect 452 755 456 759
rect 468 755 472 759
rect 484 755 488 759
rect 500 755 504 759
rect 516 755 520 759
rect 532 755 536 759
rect 548 755 552 759
rect 564 755 568 759
rect 580 755 584 759
rect 30 744 34 748
rect 62 742 66 746
rect 80 743 84 747
rect 112 743 116 747
rect 144 743 148 747
rect 176 743 180 747
rect 208 744 212 748
rect 288 746 292 750
rect 304 746 308 750
rect 240 742 244 746
rect 4 738 8 742
rect 256 740 260 744
rect 272 742 276 746
rect 404 744 408 748
rect 420 742 424 746
rect 436 744 440 748
rect 468 745 472 749
rect 500 745 504 749
rect 532 745 536 749
rect 564 745 568 749
rect 592 747 596 751
rect 30 734 34 738
rect 46 734 50 738
rect 62 732 66 736
rect 80 733 84 737
rect 4 728 8 732
rect 96 730 100 734
rect 112 733 116 737
rect 128 730 132 734
rect 144 733 148 737
rect 160 730 164 734
rect 176 733 180 737
rect 208 734 212 738
rect 192 730 196 734
rect 224 730 228 734
rect 240 732 244 736
rect 256 730 260 734
rect 272 732 276 736
rect 288 734 292 738
rect 304 735 308 739
rect 388 734 392 738
rect 404 734 408 738
rect 420 732 424 736
rect 436 734 440 738
rect 452 735 456 739
rect 468 735 472 739
rect 484 735 488 739
rect 500 735 504 739
rect 516 735 520 739
rect 532 735 536 739
rect 548 735 552 739
rect 564 735 568 739
rect 580 735 584 739
rect 30 724 34 728
rect 62 722 66 726
rect 80 723 84 727
rect 112 723 116 727
rect 144 723 148 727
rect 176 723 180 727
rect 208 724 212 728
rect 4 718 8 722
rect 256 720 260 724
rect 288 722 292 726
rect 304 722 308 726
rect 404 724 408 728
rect 436 724 440 728
rect 468 725 472 729
rect 500 725 504 729
rect 532 725 536 729
rect 564 725 568 729
rect 592 727 596 731
rect 46 714 50 718
rect 62 712 66 716
rect 4 708 8 712
rect 96 710 100 714
rect 112 713 116 717
rect 128 710 132 714
rect 144 713 148 717
rect 160 710 164 714
rect 176 713 180 717
rect 208 714 212 718
rect 192 710 196 714
rect 224 710 228 714
rect 256 710 260 714
rect 272 712 276 716
rect 388 714 392 718
rect 404 714 408 718
rect 304 710 308 714
rect 420 711 424 715
rect 436 714 440 718
rect 452 715 456 719
rect 468 715 472 719
rect 484 715 488 719
rect 500 715 504 719
rect 516 715 520 719
rect 532 715 536 719
rect 548 715 552 719
rect 564 715 568 719
rect 580 715 584 719
rect 592 707 596 711
rect 4 698 8 702
rect 20 696 24 700
rect 52 696 56 700
rect 106 695 110 699
rect 116 695 120 699
rect 174 696 178 700
rect 184 696 188 700
rect 276 696 280 700
rect 286 696 290 700
rect 462 697 466 701
rect 472 697 476 701
rect 558 697 562 701
rect 568 697 572 701
rect 4 688 8 692
rect 36 688 40 692
rect 78 687 82 691
rect 92 687 96 691
rect 130 687 134 691
rect 140 687 144 691
rect 150 687 154 691
rect 160 687 164 691
rect 200 689 204 693
rect 218 689 222 693
rect 250 689 254 693
rect 390 687 394 691
rect 400 687 404 691
rect 410 687 414 691
rect 420 687 424 691
rect 448 688 452 692
rect 486 687 490 691
rect 496 687 500 691
rect 516 687 520 691
rect 544 686 548 690
rect 582 687 586 691
rect 592 687 596 691
rect 66 672 70 676
rect 76 672 80 676
rect 162 672 166 676
rect 172 672 176 676
rect 276 672 280 676
rect 286 672 290 676
rect 4 656 8 660
rect 36 657 40 661
rect 78 657 82 661
rect 92 657 96 661
rect 130 657 134 661
rect 150 657 154 661
rect 160 657 164 661
rect 198 657 202 661
rect 220 657 224 661
rect 276 657 280 661
rect 390 657 394 661
rect 400 657 404 661
rect 420 657 424 661
rect 448 657 452 661
rect 486 657 490 661
rect 496 657 500 661
rect 516 657 520 661
rect 544 657 548 661
rect 582 658 586 662
rect 592 658 596 662
rect 4 646 8 650
rect 20 649 24 653
rect 52 649 56 653
rect 106 649 110 653
rect 116 649 120 653
rect 174 649 178 653
rect 184 649 188 653
rect 250 649 254 653
rect 260 649 264 653
rect 462 649 466 653
rect 472 649 476 653
rect 558 649 562 653
rect 568 649 572 653
rect 592 648 596 652
rect 46 635 50 639
rect 62 633 66 637
rect 96 635 100 639
rect 112 633 116 637
rect 144 633 148 637
rect 176 634 180 638
rect 208 633 212 637
rect 224 635 228 639
rect 240 634 244 638
rect 272 634 276 638
rect 288 635 292 639
rect 4 626 8 630
rect 128 627 132 631
rect 160 627 164 631
rect 30 623 34 627
rect 62 623 66 627
rect 80 623 84 627
rect 112 623 116 627
rect 144 623 148 627
rect 176 624 180 628
rect 192 627 196 631
rect 208 623 212 627
rect 240 624 244 628
rect 288 625 292 629
rect 388 627 392 631
rect 404 627 408 631
rect 420 627 424 631
rect 436 627 440 631
rect 452 627 456 631
rect 468 627 472 631
rect 484 627 488 631
rect 500 627 504 631
rect 516 627 520 631
rect 532 627 536 631
rect 548 627 552 631
rect 564 627 568 631
rect 580 627 584 631
rect 592 628 596 632
rect 30 613 34 617
rect 46 615 50 619
rect 62 613 66 617
rect 80 613 84 617
rect 96 615 100 619
rect 112 613 116 617
rect 144 613 148 617
rect 176 614 180 618
rect 208 613 212 617
rect 224 615 228 619
rect 240 614 244 618
rect 256 617 260 621
rect 288 615 292 619
rect 404 617 408 621
rect 436 617 440 621
rect 468 617 472 621
rect 500 617 504 621
rect 532 617 536 621
rect 564 617 568 621
rect 304 613 308 617
rect 4 606 8 610
rect 128 607 132 611
rect 160 607 164 611
rect 30 603 34 607
rect 62 603 66 607
rect 80 603 84 607
rect 112 603 116 607
rect 144 603 148 607
rect 176 604 180 608
rect 192 607 196 611
rect 208 603 212 607
rect 240 604 244 608
rect 256 607 260 611
rect 272 608 276 612
rect 288 605 292 609
rect 388 607 392 611
rect 404 607 408 611
rect 420 607 424 611
rect 436 607 440 611
rect 452 607 456 611
rect 468 607 472 611
rect 484 607 488 611
rect 500 607 504 611
rect 516 607 520 611
rect 532 607 536 611
rect 548 607 552 611
rect 564 607 568 611
rect 580 607 584 611
rect 592 608 596 612
rect 304 603 308 607
rect 30 593 34 597
rect 46 595 50 599
rect 62 593 66 597
rect 80 593 84 597
rect 96 595 100 599
rect 112 593 116 597
rect 144 593 148 597
rect 176 594 180 598
rect 208 593 212 597
rect 224 595 228 599
rect 240 594 244 598
rect 256 597 260 601
rect 272 598 276 602
rect 288 595 292 599
rect 404 597 408 601
rect 436 597 440 601
rect 468 597 472 601
rect 500 597 504 601
rect 532 597 536 601
rect 564 597 568 601
rect 304 593 308 597
rect 4 586 8 590
rect 128 587 132 591
rect 30 583 34 587
rect 62 583 66 587
rect 80 583 84 587
rect 112 583 116 587
rect 144 583 148 587
rect 176 584 180 588
rect 192 587 196 591
rect 208 583 212 587
rect 240 584 244 588
rect 256 587 260 591
rect 272 588 276 592
rect 288 585 292 589
rect 404 587 408 591
rect 436 587 440 591
rect 468 587 472 591
rect 500 587 504 591
rect 532 587 536 591
rect 564 587 568 591
rect 580 587 584 591
rect 592 588 596 592
rect 304 583 308 587
rect 30 573 34 577
rect 46 575 50 579
rect 62 573 66 577
rect 80 573 84 577
rect 96 575 100 579
rect 160 577 164 581
rect 112 573 116 577
rect 144 573 148 577
rect 176 574 180 578
rect 208 573 212 577
rect 224 575 228 579
rect 240 574 244 578
rect 256 577 260 581
rect 272 578 276 582
rect 288 575 292 579
rect 388 577 392 581
rect 404 577 408 581
rect 420 577 424 581
rect 436 577 440 581
rect 452 577 456 581
rect 468 577 472 581
rect 484 577 488 581
rect 500 577 504 581
rect 516 577 520 581
rect 532 577 536 581
rect 548 577 552 581
rect 564 577 568 581
rect 304 573 308 577
rect 4 566 8 570
rect 128 567 132 571
rect 160 567 164 571
rect 30 563 34 567
rect 62 563 66 567
rect 80 563 84 567
rect 112 563 116 567
rect 144 563 148 567
rect 176 564 180 568
rect 192 567 196 571
rect 208 563 212 567
rect 240 564 244 568
rect 256 567 260 571
rect 272 568 276 572
rect 288 565 292 569
rect 388 567 392 571
rect 404 567 408 571
rect 420 567 424 571
rect 436 567 440 571
rect 452 567 456 571
rect 468 567 472 571
rect 484 567 488 571
rect 500 567 504 571
rect 516 567 520 571
rect 532 567 536 571
rect 548 567 552 571
rect 564 567 568 571
rect 580 567 584 571
rect 592 568 596 572
rect 304 563 308 567
rect 30 553 34 557
rect 46 555 50 559
rect 62 553 66 557
rect 80 553 84 557
rect 96 555 100 559
rect 112 553 116 557
rect 144 553 148 557
rect 176 554 180 558
rect 208 553 212 557
rect 224 555 228 559
rect 240 554 244 558
rect 256 557 260 561
rect 272 558 276 562
rect 288 555 292 559
rect 404 557 408 561
rect 436 557 440 561
rect 468 557 472 561
rect 500 557 504 561
rect 532 557 536 561
rect 564 557 568 561
rect 304 553 308 557
rect 4 546 8 550
rect 160 547 164 551
rect 30 543 34 547
rect 62 543 66 547
rect 80 543 84 547
rect 112 543 116 547
rect 144 543 148 547
rect 176 544 180 548
rect 192 547 196 551
rect 208 543 212 547
rect 240 544 244 548
rect 256 547 260 551
rect 288 545 292 549
rect 388 547 392 551
rect 404 547 408 551
rect 420 547 424 551
rect 436 547 440 551
rect 452 547 456 551
rect 468 547 472 551
rect 484 547 488 551
rect 500 547 504 551
rect 516 547 520 551
rect 532 547 536 551
rect 548 547 552 551
rect 564 547 568 551
rect 580 547 584 551
rect 592 548 596 552
rect 304 543 308 547
rect 4 526 8 530
rect 24 529 28 533
rect 34 529 38 533
rect 52 529 56 533
rect 62 529 66 533
rect 92 529 96 533
rect 102 529 106 533
rect 120 520 124 524
rect 130 520 134 524
rect 140 520 144 524
rect 150 520 154 524
rect 160 520 164 524
rect 170 520 174 524
rect 180 520 184 524
rect 190 520 194 524
rect 200 520 204 524
rect 210 520 214 524
rect 220 520 224 524
rect 388 523 392 527
rect 484 523 488 527
rect 582 525 586 529
rect 592 528 596 532
rect 36 510 40 514
rect 46 510 50 514
rect 56 510 60 514
rect 66 510 70 514
rect 6 506 10 510
rect 110 508 114 512
rect 120 508 124 512
rect 130 508 134 512
rect 140 508 144 512
rect 150 508 154 512
rect 160 508 164 512
rect 170 508 174 512
rect 180 508 184 512
rect 190 508 194 512
rect 200 508 204 512
rect 210 508 214 512
rect 220 510 224 514
rect 391 510 395 514
rect 401 510 405 514
rect 411 510 415 514
rect 421 510 425 514
rect 431 510 435 514
rect 441 510 445 514
rect 451 510 455 514
rect 482 513 486 517
rect 492 513 496 517
rect 502 513 506 517
rect 529 515 533 519
rect 542 515 546 519
rect 552 515 556 519
rect 562 515 566 519
rect 572 515 576 519
rect 582 515 586 519
rect 592 506 596 510
rect 6 496 10 500
rect 582 496 586 500
rect 592 496 596 500
rect 6 486 10 490
rect 582 486 586 490
rect 592 486 596 490
rect 6 476 10 480
rect 36 478 40 482
rect 46 478 50 482
rect 56 478 60 482
rect 66 478 70 482
rect 108 480 112 484
rect 118 480 122 484
rect 128 480 132 484
rect 138 480 142 484
rect 148 480 152 484
rect 158 480 162 484
rect 168 480 172 484
rect 178 480 182 484
rect 188 480 192 484
rect 198 480 202 484
rect 208 480 212 484
rect 218 480 222 484
rect 228 480 232 484
rect 366 480 370 484
rect 376 480 380 484
rect 386 480 390 484
rect 396 480 400 484
rect 406 480 410 484
rect 416 480 420 484
rect 426 480 430 484
rect 436 480 440 484
rect 446 480 450 484
rect 456 480 460 484
rect 466 480 470 484
rect 476 480 480 484
rect 486 480 490 484
rect 544 478 548 482
rect 554 478 558 482
rect 582 476 586 480
rect 592 476 596 480
rect 6 466 10 470
rect 36 468 40 472
rect 46 468 50 472
rect 56 468 60 472
rect 66 468 70 472
rect 108 470 112 474
rect 118 470 122 474
rect 128 470 132 474
rect 138 470 142 474
rect 148 470 152 474
rect 158 470 162 474
rect 168 470 172 474
rect 178 470 182 474
rect 188 470 192 474
rect 198 470 202 474
rect 208 470 212 474
rect 218 470 222 474
rect 228 470 232 474
rect 298 472 302 476
rect 366 470 370 474
rect 376 470 380 474
rect 386 470 390 474
rect 396 470 400 474
rect 406 470 410 474
rect 416 470 420 474
rect 426 470 430 474
rect 436 470 440 474
rect 446 470 450 474
rect 456 470 460 474
rect 466 470 470 474
rect 476 470 480 474
rect 486 470 490 474
rect 544 468 548 472
rect 554 468 558 472
rect 582 466 586 470
rect 592 466 596 470
rect 6 456 10 460
rect 36 458 40 462
rect 46 458 50 462
rect 110 460 114 464
rect 120 460 124 464
rect 140 460 144 464
rect 150 460 154 464
rect 170 460 174 464
rect 180 460 184 464
rect 200 460 204 464
rect 210 460 214 464
rect 230 460 234 464
rect 298 462 302 466
rect 366 460 370 464
rect 376 460 380 464
rect 396 460 400 464
rect 406 460 410 464
rect 426 460 430 464
rect 436 460 440 464
rect 456 460 460 464
rect 466 460 470 464
rect 486 460 490 464
rect 544 455 548 459
rect 554 455 558 459
rect 582 456 586 460
rect 592 456 596 460
rect 6 446 10 450
rect 110 448 114 452
rect 120 448 124 452
rect 140 448 144 452
rect 150 448 154 452
rect 170 448 174 452
rect 180 448 184 452
rect 200 448 204 452
rect 210 448 214 452
rect 230 448 234 452
rect 366 448 370 452
rect 376 448 380 452
rect 396 448 400 452
rect 406 448 410 452
rect 426 448 430 452
rect 436 448 440 452
rect 456 448 460 452
rect 466 448 470 452
rect 486 448 490 452
rect 582 446 586 450
rect 592 446 596 450
rect 298 442 302 446
rect 6 436 10 440
rect 36 438 40 442
rect 46 438 50 442
rect 298 432 302 436
rect 544 435 548 439
rect 554 435 558 439
rect 582 436 586 440
rect 592 436 596 440
rect 6 426 10 430
rect 36 428 40 432
rect 46 428 50 432
rect 66 428 70 432
rect 530 428 534 432
rect 544 425 548 429
rect 554 425 558 429
rect 582 426 586 430
rect 592 426 596 430
rect 6 416 10 420
rect 36 418 40 422
rect 46 418 50 422
rect 66 418 70 422
rect 530 418 534 422
rect 298 412 302 416
rect 544 415 548 419
rect 554 415 558 419
rect 582 416 586 420
rect 592 416 596 420
rect 6 406 10 410
rect 66 408 70 412
rect 530 408 534 412
rect 582 406 586 410
rect 592 406 596 410
rect 298 402 302 406
rect 6 396 10 400
rect 36 398 40 402
rect 46 398 50 402
rect 66 398 70 402
rect 530 398 534 402
rect 114 394 118 398
rect 124 394 128 398
rect 134 394 138 398
rect 144 394 148 398
rect 154 394 158 398
rect 164 394 168 398
rect 174 394 178 398
rect 184 394 188 398
rect 194 394 198 398
rect 204 394 208 398
rect 214 394 218 398
rect 224 394 228 398
rect 234 394 238 398
rect 362 394 366 398
rect 372 394 376 398
rect 382 394 386 398
rect 392 394 396 398
rect 402 394 406 398
rect 412 394 416 398
rect 422 394 426 398
rect 432 394 436 398
rect 442 394 446 398
rect 452 394 456 398
rect 462 394 466 398
rect 472 394 476 398
rect 482 394 486 398
rect 544 395 548 399
rect 554 395 558 399
rect 582 396 586 400
rect 592 396 596 400
rect 6 386 10 390
rect 36 388 40 392
rect 46 388 50 392
rect 66 388 70 392
rect 530 388 534 392
rect 114 382 118 386
rect 124 382 128 386
rect 134 382 138 386
rect 144 382 148 386
rect 154 382 158 386
rect 164 382 168 386
rect 174 382 178 386
rect 184 382 188 386
rect 194 382 198 386
rect 204 382 208 386
rect 214 382 218 386
rect 224 382 228 386
rect 234 382 238 386
rect 298 382 302 386
rect 362 382 366 386
rect 372 382 376 386
rect 382 382 386 386
rect 392 382 396 386
rect 402 382 406 386
rect 412 382 416 386
rect 422 382 426 386
rect 432 382 436 386
rect 442 382 446 386
rect 452 382 456 386
rect 462 382 466 386
rect 472 382 476 386
rect 482 382 486 386
rect 544 385 548 389
rect 554 385 558 389
rect 582 386 586 390
rect 592 386 596 390
rect 6 376 10 380
rect 36 378 40 382
rect 46 378 50 382
rect 66 378 70 382
rect 530 378 534 382
rect 298 372 302 376
rect 544 375 548 379
rect 554 375 558 379
rect 582 376 586 380
rect 592 376 596 380
rect 6 366 10 370
rect 66 368 70 372
rect 530 368 534 372
rect 582 366 586 370
rect 592 366 596 370
rect 6 356 10 360
rect 36 358 40 362
rect 46 358 50 362
rect 66 358 70 362
rect 530 358 534 362
rect 298 352 302 356
rect 544 355 548 359
rect 554 355 558 359
rect 582 356 586 360
rect 592 356 596 360
rect 6 346 10 350
rect 36 348 40 352
rect 46 348 50 352
rect 66 348 70 352
rect 530 348 534 352
rect 298 342 302 346
rect 544 345 548 349
rect 554 345 558 349
rect 582 346 586 350
rect 592 346 596 350
rect 6 336 10 340
rect 36 338 40 342
rect 46 338 50 342
rect 66 338 70 342
rect 530 338 534 342
rect 544 335 548 339
rect 554 335 558 339
rect 582 336 586 340
rect 592 336 596 340
rect 6 326 10 330
rect 66 328 70 332
rect 112 328 116 332
rect 122 328 126 332
rect 142 328 146 332
rect 152 328 156 332
rect 172 328 176 332
rect 182 328 186 332
rect 202 328 206 332
rect 212 328 216 332
rect 232 328 236 332
rect 365 329 369 333
rect 375 329 379 333
rect 395 329 399 333
rect 405 329 409 333
rect 425 329 429 333
rect 435 329 439 333
rect 455 329 459 333
rect 465 329 469 333
rect 485 329 489 333
rect 530 328 534 332
rect 582 326 586 330
rect 592 326 596 330
rect 298 322 302 326
rect 6 316 10 320
rect 36 318 40 322
rect 46 318 50 322
rect 66 318 70 322
rect 112 316 116 320
rect 122 316 126 320
rect 142 316 146 320
rect 152 316 156 320
rect 172 316 176 320
rect 182 316 186 320
rect 202 316 206 320
rect 212 316 216 320
rect 232 316 236 320
rect 365 317 369 321
rect 375 317 379 321
rect 395 317 399 321
rect 405 317 409 321
rect 425 317 429 321
rect 435 317 439 321
rect 455 317 459 321
rect 465 317 469 321
rect 485 317 489 321
rect 530 318 534 322
rect 298 312 302 316
rect 544 315 548 319
rect 554 315 558 319
rect 582 316 586 320
rect 592 316 596 320
rect 6 306 10 310
rect 36 308 40 312
rect 46 308 50 312
rect 66 308 70 312
rect 530 308 534 312
rect 544 305 548 309
rect 554 305 558 309
rect 582 306 586 310
rect 592 306 596 310
rect 6 296 10 300
rect 36 298 40 302
rect 46 298 50 302
rect 66 298 70 302
rect 530 298 534 302
rect 544 295 548 299
rect 554 295 558 299
rect 582 296 586 300
rect 592 296 596 300
rect 6 286 10 290
rect 66 288 70 292
rect 530 288 534 292
rect 582 286 586 290
rect 592 286 596 290
rect 298 282 302 286
rect 6 276 10 280
rect 36 278 40 282
rect 46 278 50 282
rect 66 278 70 282
rect 530 278 534 282
rect 544 275 548 279
rect 554 275 558 279
rect 582 276 586 280
rect 592 276 596 280
rect 6 266 10 270
rect 36 268 40 272
rect 46 268 50 272
rect 66 268 70 272
rect 530 268 534 272
rect 114 262 118 266
rect 124 262 128 266
rect 134 262 138 266
rect 144 262 148 266
rect 154 262 158 266
rect 164 262 168 266
rect 174 262 178 266
rect 184 262 188 266
rect 194 262 198 266
rect 204 262 208 266
rect 214 262 218 266
rect 224 262 228 266
rect 234 262 238 266
rect 298 262 302 266
rect 362 262 366 266
rect 372 262 376 266
rect 382 262 386 266
rect 392 262 396 266
rect 402 262 406 266
rect 412 262 416 266
rect 422 262 426 266
rect 432 262 436 266
rect 442 262 446 266
rect 452 262 456 266
rect 462 262 466 266
rect 472 262 476 266
rect 482 262 486 266
rect 544 265 548 269
rect 554 265 558 269
rect 582 266 586 270
rect 592 266 596 270
rect 6 256 10 260
rect 36 258 40 262
rect 46 258 50 262
rect 66 258 70 262
rect 530 258 534 262
rect 114 252 118 256
rect 124 252 128 256
rect 134 252 138 256
rect 144 252 148 256
rect 154 252 158 256
rect 164 252 168 256
rect 174 252 178 256
rect 184 252 188 256
rect 194 252 198 256
rect 204 252 208 256
rect 214 252 218 256
rect 224 252 228 256
rect 234 252 238 256
rect 298 252 302 256
rect 362 252 366 256
rect 372 252 376 256
rect 382 252 386 256
rect 392 252 396 256
rect 402 252 406 256
rect 412 252 416 256
rect 422 252 426 256
rect 432 252 436 256
rect 442 252 446 256
rect 452 252 456 256
rect 462 252 466 256
rect 472 252 476 256
rect 482 252 486 256
rect 544 255 548 259
rect 554 255 558 259
rect 582 256 586 260
rect 592 256 596 260
rect 6 246 10 250
rect 66 248 70 252
rect 530 248 534 252
rect 582 246 586 250
rect 592 246 596 250
rect 6 236 10 240
rect 36 238 40 242
rect 46 238 50 242
rect 66 238 70 242
rect 530 238 534 242
rect 298 232 302 236
rect 544 235 548 239
rect 554 235 558 239
rect 582 236 586 240
rect 592 236 596 240
rect 6 226 10 230
rect 36 228 40 232
rect 46 228 50 232
rect 66 228 70 232
rect 530 228 534 232
rect 298 222 302 226
rect 544 225 548 229
rect 554 225 558 229
rect 582 226 586 230
rect 592 226 596 230
rect 6 216 10 220
rect 36 218 40 222
rect 46 218 50 222
rect 66 218 70 222
rect 530 218 534 222
rect 544 215 548 219
rect 554 215 558 219
rect 582 216 586 220
rect 592 216 596 220
rect 6 206 10 210
rect 66 208 70 212
rect 530 208 534 212
rect 582 206 586 210
rect 592 206 596 210
rect 298 202 302 206
rect 6 196 10 200
rect 36 198 40 202
rect 46 198 50 202
rect 66 198 70 202
rect 111 198 115 202
rect 121 198 125 202
rect 141 198 145 202
rect 151 198 155 202
rect 171 198 175 202
rect 181 198 185 202
rect 201 198 205 202
rect 211 198 215 202
rect 231 198 235 202
rect 366 198 370 202
rect 376 198 380 202
rect 396 198 400 202
rect 406 198 410 202
rect 426 198 430 202
rect 436 198 440 202
rect 456 198 460 202
rect 466 198 470 202
rect 486 198 490 202
rect 530 198 534 202
rect 298 192 302 196
rect 544 195 548 199
rect 554 195 558 199
rect 582 196 586 200
rect 592 196 596 200
rect 6 186 10 190
rect 36 188 40 192
rect 46 188 50 192
rect 66 188 70 192
rect 111 186 115 190
rect 121 186 125 190
rect 141 186 145 190
rect 151 186 155 190
rect 171 186 175 190
rect 181 186 185 190
rect 201 186 205 190
rect 211 186 215 190
rect 231 186 235 190
rect 366 186 370 190
rect 376 186 380 190
rect 396 186 400 190
rect 406 186 410 190
rect 426 186 430 190
rect 436 186 440 190
rect 456 186 460 190
rect 466 186 470 190
rect 486 186 490 190
rect 530 188 534 192
rect 544 185 548 189
rect 554 185 558 189
rect 582 186 586 190
rect 592 186 596 190
rect 6 176 10 180
rect 36 178 40 182
rect 46 178 50 182
rect 66 178 70 182
rect 530 178 534 182
rect 298 172 302 176
rect 544 175 548 179
rect 554 175 558 179
rect 582 176 586 180
rect 592 176 596 180
rect 6 166 10 170
rect 66 168 70 172
rect 530 168 534 172
rect 582 166 586 170
rect 592 166 596 170
rect 6 156 10 160
rect 36 158 40 162
rect 46 158 50 162
rect 66 158 70 162
rect 530 158 534 162
rect 544 155 548 159
rect 554 155 558 159
rect 582 156 586 160
rect 592 156 596 160
rect 6 146 10 150
rect 36 148 40 152
rect 46 148 50 152
rect 66 148 70 152
rect 530 148 534 152
rect 298 142 302 146
rect 544 145 548 149
rect 554 145 558 149
rect 582 146 586 150
rect 592 146 596 150
rect 6 136 10 140
rect 36 138 40 142
rect 46 138 50 142
rect 66 138 70 142
rect 530 138 534 142
rect 114 132 118 136
rect 124 132 128 136
rect 134 132 138 136
rect 144 132 148 136
rect 154 132 158 136
rect 164 132 168 136
rect 174 132 178 136
rect 184 132 188 136
rect 194 132 198 136
rect 204 132 208 136
rect 214 132 218 136
rect 224 132 228 136
rect 234 132 238 136
rect 298 132 302 136
rect 362 132 366 136
rect 372 132 376 136
rect 382 132 386 136
rect 392 132 396 136
rect 402 132 406 136
rect 412 132 416 136
rect 422 132 426 136
rect 432 132 436 136
rect 442 132 446 136
rect 452 132 456 136
rect 462 132 466 136
rect 472 132 476 136
rect 482 132 486 136
rect 544 135 548 139
rect 554 135 558 139
rect 582 136 586 140
rect 592 136 596 140
rect 6 126 10 130
rect 66 128 70 132
rect 530 128 534 132
rect 582 126 586 130
rect 592 126 596 130
rect 114 122 118 126
rect 124 122 128 126
rect 134 122 138 126
rect 144 122 148 126
rect 154 122 158 126
rect 164 122 168 126
rect 174 122 178 126
rect 184 122 188 126
rect 194 122 198 126
rect 204 122 208 126
rect 214 122 218 126
rect 224 122 228 126
rect 234 122 238 126
rect 362 122 366 126
rect 372 122 376 126
rect 382 122 386 126
rect 392 122 396 126
rect 402 122 406 126
rect 412 122 416 126
rect 422 122 426 126
rect 432 122 436 126
rect 442 122 446 126
rect 452 122 456 126
rect 462 122 466 126
rect 472 122 476 126
rect 482 122 486 126
rect 6 116 10 120
rect 36 118 40 122
rect 46 118 50 122
rect 66 118 70 122
rect 530 118 534 122
rect 298 112 302 116
rect 544 115 548 119
rect 554 115 558 119
rect 582 116 586 120
rect 592 116 596 120
rect 6 106 10 110
rect 36 108 40 112
rect 46 108 50 112
rect 66 108 70 112
rect 530 108 534 112
rect 544 105 548 109
rect 554 105 558 109
rect 582 106 586 110
rect 592 106 596 110
rect 6 96 10 100
rect 36 98 40 102
rect 46 98 50 102
rect 66 98 70 102
rect 530 98 534 102
rect 544 95 548 99
rect 554 95 558 99
rect 582 96 586 100
rect 592 96 596 100
rect 6 86 10 90
rect 66 88 70 92
rect 530 88 534 92
rect 582 86 586 90
rect 592 86 596 90
rect 6 76 10 80
rect 36 78 40 82
rect 46 78 50 82
rect 544 75 548 79
rect 554 75 558 79
rect 582 76 586 80
rect 592 76 596 80
rect 6 66 10 70
rect 36 68 40 72
rect 46 68 50 72
rect 80 69 84 73
rect 109 68 113 72
rect 120 68 124 72
rect 130 68 134 72
rect 140 68 144 72
rect 150 68 154 72
rect 160 68 164 72
rect 170 68 174 72
rect 180 68 184 72
rect 190 68 194 72
rect 200 68 204 72
rect 210 68 214 72
rect 220 68 224 72
rect 230 68 234 72
rect 366 68 370 72
rect 376 68 380 72
rect 386 68 390 72
rect 396 68 400 72
rect 406 68 410 72
rect 416 68 420 72
rect 426 68 430 72
rect 436 68 440 72
rect 446 68 450 72
rect 456 68 460 72
rect 466 68 470 72
rect 476 68 480 72
rect 486 68 490 72
rect 544 65 548 69
rect 554 65 558 69
rect 582 66 586 70
rect 592 66 596 70
rect 6 56 10 60
rect 80 58 84 62
rect 109 58 113 62
rect 130 56 134 60
rect 150 56 154 60
rect 170 56 174 60
rect 190 56 194 60
rect 210 56 214 60
rect 230 56 234 60
rect 366 56 370 60
rect 386 56 390 60
rect 406 56 410 60
rect 426 56 430 60
rect 446 56 450 60
rect 466 56 470 60
rect 486 58 490 62
rect 582 56 586 60
rect 592 56 596 60
rect 36 52 40 56
rect 50 52 54 56
rect 60 52 64 56
rect 70 52 74 56
rect 528 52 532 56
rect 538 52 542 56
rect 554 52 558 56
rect 6 46 10 50
rect 109 48 113 52
rect 130 46 134 50
rect 150 46 154 50
rect 170 46 174 50
rect 190 46 194 50
rect 210 46 214 50
rect 230 46 234 50
rect 366 46 370 50
rect 386 46 390 50
rect 406 46 410 50
rect 426 46 430 50
rect 446 46 450 50
rect 466 46 470 50
rect 486 48 490 52
rect 582 46 586 50
rect 592 46 596 50
rect 6 36 10 40
rect 80 38 84 42
rect 109 38 113 42
rect 130 36 134 40
rect 150 36 154 40
rect 170 36 174 40
rect 190 36 194 40
rect 210 36 214 40
rect 230 36 234 40
rect 366 36 370 40
rect 386 36 390 40
rect 406 36 410 40
rect 426 36 430 40
rect 446 36 450 40
rect 466 36 470 40
rect 486 38 490 42
rect 50 32 54 36
rect 60 32 64 36
rect 70 32 74 36
rect 528 34 532 38
rect 582 36 586 40
rect 592 36 596 40
rect 554 32 558 36
rect 6 26 10 30
rect 582 26 586 30
rect 592 26 596 30
rect 6 16 10 20
rect 582 16 586 20
rect 592 16 596 20
rect 6 6 10 10
rect 16 4 20 8
rect 26 4 30 8
rect 36 4 40 8
rect 48 4 52 8
rect 58 6 62 10
rect 68 6 72 10
rect 78 4 82 8
rect 88 4 92 8
rect 98 4 102 8
rect 108 4 112 8
rect 118 6 122 10
rect 128 6 132 10
rect 138 6 142 10
rect 148 6 152 10
rect 158 6 162 10
rect 168 6 172 10
rect 178 6 182 10
rect 188 6 192 10
rect 198 6 202 10
rect 208 6 212 10
rect 218 6 222 10
rect 228 6 232 10
rect 238 6 242 10
rect 248 6 252 10
rect 258 6 262 10
rect 268 6 272 10
rect 278 6 282 10
rect 288 6 292 10
rect 298 6 302 10
rect 308 6 312 10
rect 318 6 322 10
rect 328 6 332 10
rect 340 6 344 10
rect 350 6 354 10
rect 360 6 364 10
rect 370 6 374 10
rect 380 6 384 10
rect 390 6 394 10
rect 400 6 404 10
rect 410 6 414 10
rect 420 6 424 10
rect 430 6 434 10
rect 440 6 444 10
rect 450 6 454 10
rect 460 6 464 10
rect 470 6 474 10
rect 480 4 484 8
rect 490 4 494 8
rect 500 4 504 8
rect 510 4 514 8
rect 520 4 524 8
rect 530 4 534 8
rect 540 6 544 10
rect 550 6 554 10
rect 560 6 564 10
rect 570 6 574 10
rect 580 6 584 10
rect 592 6 596 10
<< gv1 >>
rect 30 1302 34 1306
rect 40 1302 44 1306
rect 50 1302 54 1306
rect 60 1302 64 1306
rect 70 1302 74 1306
rect 80 1302 84 1306
rect 90 1302 94 1306
rect 100 1302 104 1306
rect 110 1302 114 1306
rect 120 1302 124 1306
rect 130 1302 134 1306
rect 140 1302 144 1306
rect 150 1302 154 1306
rect 160 1302 164 1306
rect 170 1302 174 1306
rect 180 1302 184 1306
rect 190 1302 194 1306
rect 200 1302 204 1306
rect 210 1302 214 1306
rect 220 1302 224 1306
rect 376 1304 380 1308
rect 386 1304 390 1308
rect 396 1304 400 1308
rect 406 1304 410 1308
rect 416 1304 420 1308
rect 426 1304 430 1308
rect 436 1304 440 1308
rect 446 1304 450 1308
rect 456 1304 460 1308
rect 466 1304 470 1308
rect 476 1304 480 1308
rect 486 1304 490 1308
rect 496 1304 500 1308
rect 506 1304 510 1308
rect 516 1304 520 1308
rect 526 1304 530 1308
rect 536 1304 540 1308
rect 546 1304 550 1308
rect 556 1304 560 1308
rect 566 1304 570 1308
rect 30 1292 34 1296
rect 566 1294 570 1298
rect 30 1282 34 1286
rect 42 1284 46 1288
rect 52 1284 56 1288
rect 62 1284 66 1288
rect 72 1284 76 1288
rect 82 1284 86 1288
rect 124 1284 128 1288
rect 154 1284 158 1288
rect 184 1284 188 1288
rect 214 1284 218 1288
rect 378 1284 382 1288
rect 408 1284 412 1288
rect 438 1284 442 1288
rect 468 1284 472 1288
rect 510 1284 514 1288
rect 520 1284 524 1288
rect 530 1284 534 1288
rect 544 1284 548 1288
rect 554 1284 558 1288
rect 566 1284 570 1288
rect 298 1278 302 1282
rect 30 1272 34 1276
rect 62 1274 66 1278
rect 72 1274 76 1278
rect 82 1274 86 1278
rect 124 1274 128 1278
rect 154 1274 158 1278
rect 184 1274 188 1278
rect 214 1274 218 1278
rect 378 1274 382 1278
rect 408 1274 412 1278
rect 438 1274 442 1278
rect 468 1274 472 1278
rect 510 1274 514 1278
rect 520 1274 524 1278
rect 530 1274 534 1278
rect 566 1274 570 1278
rect 30 1262 34 1266
rect 62 1264 66 1268
rect 72 1264 76 1268
rect 82 1264 86 1268
rect 124 1264 128 1268
rect 154 1264 158 1268
rect 184 1264 188 1268
rect 214 1264 218 1268
rect 378 1264 382 1268
rect 408 1264 412 1268
rect 438 1264 442 1268
rect 468 1264 472 1268
rect 510 1264 514 1268
rect 520 1264 524 1268
rect 530 1264 534 1268
rect 566 1264 570 1268
rect 30 1252 34 1256
rect 566 1254 570 1258
rect 30 1242 34 1246
rect 42 1244 46 1248
rect 52 1244 56 1248
rect 66 1245 70 1249
rect 530 1244 534 1248
rect 544 1244 548 1248
rect 554 1244 558 1248
rect 566 1244 570 1248
rect 86 1238 90 1242
rect 96 1238 100 1242
rect 106 1238 110 1242
rect 116 1238 120 1242
rect 126 1238 130 1242
rect 136 1238 140 1242
rect 146 1238 150 1242
rect 156 1238 160 1242
rect 166 1238 170 1242
rect 176 1238 180 1242
rect 186 1238 190 1242
rect 196 1238 200 1242
rect 206 1238 210 1242
rect 216 1238 220 1242
rect 226 1238 230 1242
rect 298 1238 302 1242
rect 370 1238 374 1242
rect 380 1238 384 1242
rect 390 1238 394 1242
rect 400 1238 404 1242
rect 410 1238 414 1242
rect 420 1238 424 1242
rect 430 1238 434 1242
rect 440 1238 444 1242
rect 450 1238 454 1242
rect 460 1238 464 1242
rect 470 1238 474 1242
rect 480 1238 484 1242
rect 490 1238 494 1242
rect 500 1238 504 1242
rect 510 1238 514 1242
rect 30 1232 34 1236
rect 566 1234 570 1238
rect 84 1227 88 1231
rect 94 1227 98 1231
rect 30 1222 34 1226
rect 500 1223 504 1227
rect 510 1223 514 1227
rect 566 1224 570 1228
rect 84 1217 88 1221
rect 94 1217 98 1221
rect 30 1212 34 1216
rect 500 1213 504 1217
rect 510 1213 514 1217
rect 566 1214 570 1218
rect 30 1202 34 1206
rect 42 1204 46 1208
rect 52 1204 56 1208
rect 84 1207 88 1211
rect 94 1207 98 1211
rect 500 1203 504 1207
rect 510 1203 514 1207
rect 544 1204 548 1208
rect 554 1204 558 1208
rect 566 1204 570 1208
rect 84 1197 88 1201
rect 94 1197 98 1201
rect 298 1198 302 1202
rect 30 1192 34 1196
rect 500 1193 504 1197
rect 510 1193 514 1197
rect 566 1194 570 1198
rect 84 1187 88 1191
rect 94 1187 98 1191
rect 30 1182 34 1186
rect 500 1183 504 1187
rect 510 1183 514 1187
rect 566 1184 570 1188
rect 30 1172 34 1176
rect 66 1173 70 1177
rect 86 1174 90 1178
rect 96 1174 100 1178
rect 106 1174 110 1178
rect 116 1174 120 1178
rect 126 1174 130 1178
rect 136 1174 140 1178
rect 146 1174 150 1178
rect 156 1174 160 1178
rect 166 1174 170 1178
rect 176 1174 180 1178
rect 186 1174 190 1178
rect 196 1174 200 1178
rect 206 1174 210 1178
rect 216 1174 220 1178
rect 226 1174 230 1178
rect 370 1172 374 1176
rect 380 1172 384 1176
rect 390 1172 394 1176
rect 400 1172 404 1176
rect 410 1172 414 1176
rect 420 1172 424 1176
rect 430 1172 434 1176
rect 440 1172 444 1176
rect 450 1172 454 1176
rect 460 1172 464 1176
rect 470 1172 474 1176
rect 480 1172 484 1176
rect 490 1172 494 1176
rect 500 1172 504 1176
rect 510 1172 514 1176
rect 566 1174 570 1178
rect 530 1170 534 1174
rect 30 1162 34 1166
rect 42 1164 46 1168
rect 52 1164 56 1168
rect 66 1163 70 1167
rect 544 1164 548 1168
rect 554 1164 558 1168
rect 566 1164 570 1168
rect 298 1158 302 1162
rect 530 1160 534 1164
rect 30 1152 34 1156
rect 66 1153 70 1157
rect 566 1154 570 1158
rect 530 1150 534 1154
rect 30 1142 34 1146
rect 66 1143 70 1147
rect 85 1146 89 1150
rect 95 1146 99 1150
rect 105 1146 109 1150
rect 115 1146 119 1150
rect 145 1146 149 1150
rect 175 1146 179 1150
rect 205 1146 209 1150
rect 390 1146 394 1150
rect 420 1146 424 1150
rect 450 1146 454 1150
rect 480 1146 484 1150
rect 490 1146 494 1150
rect 500 1146 504 1150
rect 510 1146 514 1150
rect 566 1144 570 1148
rect 530 1140 534 1144
rect 30 1132 34 1136
rect 66 1133 70 1137
rect 85 1134 89 1138
rect 95 1134 99 1138
rect 105 1134 109 1138
rect 115 1134 119 1138
rect 145 1134 149 1138
rect 175 1134 179 1138
rect 205 1134 209 1138
rect 390 1134 394 1138
rect 420 1134 424 1138
rect 450 1134 454 1138
rect 480 1134 484 1138
rect 490 1134 494 1138
rect 500 1134 504 1138
rect 510 1134 514 1138
rect 566 1134 570 1138
rect 530 1130 534 1134
rect 30 1122 34 1126
rect 42 1124 46 1128
rect 52 1124 56 1128
rect 66 1123 70 1127
rect 544 1124 548 1128
rect 554 1124 558 1128
rect 566 1124 570 1128
rect 298 1118 302 1122
rect 530 1120 534 1124
rect 30 1112 34 1116
rect 66 1113 70 1117
rect 566 1114 570 1118
rect 86 1107 90 1111
rect 96 1107 100 1111
rect 106 1107 110 1111
rect 116 1107 120 1111
rect 126 1107 130 1111
rect 136 1107 140 1111
rect 146 1107 150 1111
rect 156 1107 160 1111
rect 166 1107 170 1111
rect 176 1107 180 1111
rect 186 1107 190 1111
rect 196 1107 200 1111
rect 206 1107 210 1111
rect 216 1107 220 1111
rect 226 1107 230 1111
rect 370 1108 374 1112
rect 380 1108 384 1112
rect 390 1108 394 1112
rect 400 1108 404 1112
rect 410 1108 414 1112
rect 420 1108 424 1112
rect 430 1108 434 1112
rect 440 1108 444 1112
rect 450 1108 454 1112
rect 460 1108 464 1112
rect 470 1108 474 1112
rect 480 1108 484 1112
rect 490 1108 494 1112
rect 500 1108 504 1112
rect 510 1108 514 1112
rect 530 1110 534 1114
rect 30 1102 34 1106
rect 566 1104 570 1108
rect 86 1097 90 1101
rect 96 1097 100 1101
rect 500 1097 504 1101
rect 510 1097 514 1101
rect 30 1092 34 1096
rect 566 1094 570 1098
rect 30 1082 34 1086
rect 42 1084 46 1088
rect 52 1084 56 1088
rect 86 1087 90 1091
rect 96 1087 100 1091
rect 500 1087 504 1091
rect 510 1087 514 1091
rect 544 1084 548 1088
rect 554 1084 558 1088
rect 566 1084 570 1088
rect 86 1077 90 1081
rect 96 1077 100 1081
rect 298 1078 302 1082
rect 500 1077 504 1081
rect 510 1077 514 1081
rect 30 1072 34 1076
rect 566 1074 570 1078
rect 86 1067 90 1071
rect 96 1067 100 1071
rect 500 1067 504 1071
rect 510 1067 514 1071
rect 30 1062 34 1066
rect 566 1064 570 1068
rect 86 1057 90 1061
rect 96 1057 100 1061
rect 500 1057 504 1061
rect 510 1057 514 1061
rect 30 1052 34 1056
rect 566 1054 570 1058
rect 30 1042 34 1046
rect 42 1044 46 1048
rect 52 1044 56 1048
rect 66 1043 70 1047
rect 86 1046 90 1050
rect 96 1046 100 1050
rect 106 1046 110 1050
rect 116 1046 120 1050
rect 126 1046 130 1050
rect 136 1046 140 1050
rect 146 1046 150 1050
rect 156 1046 160 1050
rect 166 1046 170 1050
rect 176 1046 180 1050
rect 186 1046 190 1050
rect 196 1046 200 1050
rect 206 1046 210 1050
rect 216 1046 220 1050
rect 226 1046 230 1050
rect 370 1046 374 1050
rect 380 1046 384 1050
rect 390 1046 394 1050
rect 400 1046 404 1050
rect 410 1046 414 1050
rect 420 1046 424 1050
rect 430 1046 434 1050
rect 440 1046 444 1050
rect 450 1046 454 1050
rect 460 1046 464 1050
rect 470 1046 474 1050
rect 480 1046 484 1050
rect 490 1046 494 1050
rect 500 1046 504 1050
rect 510 1046 514 1050
rect 530 1043 534 1047
rect 544 1044 548 1048
rect 554 1044 558 1048
rect 566 1044 570 1048
rect 298 1038 302 1042
rect 30 1032 34 1036
rect 66 1033 70 1037
rect 530 1033 534 1037
rect 566 1034 570 1038
rect 30 1022 34 1026
rect 66 1023 70 1027
rect 530 1023 534 1027
rect 566 1024 570 1028
rect 84 1018 88 1022
rect 94 1018 98 1022
rect 104 1018 108 1022
rect 114 1018 118 1022
rect 144 1018 148 1022
rect 174 1018 178 1022
rect 204 1018 208 1022
rect 389 1018 393 1022
rect 419 1018 423 1022
rect 449 1018 453 1022
rect 479 1018 483 1022
rect 489 1018 493 1022
rect 499 1018 503 1022
rect 509 1018 513 1022
rect 30 1012 34 1016
rect 66 1013 70 1017
rect 530 1013 534 1017
rect 566 1014 570 1018
rect 30 1002 34 1006
rect 42 1004 46 1008
rect 52 1004 56 1008
rect 66 1003 70 1007
rect 84 1006 88 1010
rect 94 1006 98 1010
rect 104 1006 108 1010
rect 114 1006 118 1010
rect 144 1006 148 1010
rect 174 1006 178 1010
rect 204 1006 208 1010
rect 389 1006 393 1010
rect 419 1006 423 1010
rect 449 1006 453 1010
rect 479 1006 483 1010
rect 489 1006 493 1010
rect 499 1006 503 1010
rect 509 1006 513 1010
rect 530 1003 534 1007
rect 544 1004 548 1008
rect 554 1004 558 1008
rect 566 1004 570 1008
rect 298 998 302 1002
rect 30 992 34 996
rect 66 993 70 997
rect 530 993 534 997
rect 566 994 570 998
rect 30 982 34 986
rect 66 983 70 987
rect 86 980 90 984
rect 96 980 100 984
rect 106 980 110 984
rect 116 980 120 984
rect 126 980 130 984
rect 136 980 140 984
rect 146 980 150 984
rect 156 980 160 984
rect 166 980 170 984
rect 176 980 180 984
rect 186 980 190 984
rect 196 980 200 984
rect 206 980 210 984
rect 216 980 220 984
rect 226 980 230 984
rect 370 980 374 984
rect 380 980 384 984
rect 390 980 394 984
rect 400 980 404 984
rect 410 980 414 984
rect 420 980 424 984
rect 430 980 434 984
rect 440 980 444 984
rect 450 980 454 984
rect 460 980 464 984
rect 470 980 474 984
rect 480 980 484 984
rect 490 980 494 984
rect 500 980 504 984
rect 510 980 514 984
rect 530 983 534 987
rect 566 984 570 988
rect 30 972 34 976
rect 566 974 570 978
rect 86 969 90 973
rect 96 969 100 973
rect 502 968 506 972
rect 512 968 516 972
rect 30 962 34 966
rect 42 964 46 968
rect 52 964 56 968
rect 544 964 548 968
rect 554 964 558 968
rect 566 964 570 968
rect 86 959 90 963
rect 96 959 100 963
rect 298 958 302 962
rect 502 958 506 962
rect 512 958 516 962
rect 30 952 34 956
rect 566 954 570 958
rect 86 949 90 953
rect 96 949 100 953
rect 502 948 506 952
rect 512 948 516 952
rect 30 942 34 946
rect 566 944 570 948
rect 86 939 90 943
rect 96 939 100 943
rect 502 938 506 942
rect 512 938 516 942
rect 30 932 34 936
rect 566 934 570 938
rect 86 929 90 933
rect 96 929 100 933
rect 502 928 506 932
rect 512 928 516 932
rect 30 922 34 926
rect 42 924 46 928
rect 52 924 56 928
rect 544 924 548 928
rect 554 924 558 928
rect 566 924 570 928
rect 84 916 88 920
rect 94 916 98 920
rect 104 916 108 920
rect 114 916 118 920
rect 124 916 128 920
rect 134 916 138 920
rect 144 916 148 920
rect 154 916 158 920
rect 164 916 168 920
rect 174 916 178 920
rect 184 916 188 920
rect 194 916 198 920
rect 204 916 208 920
rect 214 916 218 920
rect 224 916 228 920
rect 298 918 302 922
rect 372 916 376 920
rect 382 916 386 920
rect 392 916 396 920
rect 402 916 406 920
rect 412 916 416 920
rect 422 916 426 920
rect 432 916 436 920
rect 442 916 446 920
rect 452 916 456 920
rect 462 916 466 920
rect 472 916 476 920
rect 482 916 486 920
rect 492 916 496 920
rect 502 916 506 920
rect 512 916 516 920
rect 30 912 34 916
rect 566 914 570 918
rect 30 902 34 906
rect 566 904 570 908
rect 30 892 34 896
rect 566 894 570 898
rect 82 888 86 892
rect 93 888 97 892
rect 104 888 108 892
rect 115 888 119 892
rect 145 888 149 892
rect 175 888 179 892
rect 205 888 209 892
rect 391 888 395 892
rect 421 888 425 892
rect 451 888 455 892
rect 481 888 485 892
rect 492 888 496 892
rect 503 888 507 892
rect 514 888 518 892
rect 30 882 34 886
rect 42 884 46 888
rect 52 884 56 888
rect 544 884 548 888
rect 554 884 558 888
rect 566 884 570 888
rect 95 876 99 880
rect 115 876 119 880
rect 145 876 149 880
rect 175 876 179 880
rect 205 876 209 880
rect 298 878 302 882
rect 391 876 395 880
rect 421 876 425 880
rect 451 876 455 880
rect 481 876 485 880
rect 501 876 505 880
rect 66 864 70 868
rect 76 864 80 868
rect 520 864 524 868
rect 530 864 534 868
rect 32 844 36 848
rect 42 844 46 848
rect 52 844 56 848
rect 80 844 84 848
rect 90 844 94 848
rect 100 844 104 848
rect 110 844 114 848
rect 120 844 124 848
rect 130 844 134 848
rect 140 844 144 848
rect 150 844 154 848
rect 160 844 164 848
rect 170 844 174 848
rect 180 844 184 848
rect 190 844 194 848
rect 200 844 204 848
rect 210 844 214 848
rect 220 844 224 848
rect 298 844 302 848
rect 370 844 374 848
rect 380 844 384 848
rect 390 844 394 848
rect 400 844 404 848
rect 410 844 414 848
rect 420 844 424 848
rect 430 844 434 848
rect 440 844 444 848
rect 450 844 454 848
rect 460 844 464 848
rect 470 844 474 848
rect 480 844 484 848
rect 490 844 494 848
rect 500 844 504 848
rect 510 844 514 848
rect 520 844 524 848
rect 530 844 534 848
rect 540 844 544 848
rect 550 844 554 848
rect 560 844 564 848
rect 570 844 574 848
rect 592 817 596 821
rect 16 812 20 816
rect 28 812 32 816
rect 38 812 42 816
rect 48 812 52 816
rect 80 812 84 816
rect 90 812 94 816
rect 100 812 104 816
rect 110 812 114 816
rect 120 812 124 816
rect 130 812 134 816
rect 140 812 144 816
rect 150 812 154 816
rect 160 812 164 816
rect 170 812 174 816
rect 180 812 184 816
rect 190 812 194 816
rect 200 812 204 816
rect 210 812 214 816
rect 16 802 20 806
rect 592 797 596 801
rect 16 792 20 796
rect 16 780 20 784
rect 578 778 582 782
rect 592 777 596 781
rect 16 770 20 774
rect 16 760 20 764
rect 592 757 596 761
rect 16 750 20 754
rect 46 744 50 748
rect 388 744 392 748
rect 452 745 456 749
rect 484 745 488 749
rect 516 745 520 749
rect 548 745 552 749
rect 580 745 584 749
rect 16 740 20 744
rect 96 740 100 744
rect 128 740 132 744
rect 160 740 164 744
rect 192 740 196 744
rect 224 740 228 744
rect 592 737 596 741
rect 16 730 20 734
rect 46 724 50 728
rect 16 720 20 724
rect 96 720 100 724
rect 128 720 132 724
rect 160 720 164 724
rect 192 720 196 724
rect 224 720 228 724
rect 240 722 244 726
rect 272 722 276 726
rect 388 724 392 728
rect 420 722 424 726
rect 452 725 456 729
rect 484 725 488 729
rect 516 725 520 729
rect 548 725 552 729
rect 580 725 584 729
rect 592 717 596 721
rect 16 710 20 714
rect 582 699 586 703
rect 592 697 596 701
rect 208 689 212 693
rect 262 689 266 693
rect 506 687 510 691
rect 42 672 46 676
rect 52 672 56 676
rect 186 672 190 676
rect 196 672 200 676
rect 250 672 254 676
rect 260 672 264 676
rect 390 675 394 679
rect 400 675 404 679
rect 410 675 414 679
rect 420 675 424 679
rect 436 672 440 676
rect 446 672 450 676
rect 557 672 561 676
rect 567 672 571 676
rect 140 657 144 661
rect 210 657 214 661
rect 286 657 290 661
rect 410 657 414 661
rect 506 657 510 661
rect 4 636 8 640
rect 592 638 596 642
rect 16 630 20 634
rect 46 625 50 629
rect 96 625 100 629
rect 224 625 228 629
rect 16 620 20 624
rect 272 623 276 627
rect 304 623 308 627
rect 4 616 8 620
rect 128 617 132 621
rect 160 617 164 621
rect 192 617 196 621
rect 388 617 392 621
rect 420 617 424 621
rect 452 617 456 621
rect 484 617 488 621
rect 516 617 520 621
rect 548 617 552 621
rect 580 617 584 621
rect 592 618 596 622
rect 16 610 20 614
rect 46 605 50 609
rect 96 605 100 609
rect 224 605 228 609
rect 16 600 20 604
rect 4 596 8 600
rect 128 597 132 601
rect 160 597 164 601
rect 192 597 196 601
rect 388 597 392 601
rect 420 597 424 601
rect 452 597 456 601
rect 484 597 488 601
rect 516 597 520 601
rect 548 597 552 601
rect 580 597 584 601
rect 592 598 596 602
rect 16 590 20 594
rect 46 585 50 589
rect 96 585 100 589
rect 160 587 164 591
rect 224 585 228 589
rect 388 587 392 591
rect 420 587 424 591
rect 452 587 456 591
rect 484 587 488 591
rect 516 587 520 591
rect 548 587 552 591
rect 16 580 20 584
rect 4 576 8 580
rect 128 577 132 581
rect 192 577 196 581
rect 580 577 584 581
rect 592 578 596 582
rect 16 570 20 574
rect 46 565 50 569
rect 96 565 100 569
rect 224 565 228 569
rect 16 560 20 564
rect 4 556 8 560
rect 128 557 132 561
rect 160 557 164 561
rect 192 557 196 561
rect 388 557 392 561
rect 420 557 424 561
rect 452 557 456 561
rect 484 557 488 561
rect 516 557 520 561
rect 548 557 552 561
rect 580 557 584 561
rect 592 558 596 562
rect 16 550 20 554
rect 4 536 8 540
rect 582 535 586 539
rect 592 538 596 542
rect 4 516 8 520
rect 592 518 596 522
rect 36 496 40 500
rect 46 496 50 500
rect 56 496 60 500
rect 66 496 70 500
rect 108 496 112 500
rect 118 496 122 500
rect 128 496 132 500
rect 138 496 142 500
rect 148 496 152 500
rect 158 496 162 500
rect 168 496 172 500
rect 178 496 182 500
rect 188 496 192 500
rect 198 496 202 500
rect 208 496 212 500
rect 224 496 228 500
rect 234 496 238 500
rect 391 496 395 500
rect 401 496 405 500
rect 411 496 415 500
rect 421 496 425 500
rect 431 496 435 500
rect 441 496 445 500
rect 451 496 455 500
rect 529 496 533 500
rect 539 496 543 500
rect 549 496 553 500
rect 559 496 563 500
rect 569 496 573 500
rect 80 478 84 482
rect 529 478 533 482
rect 80 466 84 470
rect 529 466 533 470
rect 130 460 134 464
rect 160 460 164 464
rect 190 460 194 464
rect 220 460 224 464
rect 386 460 390 464
rect 416 460 420 464
rect 446 460 450 464
rect 476 460 480 464
rect 298 452 302 456
rect 566 453 570 457
rect 36 448 40 452
rect 46 448 50 452
rect 66 446 70 450
rect 130 448 134 452
rect 160 448 164 452
rect 190 448 194 452
rect 220 448 224 452
rect 386 448 390 452
rect 416 448 420 452
rect 446 448 450 452
rect 476 448 480 452
rect 544 445 548 449
rect 554 445 558 449
rect 566 443 570 447
rect 566 433 570 437
rect 110 423 114 427
rect 120 423 124 427
rect 130 423 134 427
rect 140 423 144 427
rect 150 423 154 427
rect 160 423 164 427
rect 170 423 174 427
rect 180 423 184 427
rect 190 423 194 427
rect 200 423 204 427
rect 210 423 214 427
rect 220 423 224 427
rect 230 423 234 427
rect 298 422 302 426
rect 366 423 370 427
rect 376 423 380 427
rect 386 423 390 427
rect 396 423 400 427
rect 406 423 410 427
rect 416 423 420 427
rect 426 423 430 427
rect 436 423 440 427
rect 446 423 450 427
rect 456 423 460 427
rect 466 423 470 427
rect 476 423 480 427
rect 486 423 490 427
rect 566 423 570 427
rect 566 413 570 417
rect 36 408 40 412
rect 46 408 50 412
rect 544 405 548 409
rect 554 405 558 409
rect 566 403 570 407
rect 298 392 302 396
rect 566 393 570 397
rect 566 383 570 387
rect 566 373 570 377
rect 36 368 40 372
rect 46 368 50 372
rect 298 362 302 366
rect 544 365 548 369
rect 554 365 558 369
rect 566 363 570 367
rect 114 356 118 360
rect 124 356 128 360
rect 134 356 138 360
rect 144 356 148 360
rect 154 356 158 360
rect 164 356 168 360
rect 174 356 178 360
rect 184 356 188 360
rect 194 356 198 360
rect 204 356 208 360
rect 214 356 218 360
rect 224 356 228 360
rect 234 356 238 360
rect 366 356 370 360
rect 376 356 380 360
rect 386 356 390 360
rect 396 356 400 360
rect 406 356 410 360
rect 416 356 420 360
rect 426 356 430 360
rect 436 356 440 360
rect 446 356 450 360
rect 456 356 460 360
rect 466 356 470 360
rect 476 356 480 360
rect 486 356 490 360
rect 566 353 570 357
rect 566 343 570 347
rect 298 332 302 336
rect 566 333 570 337
rect 36 328 40 332
rect 46 328 50 332
rect 132 328 136 332
rect 162 328 166 332
rect 192 328 196 332
rect 222 328 226 332
rect 385 329 389 333
rect 415 329 419 333
rect 445 329 449 333
rect 475 329 479 333
rect 544 325 548 329
rect 554 325 558 329
rect 566 323 570 327
rect 132 316 136 320
rect 162 316 166 320
rect 192 316 196 320
rect 222 316 226 320
rect 385 317 389 321
rect 415 317 419 321
rect 445 317 449 321
rect 475 317 479 321
rect 566 313 570 317
rect 298 302 302 306
rect 566 303 570 307
rect 36 288 40 292
rect 46 288 50 292
rect 112 290 116 294
rect 122 290 126 294
rect 132 290 136 294
rect 142 290 146 294
rect 152 290 156 294
rect 162 290 166 294
rect 172 290 176 294
rect 182 290 186 294
rect 192 290 196 294
rect 202 290 206 294
rect 212 290 216 294
rect 222 290 226 294
rect 232 290 236 294
rect 365 290 369 294
rect 375 290 379 294
rect 385 290 389 294
rect 395 290 399 294
rect 405 290 409 294
rect 415 290 419 294
rect 425 290 429 294
rect 435 290 439 294
rect 445 290 449 294
rect 455 290 459 294
rect 465 290 469 294
rect 475 290 479 294
rect 485 290 489 294
rect 566 293 570 297
rect 544 285 548 289
rect 554 285 558 289
rect 566 283 570 287
rect 298 272 302 276
rect 566 273 570 277
rect 566 263 570 267
rect 566 253 570 257
rect 36 248 40 252
rect 46 248 50 252
rect 298 242 302 246
rect 544 245 548 249
rect 554 245 558 249
rect 566 243 570 247
rect 566 233 570 237
rect 112 226 116 230
rect 122 226 126 230
rect 132 226 136 230
rect 142 226 146 230
rect 152 226 156 230
rect 162 226 166 230
rect 172 226 176 230
rect 182 226 186 230
rect 192 226 196 230
rect 202 226 206 230
rect 212 226 216 230
rect 222 226 226 230
rect 232 226 236 230
rect 366 225 370 229
rect 376 225 380 229
rect 386 225 390 229
rect 396 225 400 229
rect 406 225 410 229
rect 416 225 420 229
rect 426 225 430 229
rect 436 225 440 229
rect 446 225 450 229
rect 456 225 460 229
rect 466 225 470 229
rect 476 225 480 229
rect 486 225 490 229
rect 566 223 570 227
rect 298 212 302 216
rect 566 213 570 217
rect 36 208 40 212
rect 46 208 50 212
rect 544 205 548 209
rect 554 205 558 209
rect 566 203 570 207
rect 131 198 135 202
rect 161 198 165 202
rect 191 198 195 202
rect 221 198 225 202
rect 386 198 390 202
rect 416 198 420 202
rect 446 198 450 202
rect 476 198 480 202
rect 566 193 570 197
rect 131 186 135 190
rect 161 186 165 190
rect 191 186 195 190
rect 221 186 225 190
rect 386 186 390 190
rect 416 186 420 190
rect 446 186 450 190
rect 476 186 480 190
rect 298 182 302 186
rect 566 183 570 187
rect 566 173 570 177
rect 36 168 40 172
rect 46 168 50 172
rect 112 162 116 166
rect 122 162 126 166
rect 132 162 136 166
rect 142 162 146 166
rect 152 162 156 166
rect 162 162 166 166
rect 172 162 176 166
rect 182 162 186 166
rect 192 162 196 166
rect 202 162 206 166
rect 212 162 216 166
rect 222 162 226 166
rect 232 162 236 166
rect 366 162 370 166
rect 376 162 380 166
rect 386 162 390 166
rect 396 162 400 166
rect 406 162 410 166
rect 416 162 420 166
rect 426 162 430 166
rect 436 162 440 166
rect 446 162 450 166
rect 456 162 460 166
rect 466 162 470 166
rect 476 162 480 166
rect 486 162 490 166
rect 544 165 548 169
rect 554 165 558 169
rect 566 163 570 167
rect 298 152 302 156
rect 566 153 570 157
rect 566 143 570 147
rect 566 133 570 137
rect 36 128 40 132
rect 46 128 50 132
rect 298 122 302 126
rect 544 125 548 129
rect 554 125 558 129
rect 566 123 570 127
rect 566 113 570 117
rect 566 103 570 107
rect 110 96 114 100
rect 120 96 124 100
rect 130 96 134 100
rect 140 96 144 100
rect 150 96 154 100
rect 160 96 164 100
rect 170 96 174 100
rect 180 96 184 100
rect 190 96 194 100
rect 200 96 204 100
rect 210 96 214 100
rect 220 96 224 100
rect 230 96 234 100
rect 366 97 370 101
rect 376 97 380 101
rect 386 97 390 101
rect 396 97 400 101
rect 406 97 410 101
rect 416 97 420 101
rect 426 97 430 101
rect 436 97 440 101
rect 446 97 450 101
rect 456 97 460 101
rect 466 97 470 101
rect 476 97 480 101
rect 486 97 490 101
rect 566 93 570 97
rect 36 88 40 92
rect 46 88 50 92
rect 544 85 548 89
rect 554 85 558 89
rect 566 83 570 87
rect 566 73 570 77
rect 66 66 70 70
rect 530 67 534 71
rect 566 63 570 67
rect 120 56 124 60
rect 140 56 144 60
rect 160 56 164 60
rect 180 56 184 60
rect 200 56 204 60
rect 220 56 224 60
rect 376 56 380 60
rect 396 56 400 60
rect 416 56 420 60
rect 436 56 440 60
rect 456 56 460 60
rect 476 58 480 62
rect 566 53 570 57
rect 80 48 84 52
rect 120 46 124 50
rect 140 46 144 50
rect 160 46 164 50
rect 180 46 184 50
rect 200 46 204 50
rect 220 46 224 50
rect 376 46 380 50
rect 396 46 400 50
rect 416 46 420 50
rect 436 46 440 50
rect 456 46 460 50
rect 476 48 480 52
rect 36 42 40 46
rect 50 42 54 46
rect 60 42 64 46
rect 70 42 74 46
rect 538 42 542 46
rect 554 42 558 46
rect 566 43 570 47
rect 120 36 124 40
rect 140 36 144 40
rect 160 36 164 40
rect 180 36 184 40
rect 200 36 204 40
rect 220 36 224 40
rect 376 36 380 40
rect 396 36 400 40
rect 416 36 420 40
rect 436 36 440 40
rect 456 36 460 40
rect 476 38 480 42
rect 258 32 262 36
rect 268 32 272 36
rect 278 32 282 36
rect 288 32 292 36
rect 298 32 302 36
rect 308 32 312 36
rect 318 32 322 36
rect 328 32 332 36
rect 338 32 342 36
rect 566 33 570 37
rect 24 20 28 24
rect 34 20 38 24
rect 90 20 94 24
rect 100 20 104 24
rect 490 20 494 24
rect 500 20 504 24
rect 516 20 520 24
rect 526 20 530 24
<< end >>
