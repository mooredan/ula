magic
tech scmos
timestamp 1591539889
<< nwell >>
rect -1 29 29 81
<< nselect >>
rect 8 2 22 25
<< pselect >>
rect 8 33 22 77
<< ntransistor >>
rect 14 4 16 23
<< ptransistor >>
rect 14 35 16 75
<< ndiffusion >>
rect 10 4 14 23
rect 16 4 20 23
<< pdiffusion >>
rect 10 35 14 75
rect 16 35 20 75
<< polysilicon >>
rect 14 75 16 77
rect 14 33 16 35
rect 14 23 16 30
rect 14 2 16 4
<< metal1 >>
rect 5 76 23 79
rect 6 69 9 73
rect 19 69 22 73
rect 6 62 9 66
rect 19 62 22 66
rect 6 55 9 59
rect 19 55 22 59
rect 6 48 9 52
rect 19 48 22 52
rect 6 41 9 45
rect 19 41 22 45
rect 6 34 9 38
rect 19 34 22 38
rect 6 27 9 31
rect 19 27 22 31
rect 6 20 9 24
rect 19 20 22 24
rect 6 13 9 17
rect 19 13 22 17
rect 6 6 9 10
rect 19 6 22 10
rect 5 0 23 3
rect -2 -10 2 -3
rect 5 -10 9 -3
rect 12 -10 16 -3
rect 19 -10 23 -3
rect 26 -10 30 -3
<< bb >>
rect 0 0 28 79
<< labels >>
rlabel metal1 5 0 5 0 2 Gnd
port 3 ne
rlabel nwell 5 30 5 30 2 Vdd
rlabel metal1 5 76 5 76 2 Vdd
port 2 ne
<< end >>
