magic
tech amic5n
timestamp 1622292512
use inv_b  inv_b_0
timestamp 1622291139
transform 1 0 0 0 1 0
box -130 -45 580 1495
use inv_b  inv_b_1
timestamp 1622291139
transform 1 0 450 0 1 0
box -130 -45 580 1495
use inv_b  inv_b_5
timestamp 1622291139
transform 1 0 450 0 -1 2880
box -130 -45 580 1495
use inv_b  inv_b_4
timestamp 1622291139
transform 1 0 0 0 -1 2880
box -130 -45 580 1495
use inv_b  inv_b_2
timestamp 1622291139
transform -1 0 1350 0 1 0
box -130 -45 580 1495
use inv_b  inv_b_3
timestamp 1622291139
transform 1 0 1350 0 1 0
box -130 -45 580 1495
use inv_b  inv_b_7
timestamp 1622291139
transform 1 0 1350 0 -1 2880
box -130 -45 580 1495
use inv_b  inv_b_6
timestamp 1622291139
transform 1 0 900 0 -1 2880
box -130 -45 580 1495
use inv_b  inv_b_8
timestamp 1622291139
transform 1 0 0 0 1 2880
box -130 -45 580 1495
use inv_b  inv_b_9
timestamp 1622291139
transform 1 0 450 0 1 2880
box -130 -45 580 1495
use inv_b  inv_b_11
timestamp 1622291139
transform 1 0 1350 0 1 2880
box -130 -45 580 1495
use inv_b  inv_b_10
timestamp 1622291139
transform 1 0 900 0 1 2880
box -130 -45 580 1495
<< end >>
