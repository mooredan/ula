magic
tech amic5n
timestamp 1625354835
<< nwell >>
rect -130 550 580 1495
<< ntransistor >>
rect 165 95 285 400
<< ptransistor >>
rect 165 710 285 1345
<< nselect >>
rect -10 0 460 430
<< pselect >>
rect -10 680 460 1440
rect -10 670 165 680
rect 285 670 460 680
<< ndiffusion >>
rect 45 370 165 400
rect 45 320 75 370
rect 125 320 165 370
rect 45 175 165 320
rect 45 125 75 175
rect 125 125 165 175
rect 45 95 165 125
rect 285 355 405 400
rect 285 305 325 355
rect 375 305 405 355
rect 285 175 405 305
rect 285 125 325 175
rect 375 125 405 175
rect 285 95 405 125
<< pdiffusion >>
rect 45 1315 165 1345
rect 45 1265 75 1315
rect 125 1265 165 1315
rect 45 1190 165 1265
rect 45 1140 75 1190
rect 125 1140 165 1190
rect 45 1090 165 1140
rect 45 1040 75 1090
rect 125 1040 165 1090
rect 45 990 165 1040
rect 45 940 75 990
rect 125 940 165 990
rect 45 890 165 940
rect 45 840 75 890
rect 125 840 165 890
rect 45 710 165 840
rect 285 1315 405 1345
rect 285 1265 325 1315
rect 375 1265 405 1315
rect 285 1190 405 1265
rect 285 1140 325 1190
rect 375 1140 405 1190
rect 285 1090 405 1140
rect 285 1040 325 1090
rect 375 1040 405 1090
rect 285 990 405 1040
rect 285 940 325 990
rect 375 940 405 990
rect 285 890 405 940
rect 285 840 325 890
rect 375 840 405 890
rect 285 790 405 840
rect 285 740 325 790
rect 375 740 405 790
rect 285 710 405 740
<< ndcontact >>
rect 75 320 125 370
rect 75 125 125 175
rect 325 305 375 355
rect 325 125 375 175
<< pdcontact >>
rect 75 1265 125 1315
rect 75 1140 125 1190
rect 75 1040 125 1090
rect 75 940 125 990
rect 75 840 125 890
rect 325 1265 375 1315
rect 325 1140 375 1190
rect 325 1040 375 1090
rect 325 940 375 990
rect 325 840 375 890
rect 325 740 375 790
<< polysilicon >>
rect 165 1345 285 1410
rect 165 675 285 710
rect 55 655 285 675
rect 55 605 75 655
rect 125 605 175 655
rect 225 605 285 655
rect 55 585 285 605
rect 165 505 395 525
rect 165 455 225 505
rect 275 455 325 505
rect 375 455 395 505
rect 165 435 395 455
rect 165 400 285 435
rect 165 30 285 95
<< polycontact >>
rect 75 605 125 655
rect 175 605 225 655
rect 225 455 275 505
rect 325 455 375 505
<< metal1 >>
rect 0 1395 450 1485
rect 55 1315 145 1395
rect 55 1265 75 1315
rect 125 1265 145 1315
rect 55 1190 145 1265
rect 55 1140 75 1190
rect 125 1140 145 1190
rect 55 1090 145 1140
rect 55 1040 75 1090
rect 125 1040 145 1090
rect 55 990 145 1040
rect 55 940 75 990
rect 125 940 145 990
rect 55 890 145 940
rect 55 840 75 890
rect 125 840 145 890
rect 55 735 145 840
rect 305 1315 395 1395
rect 305 1265 325 1315
rect 375 1265 395 1315
rect 305 1190 395 1265
rect 305 1140 325 1190
rect 375 1140 395 1190
rect 305 1090 395 1140
rect 305 1040 325 1090
rect 375 1040 395 1090
rect 305 990 395 1040
rect 305 940 325 990
rect 375 940 395 990
rect 305 890 395 940
rect 305 840 325 890
rect 375 840 395 890
rect 305 790 395 840
rect 305 740 325 790
rect 375 740 395 790
rect 55 655 245 675
rect 55 605 75 655
rect 125 605 175 655
rect 225 605 245 655
rect 55 585 245 605
rect 55 370 145 585
rect 305 525 395 740
rect 205 505 395 525
rect 205 455 225 505
rect 275 455 325 505
rect 375 455 395 505
rect 205 435 395 455
rect 55 320 75 370
rect 125 320 145 370
rect 55 175 145 320
rect 55 125 75 175
rect 125 125 145 175
rect 55 45 145 125
rect 305 355 395 375
rect 305 305 325 355
rect 375 305 395 355
rect 305 175 395 305
rect 305 125 325 175
rect 375 125 395 175
rect 305 45 395 125
rect 0 -45 450 45
<< labels >>
flabel metal1 s 5 5 5 5 2 FreeSans 400 0 0 0 vss
port 1 ne
flabel metal1 s 20 1415 20 1415 2 FreeSans 400 0 0 0 vdd
port 0 ne
flabel nwell 5 600 5 600 2 FreeSans 400 0 0 0 vdd
<< properties >>
string LEFsite core
string LEFclass CORE
string FIXED_BBOX 0 0 450 1440
string LEFsymmetry X Y
<< end >>
