magic
tech scmos
timestamp 1594330712
<< nwell >>
rect 14 452 346 681
rect -3 418 363 435
rect -3 373 363 390
rect -3 144 14 373
rect 346 144 363 373
rect -3 127 363 144
<< nselect >>
rect 22 13 74 94
rect 286 13 338 94
<< pselect >>
rect -2 111 362 126
rect -2 13 13 111
rect 347 13 362 111
rect -2 -2 362 13
<< ntransistor >>
rect 45 344 159 347
rect 45 300 159 303
rect 45 279 159 282
rect 45 235 159 238
rect 45 214 159 217
rect 45 170 159 173
rect 201 344 315 347
rect 201 300 315 303
rect 201 279 315 282
rect 201 235 315 238
rect 201 214 315 217
rect 201 170 315 173
rect 29 84 72 86
rect 288 84 331 86
rect 29 76 72 78
rect 288 76 331 78
rect 29 68 72 70
rect 29 60 72 62
rect 29 52 72 54
rect 288 68 331 70
rect 288 60 331 62
rect 288 52 331 54
rect 29 44 72 46
rect 29 36 72 38
rect 288 44 331 46
rect 288 36 331 38
rect 29 28 72 30
rect 29 20 72 22
rect 288 28 331 30
rect 288 20 331 22
<< ptransistor >>
rect 38 652 166 655
rect 38 608 166 611
rect 38 587 166 590
rect 38 543 166 546
rect 38 522 166 525
rect 38 478 166 481
rect 194 652 322 655
rect 194 608 322 611
rect 194 587 322 590
rect 194 543 322 546
rect 194 522 322 525
rect 194 478 322 481
<< ndiffusion >>
rect 43 350 161 356
rect 199 350 317 356
rect 45 347 159 350
rect 45 303 159 344
rect 45 282 159 300
rect 45 238 159 279
rect 45 217 159 235
rect 45 173 159 214
rect 45 167 159 170
rect 201 347 315 350
rect 201 303 315 344
rect 201 282 315 300
rect 201 238 315 279
rect 201 217 315 235
rect 201 173 315 214
rect 201 167 315 170
rect 43 161 161 167
rect 199 161 317 167
rect 29 86 72 92
rect 288 86 331 92
rect 29 78 72 84
rect 29 70 72 76
rect 288 78 331 84
rect 29 62 72 68
rect 29 54 72 60
rect 29 46 72 52
rect 288 70 331 76
rect 288 62 331 68
rect 288 54 331 60
rect 29 38 72 44
rect 288 46 331 52
rect 288 38 331 44
rect 29 30 72 36
rect 29 22 72 28
rect 288 30 331 36
rect 288 22 331 28
rect 29 15 72 20
rect 288 15 331 20
<< pdiffusion >>
rect 36 658 168 664
rect 192 658 324 664
rect 38 655 166 658
rect 38 611 166 652
rect 38 590 166 608
rect 38 546 166 587
rect 38 525 166 543
rect 38 481 166 522
rect 38 475 166 478
rect 194 655 322 658
rect 194 611 322 652
rect 194 590 322 608
rect 194 546 322 587
rect 194 525 322 543
rect 194 481 322 522
rect 194 475 322 478
rect 36 469 168 475
rect 192 469 324 475
<< psubstratepdiff >>
rect 0 684 360 695
rect 0 449 11 684
rect 349 449 360 684
rect 0 438 360 449
rect 0 393 360 404
rect 19 356 341 368
rect 19 350 43 356
rect 161 350 199 356
rect 317 350 341 356
rect 19 167 37 350
rect 167 167 193 350
rect 323 167 341 350
rect 19 161 43 167
rect 161 161 199 167
rect 317 161 341 167
rect 19 149 341 161
rect 0 113 360 124
rect 0 11 11 113
rect 349 11 360 113
rect 0 0 360 11
<< nsubstratendiff >>
rect 19 664 341 676
rect 19 658 36 664
rect 168 658 192 664
rect 324 658 341 664
rect 19 475 30 658
rect 174 475 186 658
rect 330 475 341 658
rect 19 469 36 475
rect 168 469 192 475
rect 324 469 341 475
rect 19 457 341 469
rect 0 421 360 432
rect 0 376 360 387
rect 0 141 11 376
rect 349 141 360 376
rect 0 130 360 141
rect 81 71 279 82
rect 81 36 279 47
<< polysilicon >>
rect 31 652 38 655
rect 166 652 173 655
rect 31 611 37 652
rect 167 611 173 652
rect 31 608 38 611
rect 166 608 173 611
rect 31 590 37 608
rect 167 590 173 608
rect 31 587 38 590
rect 166 587 173 590
rect 31 546 37 587
rect 167 546 173 587
rect 31 543 38 546
rect 166 543 173 546
rect 31 525 37 543
rect 167 525 173 543
rect 31 522 38 525
rect 166 522 173 525
rect 31 481 37 522
rect 167 481 173 522
rect 31 478 38 481
rect 166 478 173 481
rect 187 652 194 655
rect 322 652 329 655
rect 187 611 193 652
rect 323 611 329 652
rect 187 608 194 611
rect 322 608 329 611
rect 187 590 193 608
rect 323 590 329 608
rect 187 587 194 590
rect 322 587 329 590
rect 187 546 193 587
rect 323 546 329 587
rect 187 543 194 546
rect 322 543 329 546
rect 187 525 193 543
rect 323 525 329 543
rect 187 522 194 525
rect 322 522 329 525
rect 187 481 193 522
rect 323 481 329 522
rect 187 478 194 481
rect 322 478 329 481
rect 38 344 45 347
rect 159 344 166 347
rect 38 303 44 344
rect 160 303 166 344
rect 38 300 45 303
rect 159 300 166 303
rect 38 282 44 300
rect 160 282 166 300
rect 38 279 45 282
rect 159 279 166 282
rect 38 238 44 279
rect 160 238 166 279
rect 38 235 45 238
rect 159 235 166 238
rect 38 228 44 235
rect 38 217 44 221
rect 160 228 166 235
rect 160 217 166 221
rect 38 214 45 217
rect 159 214 166 217
rect 38 173 44 214
rect 160 173 166 214
rect 38 170 45 173
rect 159 170 166 173
rect 194 344 201 347
rect 315 344 322 347
rect 194 303 200 344
rect 316 303 322 344
rect 194 300 201 303
rect 315 300 322 303
rect 194 282 200 300
rect 316 282 322 300
rect 194 279 201 282
rect 315 279 322 282
rect 194 264 200 279
rect 194 238 200 256
rect 316 264 322 279
rect 316 238 322 256
rect 194 235 201 238
rect 315 235 322 238
rect 194 217 200 235
rect 316 217 322 235
rect 194 214 201 217
rect 315 214 322 217
rect 194 173 200 214
rect 316 173 322 214
rect 194 170 201 173
rect 315 170 322 173
rect 22 84 29 86
rect 72 84 76 86
rect 22 78 28 84
rect 74 78 76 84
rect 284 84 288 86
rect 331 84 338 86
rect 22 76 29 78
rect 72 76 76 78
rect 22 70 28 76
rect 74 70 76 76
rect 284 78 286 84
rect 332 78 338 84
rect 284 76 288 78
rect 331 76 338 78
rect 22 68 29 70
rect 72 68 76 70
rect 22 62 28 68
rect 74 62 76 68
rect 22 60 29 62
rect 72 60 76 62
rect 22 54 28 60
rect 74 54 76 60
rect 22 52 29 54
rect 72 52 76 54
rect 22 46 28 52
rect 74 46 76 52
rect 284 70 286 76
rect 332 70 338 76
rect 284 68 288 70
rect 331 68 338 70
rect 284 62 286 68
rect 332 62 338 68
rect 284 60 288 62
rect 331 60 338 62
rect 284 54 286 60
rect 332 54 338 60
rect 284 52 288 54
rect 331 52 338 54
rect 22 44 29 46
rect 72 44 76 46
rect 22 38 28 44
rect 74 38 76 44
rect 22 36 29 38
rect 72 36 76 38
rect 284 46 286 52
rect 332 46 338 52
rect 284 44 288 46
rect 331 44 338 46
rect 284 38 286 44
rect 332 38 338 44
rect 284 36 288 38
rect 331 36 338 38
rect 22 30 28 36
rect 74 30 76 36
rect 22 28 29 30
rect 72 28 76 30
rect 22 22 28 28
rect 74 22 76 28
rect 22 20 29 22
rect 72 20 76 22
rect 284 30 286 36
rect 332 30 338 36
rect 284 28 288 30
rect 331 28 338 30
rect 284 22 286 28
rect 332 22 338 28
rect 284 20 288 22
rect 331 20 338 22
rect 22 15 28 20
rect 332 15 338 20
<< genericcontact >>
rect 9 691 11 693
rect 17 691 19 693
rect 25 691 27 693
rect 33 691 35 693
rect 41 691 43 693
rect 49 691 51 693
rect 57 691 59 693
rect 65 691 67 693
rect 73 691 75 693
rect 81 691 83 693
rect 89 691 91 693
rect 97 691 99 693
rect 105 691 107 693
rect 113 691 115 693
rect 151 691 153 693
rect 159 691 161 693
rect 167 691 169 693
rect 175 691 177 693
rect 183 691 185 693
rect 191 691 193 693
rect 199 691 201 693
rect 207 691 209 693
rect 245 691 247 693
rect 253 691 255 693
rect 261 691 263 693
rect 269 691 271 693
rect 277 691 279 693
rect 285 691 287 693
rect 293 691 295 693
rect 301 691 303 693
rect 309 691 311 693
rect 317 691 319 693
rect 325 691 327 693
rect 333 691 335 693
rect 341 691 343 693
rect 349 691 351 693
rect 9 686 11 688
rect 17 686 19 688
rect 25 686 27 688
rect 33 686 35 688
rect 41 686 43 688
rect 49 686 51 688
rect 57 686 59 688
rect 65 686 67 688
rect 73 686 75 688
rect 81 686 83 688
rect 89 686 91 688
rect 97 686 99 688
rect 105 686 107 688
rect 113 686 115 688
rect 151 686 153 688
rect 159 686 161 688
rect 167 686 169 688
rect 175 686 177 688
rect 183 686 185 688
rect 191 686 193 688
rect 199 686 201 688
rect 207 686 209 688
rect 245 686 247 688
rect 253 686 255 688
rect 261 686 263 688
rect 269 686 271 688
rect 277 686 279 688
rect 285 686 287 688
rect 293 686 295 688
rect 301 686 303 688
rect 309 686 311 688
rect 317 686 319 688
rect 325 686 327 688
rect 333 686 335 688
rect 341 686 343 688
rect 349 686 351 688
rect 2 678 4 680
rect 7 678 9 680
rect 351 678 353 680
rect 356 678 358 680
rect 2 670 4 672
rect 7 670 9 672
rect 351 670 353 672
rect 356 670 358 672
rect 30 668 32 670
rect 41 668 43 670
rect 51 668 53 670
rect 61 668 63 670
rect 71 668 73 670
rect 81 668 83 670
rect 91 668 93 670
rect 101 668 103 670
rect 111 668 113 670
rect 150 668 152 670
rect 160 668 162 670
rect 198 668 200 670
rect 208 668 210 670
rect 247 668 249 670
rect 257 668 259 670
rect 267 668 269 670
rect 277 668 279 670
rect 287 668 289 670
rect 297 668 299 670
rect 307 668 309 670
rect 317 668 319 670
rect 327 668 329 670
rect 2 662 4 664
rect 7 662 9 664
rect 30 663 32 665
rect 41 663 43 665
rect 51 663 53 665
rect 61 663 63 665
rect 71 663 73 665
rect 81 663 83 665
rect 91 663 93 665
rect 101 663 103 665
rect 111 663 113 665
rect 150 663 152 665
rect 160 663 162 665
rect 198 663 200 665
rect 208 663 210 665
rect 247 663 249 665
rect 257 663 259 665
rect 267 663 269 665
rect 277 663 279 665
rect 287 663 289 665
rect 297 663 299 665
rect 307 663 309 665
rect 317 663 319 665
rect 327 663 329 665
rect 351 662 353 664
rect 356 662 358 664
rect 41 658 43 660
rect 51 658 53 660
rect 61 658 63 660
rect 71 658 73 660
rect 81 658 83 660
rect 91 658 93 660
rect 101 658 103 660
rect 111 658 113 660
rect 150 658 152 660
rect 160 658 162 660
rect 198 658 200 660
rect 208 658 210 660
rect 247 658 249 660
rect 257 658 259 660
rect 267 658 269 660
rect 277 658 279 660
rect 287 658 289 660
rect 297 658 299 660
rect 307 658 309 660
rect 317 658 319 660
rect 2 654 4 656
rect 7 654 9 656
rect 20 653 22 655
rect 25 653 27 655
rect 177 653 179 655
rect 182 653 184 655
rect 333 653 335 655
rect 338 653 340 655
rect 351 654 353 656
rect 356 654 358 656
rect 33 650 35 652
rect 169 650 171 652
rect 189 650 191 652
rect 325 650 327 652
rect 20 648 22 650
rect 25 648 27 650
rect 42 648 44 650
rect 47 648 49 650
rect 52 648 54 650
rect 57 648 59 650
rect 62 648 64 650
rect 67 648 69 650
rect 72 648 74 650
rect 77 648 79 650
rect 82 648 84 650
rect 87 648 89 650
rect 92 648 94 650
rect 97 648 99 650
rect 102 648 104 650
rect 107 648 109 650
rect 112 648 114 650
rect 117 648 119 650
rect 122 648 124 650
rect 127 648 129 650
rect 132 648 134 650
rect 137 648 139 650
rect 142 648 144 650
rect 147 648 149 650
rect 152 648 154 650
rect 157 648 159 650
rect 162 648 164 650
rect 177 648 179 650
rect 182 648 184 650
rect 196 648 198 650
rect 201 648 203 650
rect 206 648 208 650
rect 211 648 213 650
rect 216 648 218 650
rect 221 648 223 650
rect 226 648 228 650
rect 231 648 233 650
rect 236 648 238 650
rect 241 648 243 650
rect 246 648 248 650
rect 251 648 253 650
rect 256 648 258 650
rect 261 648 263 650
rect 266 648 268 650
rect 271 648 273 650
rect 276 648 278 650
rect 281 648 283 650
rect 286 648 288 650
rect 291 648 293 650
rect 296 648 298 650
rect 301 648 303 650
rect 306 648 308 650
rect 311 648 313 650
rect 316 648 318 650
rect 333 648 335 650
rect 338 648 340 650
rect 2 646 4 648
rect 7 646 9 648
rect 33 645 35 647
rect 169 645 171 647
rect 189 645 191 647
rect 325 645 327 647
rect 351 646 353 648
rect 356 646 358 648
rect 20 643 22 645
rect 25 643 27 645
rect 42 643 44 645
rect 47 643 49 645
rect 52 643 54 645
rect 57 643 59 645
rect 62 643 64 645
rect 67 643 69 645
rect 72 643 74 645
rect 77 643 79 645
rect 82 643 84 645
rect 87 643 89 645
rect 92 643 94 645
rect 97 643 99 645
rect 102 643 104 645
rect 107 643 109 645
rect 112 643 114 645
rect 117 643 119 645
rect 122 643 124 645
rect 127 643 129 645
rect 132 643 134 645
rect 137 643 139 645
rect 142 643 144 645
rect 147 643 149 645
rect 152 643 154 645
rect 157 643 159 645
rect 162 643 164 645
rect 177 643 179 645
rect 182 643 184 645
rect 196 643 198 645
rect 201 643 203 645
rect 206 643 208 645
rect 211 643 213 645
rect 216 643 218 645
rect 221 643 223 645
rect 226 643 228 645
rect 231 643 233 645
rect 236 643 238 645
rect 241 643 243 645
rect 246 643 248 645
rect 251 643 253 645
rect 256 643 258 645
rect 261 643 263 645
rect 266 643 268 645
rect 271 643 273 645
rect 276 643 278 645
rect 281 643 283 645
rect 286 643 288 645
rect 291 643 293 645
rect 296 643 298 645
rect 301 643 303 645
rect 306 643 308 645
rect 311 643 313 645
rect 316 643 318 645
rect 333 643 335 645
rect 338 643 340 645
rect 33 640 35 642
rect 169 640 171 642
rect 189 640 191 642
rect 325 640 327 642
rect 2 638 4 640
rect 7 638 9 640
rect 20 638 22 640
rect 25 638 27 640
rect 42 638 44 640
rect 47 638 49 640
rect 52 638 54 640
rect 57 638 59 640
rect 62 638 64 640
rect 67 638 69 640
rect 72 638 74 640
rect 77 638 79 640
rect 82 638 84 640
rect 87 638 89 640
rect 92 638 94 640
rect 97 638 99 640
rect 102 638 104 640
rect 107 638 109 640
rect 112 638 114 640
rect 117 638 119 640
rect 122 638 124 640
rect 127 638 129 640
rect 132 638 134 640
rect 137 638 139 640
rect 142 638 144 640
rect 147 638 149 640
rect 152 638 154 640
rect 157 638 159 640
rect 162 638 164 640
rect 177 638 179 640
rect 182 638 184 640
rect 196 638 198 640
rect 201 638 203 640
rect 206 638 208 640
rect 211 638 213 640
rect 216 638 218 640
rect 221 638 223 640
rect 226 638 228 640
rect 231 638 233 640
rect 236 638 238 640
rect 241 638 243 640
rect 246 638 248 640
rect 251 638 253 640
rect 256 638 258 640
rect 261 638 263 640
rect 266 638 268 640
rect 271 638 273 640
rect 276 638 278 640
rect 281 638 283 640
rect 286 638 288 640
rect 291 638 293 640
rect 296 638 298 640
rect 301 638 303 640
rect 306 638 308 640
rect 311 638 313 640
rect 316 638 318 640
rect 333 638 335 640
rect 338 638 340 640
rect 351 638 353 640
rect 356 638 358 640
rect 33 635 35 637
rect 169 635 171 637
rect 189 635 191 637
rect 325 635 327 637
rect 20 633 22 635
rect 25 633 27 635
rect 42 633 44 635
rect 47 633 49 635
rect 52 633 54 635
rect 57 633 59 635
rect 62 633 64 635
rect 67 633 69 635
rect 72 633 74 635
rect 77 633 79 635
rect 82 633 84 635
rect 87 633 89 635
rect 92 633 94 635
rect 97 633 99 635
rect 102 633 104 635
rect 107 633 109 635
rect 112 633 114 635
rect 117 633 119 635
rect 122 633 124 635
rect 127 633 129 635
rect 132 633 134 635
rect 137 633 139 635
rect 142 633 144 635
rect 147 633 149 635
rect 152 633 154 635
rect 157 633 159 635
rect 162 633 164 635
rect 177 633 179 635
rect 182 633 184 635
rect 196 633 198 635
rect 201 633 203 635
rect 206 633 208 635
rect 211 633 213 635
rect 216 633 218 635
rect 221 633 223 635
rect 226 633 228 635
rect 231 633 233 635
rect 236 633 238 635
rect 241 633 243 635
rect 246 633 248 635
rect 251 633 253 635
rect 256 633 258 635
rect 261 633 263 635
rect 266 633 268 635
rect 271 633 273 635
rect 276 633 278 635
rect 281 633 283 635
rect 286 633 288 635
rect 291 633 293 635
rect 296 633 298 635
rect 301 633 303 635
rect 306 633 308 635
rect 311 633 313 635
rect 316 633 318 635
rect 333 633 335 635
rect 338 633 340 635
rect 2 630 4 632
rect 7 630 9 632
rect 33 630 35 632
rect 169 630 171 632
rect 189 630 191 632
rect 325 630 327 632
rect 351 630 353 632
rect 356 630 358 632
rect 20 628 22 630
rect 25 628 27 630
rect 42 628 44 630
rect 47 628 49 630
rect 52 628 54 630
rect 57 628 59 630
rect 62 628 64 630
rect 67 628 69 630
rect 72 628 74 630
rect 77 628 79 630
rect 82 628 84 630
rect 87 628 89 630
rect 92 628 94 630
rect 97 628 99 630
rect 102 628 104 630
rect 107 628 109 630
rect 112 628 114 630
rect 117 628 119 630
rect 122 628 124 630
rect 127 628 129 630
rect 132 628 134 630
rect 137 628 139 630
rect 142 628 144 630
rect 147 628 149 630
rect 152 628 154 630
rect 157 628 159 630
rect 162 628 164 630
rect 177 628 179 630
rect 182 628 184 630
rect 196 628 198 630
rect 201 628 203 630
rect 206 628 208 630
rect 211 628 213 630
rect 216 628 218 630
rect 221 628 223 630
rect 226 628 228 630
rect 231 628 233 630
rect 236 628 238 630
rect 241 628 243 630
rect 246 628 248 630
rect 251 628 253 630
rect 256 628 258 630
rect 261 628 263 630
rect 266 628 268 630
rect 271 628 273 630
rect 276 628 278 630
rect 281 628 283 630
rect 286 628 288 630
rect 291 628 293 630
rect 296 628 298 630
rect 301 628 303 630
rect 306 628 308 630
rect 311 628 313 630
rect 316 628 318 630
rect 333 628 335 630
rect 338 628 340 630
rect 33 625 35 627
rect 169 625 171 627
rect 189 625 191 627
rect 325 625 327 627
rect 2 622 4 624
rect 7 622 9 624
rect 20 623 22 625
rect 25 623 27 625
rect 42 623 44 625
rect 47 623 49 625
rect 52 623 54 625
rect 57 623 59 625
rect 62 623 64 625
rect 67 623 69 625
rect 72 623 74 625
rect 77 623 79 625
rect 82 623 84 625
rect 87 623 89 625
rect 92 623 94 625
rect 97 623 99 625
rect 102 623 104 625
rect 107 623 109 625
rect 112 623 114 625
rect 117 623 119 625
rect 122 623 124 625
rect 127 623 129 625
rect 132 623 134 625
rect 137 623 139 625
rect 142 623 144 625
rect 147 623 149 625
rect 152 623 154 625
rect 157 623 159 625
rect 162 623 164 625
rect 177 623 179 625
rect 182 623 184 625
rect 196 623 198 625
rect 201 623 203 625
rect 206 623 208 625
rect 211 623 213 625
rect 216 623 218 625
rect 221 623 223 625
rect 226 623 228 625
rect 231 623 233 625
rect 236 623 238 625
rect 241 623 243 625
rect 246 623 248 625
rect 251 623 253 625
rect 256 623 258 625
rect 261 623 263 625
rect 266 623 268 625
rect 271 623 273 625
rect 276 623 278 625
rect 281 623 283 625
rect 286 623 288 625
rect 291 623 293 625
rect 296 623 298 625
rect 301 623 303 625
rect 306 623 308 625
rect 311 623 313 625
rect 316 623 318 625
rect 333 623 335 625
rect 338 623 340 625
rect 351 622 353 624
rect 356 622 358 624
rect 33 620 35 622
rect 169 620 171 622
rect 189 620 191 622
rect 325 620 327 622
rect 20 618 22 620
rect 25 618 27 620
rect 42 618 44 620
rect 47 618 49 620
rect 52 618 54 620
rect 57 618 59 620
rect 62 618 64 620
rect 67 618 69 620
rect 72 618 74 620
rect 77 618 79 620
rect 82 618 84 620
rect 87 618 89 620
rect 92 618 94 620
rect 97 618 99 620
rect 102 618 104 620
rect 107 618 109 620
rect 112 618 114 620
rect 117 618 119 620
rect 122 618 124 620
rect 127 618 129 620
rect 132 618 134 620
rect 137 618 139 620
rect 142 618 144 620
rect 147 618 149 620
rect 152 618 154 620
rect 157 618 159 620
rect 162 618 164 620
rect 177 618 179 620
rect 182 618 184 620
rect 196 618 198 620
rect 201 618 203 620
rect 206 618 208 620
rect 211 618 213 620
rect 216 618 218 620
rect 221 618 223 620
rect 226 618 228 620
rect 231 618 233 620
rect 236 618 238 620
rect 241 618 243 620
rect 246 618 248 620
rect 251 618 253 620
rect 256 618 258 620
rect 261 618 263 620
rect 266 618 268 620
rect 271 618 273 620
rect 276 618 278 620
rect 281 618 283 620
rect 286 618 288 620
rect 291 618 293 620
rect 296 618 298 620
rect 301 618 303 620
rect 306 618 308 620
rect 311 618 313 620
rect 316 618 318 620
rect 333 618 335 620
rect 338 618 340 620
rect 2 614 4 616
rect 7 614 9 616
rect 33 615 35 617
rect 169 615 171 617
rect 189 615 191 617
rect 325 615 327 617
rect 20 613 22 615
rect 25 613 27 615
rect 42 613 44 615
rect 47 613 49 615
rect 52 613 54 615
rect 57 613 59 615
rect 62 613 64 615
rect 67 613 69 615
rect 72 613 74 615
rect 77 613 79 615
rect 82 613 84 615
rect 87 613 89 615
rect 92 613 94 615
rect 97 613 99 615
rect 102 613 104 615
rect 107 613 109 615
rect 112 613 114 615
rect 117 613 119 615
rect 122 613 124 615
rect 127 613 129 615
rect 132 613 134 615
rect 137 613 139 615
rect 142 613 144 615
rect 147 613 149 615
rect 152 613 154 615
rect 157 613 159 615
rect 162 613 164 615
rect 177 613 179 615
rect 182 613 184 615
rect 196 613 198 615
rect 201 613 203 615
rect 206 613 208 615
rect 211 613 213 615
rect 216 613 218 615
rect 221 613 223 615
rect 226 613 228 615
rect 231 613 233 615
rect 236 613 238 615
rect 241 613 243 615
rect 246 613 248 615
rect 251 613 253 615
rect 256 613 258 615
rect 261 613 263 615
rect 266 613 268 615
rect 271 613 273 615
rect 276 613 278 615
rect 281 613 283 615
rect 286 613 288 615
rect 291 613 293 615
rect 296 613 298 615
rect 301 613 303 615
rect 306 613 308 615
rect 311 613 313 615
rect 316 613 318 615
rect 333 613 335 615
rect 338 613 340 615
rect 351 614 353 616
rect 356 614 358 616
rect 33 610 35 612
rect 169 610 171 612
rect 189 610 191 612
rect 325 610 327 612
rect 20 608 22 610
rect 25 608 27 610
rect 177 608 179 610
rect 182 608 184 610
rect 333 608 335 610
rect 338 608 340 610
rect 2 606 4 608
rect 7 606 9 608
rect 33 605 35 607
rect 169 605 171 607
rect 189 605 191 607
rect 325 605 327 607
rect 351 606 353 608
rect 356 606 358 608
rect 41 603 43 605
rect 51 603 53 605
rect 61 603 63 605
rect 71 603 73 605
rect 81 603 83 605
rect 91 603 93 605
rect 101 603 103 605
rect 111 603 113 605
rect 150 603 152 605
rect 160 603 162 605
rect 198 603 200 605
rect 208 603 210 605
rect 247 603 249 605
rect 257 603 259 605
rect 267 603 269 605
rect 277 603 279 605
rect 287 603 289 605
rect 297 603 299 605
rect 307 603 309 605
rect 317 603 319 605
rect 33 600 35 602
rect 169 600 171 602
rect 189 600 191 602
rect 325 600 327 602
rect 2 598 4 600
rect 7 598 9 600
rect 41 598 43 600
rect 51 598 53 600
rect 61 598 63 600
rect 71 598 73 600
rect 81 598 83 600
rect 91 598 93 600
rect 101 598 103 600
rect 111 598 113 600
rect 150 598 152 600
rect 160 598 162 600
rect 198 598 200 600
rect 208 598 210 600
rect 247 598 249 600
rect 257 598 259 600
rect 267 598 269 600
rect 277 598 279 600
rect 287 598 289 600
rect 297 598 299 600
rect 307 598 309 600
rect 317 598 319 600
rect 351 598 353 600
rect 356 598 358 600
rect 33 595 35 597
rect 169 595 171 597
rect 189 595 191 597
rect 325 595 327 597
rect 41 593 43 595
rect 51 593 53 595
rect 61 593 63 595
rect 71 593 73 595
rect 81 593 83 595
rect 91 593 93 595
rect 101 593 103 595
rect 111 593 113 595
rect 150 593 152 595
rect 160 593 162 595
rect 198 593 200 595
rect 208 593 210 595
rect 247 593 249 595
rect 257 593 259 595
rect 267 593 269 595
rect 277 593 279 595
rect 287 593 289 595
rect 297 593 299 595
rect 307 593 309 595
rect 317 593 319 595
rect 2 590 4 592
rect 7 590 9 592
rect 33 590 35 592
rect 169 590 171 592
rect 189 590 191 592
rect 325 590 327 592
rect 351 590 353 592
rect 356 590 358 592
rect 20 588 22 590
rect 25 588 27 590
rect 177 588 179 590
rect 182 588 184 590
rect 333 588 335 590
rect 338 588 340 590
rect 33 585 35 587
rect 169 585 171 587
rect 189 585 191 587
rect 325 585 327 587
rect 2 582 4 584
rect 7 582 9 584
rect 20 583 22 585
rect 25 583 27 585
rect 42 583 44 585
rect 47 583 49 585
rect 52 583 54 585
rect 57 583 59 585
rect 62 583 64 585
rect 67 583 69 585
rect 72 583 74 585
rect 77 583 79 585
rect 82 583 84 585
rect 87 583 89 585
rect 92 583 94 585
rect 97 583 99 585
rect 102 583 104 585
rect 107 583 109 585
rect 112 583 114 585
rect 117 583 119 585
rect 122 583 124 585
rect 127 583 129 585
rect 132 583 134 585
rect 137 583 139 585
rect 142 583 144 585
rect 147 583 149 585
rect 152 583 154 585
rect 157 583 159 585
rect 162 583 164 585
rect 177 583 179 585
rect 182 583 184 585
rect 196 583 198 585
rect 201 583 203 585
rect 206 583 208 585
rect 211 583 213 585
rect 216 583 218 585
rect 221 583 223 585
rect 226 583 228 585
rect 231 583 233 585
rect 236 583 238 585
rect 241 583 243 585
rect 246 583 248 585
rect 251 583 253 585
rect 256 583 258 585
rect 261 583 263 585
rect 266 583 268 585
rect 271 583 273 585
rect 276 583 278 585
rect 281 583 283 585
rect 286 583 288 585
rect 291 583 293 585
rect 296 583 298 585
rect 301 583 303 585
rect 306 583 308 585
rect 311 583 313 585
rect 316 583 318 585
rect 333 583 335 585
rect 338 583 340 585
rect 351 582 353 584
rect 356 582 358 584
rect 33 580 35 582
rect 169 580 171 582
rect 189 580 191 582
rect 325 580 327 582
rect 20 578 22 580
rect 25 578 27 580
rect 42 578 44 580
rect 47 578 49 580
rect 52 578 54 580
rect 57 578 59 580
rect 62 578 64 580
rect 67 578 69 580
rect 72 578 74 580
rect 77 578 79 580
rect 82 578 84 580
rect 87 578 89 580
rect 92 578 94 580
rect 97 578 99 580
rect 102 578 104 580
rect 107 578 109 580
rect 112 578 114 580
rect 117 578 119 580
rect 122 578 124 580
rect 127 578 129 580
rect 132 578 134 580
rect 137 578 139 580
rect 142 578 144 580
rect 147 578 149 580
rect 152 578 154 580
rect 157 578 159 580
rect 162 578 164 580
rect 177 578 179 580
rect 182 578 184 580
rect 196 578 198 580
rect 201 578 203 580
rect 206 578 208 580
rect 211 578 213 580
rect 216 578 218 580
rect 221 578 223 580
rect 226 578 228 580
rect 231 578 233 580
rect 236 578 238 580
rect 241 578 243 580
rect 246 578 248 580
rect 251 578 253 580
rect 256 578 258 580
rect 261 578 263 580
rect 266 578 268 580
rect 271 578 273 580
rect 276 578 278 580
rect 281 578 283 580
rect 286 578 288 580
rect 291 578 293 580
rect 296 578 298 580
rect 301 578 303 580
rect 306 578 308 580
rect 311 578 313 580
rect 316 578 318 580
rect 333 578 335 580
rect 338 578 340 580
rect 2 574 4 576
rect 7 574 9 576
rect 33 575 35 577
rect 169 575 171 577
rect 189 575 191 577
rect 325 575 327 577
rect 20 573 22 575
rect 25 573 27 575
rect 42 573 44 575
rect 47 573 49 575
rect 52 573 54 575
rect 57 573 59 575
rect 62 573 64 575
rect 67 573 69 575
rect 72 573 74 575
rect 77 573 79 575
rect 82 573 84 575
rect 87 573 89 575
rect 92 573 94 575
rect 97 573 99 575
rect 102 573 104 575
rect 107 573 109 575
rect 112 573 114 575
rect 117 573 119 575
rect 122 573 124 575
rect 127 573 129 575
rect 132 573 134 575
rect 137 573 139 575
rect 142 573 144 575
rect 147 573 149 575
rect 152 573 154 575
rect 157 573 159 575
rect 162 573 164 575
rect 177 573 179 575
rect 182 573 184 575
rect 196 573 198 575
rect 201 573 203 575
rect 206 573 208 575
rect 211 573 213 575
rect 216 573 218 575
rect 221 573 223 575
rect 226 573 228 575
rect 231 573 233 575
rect 236 573 238 575
rect 241 573 243 575
rect 246 573 248 575
rect 251 573 253 575
rect 256 573 258 575
rect 261 573 263 575
rect 266 573 268 575
rect 271 573 273 575
rect 276 573 278 575
rect 281 573 283 575
rect 286 573 288 575
rect 291 573 293 575
rect 296 573 298 575
rect 301 573 303 575
rect 306 573 308 575
rect 311 573 313 575
rect 316 573 318 575
rect 333 573 335 575
rect 338 573 340 575
rect 351 574 353 576
rect 356 574 358 576
rect 33 570 35 572
rect 169 570 171 572
rect 189 570 191 572
rect 325 570 327 572
rect 20 568 22 570
rect 25 568 27 570
rect 42 568 44 570
rect 47 568 49 570
rect 52 568 54 570
rect 57 568 59 570
rect 62 568 64 570
rect 67 568 69 570
rect 72 568 74 570
rect 77 568 79 570
rect 82 568 84 570
rect 87 568 89 570
rect 92 568 94 570
rect 97 568 99 570
rect 102 568 104 570
rect 107 568 109 570
rect 112 568 114 570
rect 117 568 119 570
rect 122 568 124 570
rect 127 568 129 570
rect 132 568 134 570
rect 137 568 139 570
rect 142 568 144 570
rect 147 568 149 570
rect 152 568 154 570
rect 157 568 159 570
rect 162 568 164 570
rect 177 568 179 570
rect 182 568 184 570
rect 196 568 198 570
rect 201 568 203 570
rect 206 568 208 570
rect 211 568 213 570
rect 216 568 218 570
rect 221 568 223 570
rect 226 568 228 570
rect 231 568 233 570
rect 236 568 238 570
rect 241 568 243 570
rect 246 568 248 570
rect 251 568 253 570
rect 256 568 258 570
rect 261 568 263 570
rect 266 568 268 570
rect 271 568 273 570
rect 276 568 278 570
rect 281 568 283 570
rect 286 568 288 570
rect 291 568 293 570
rect 296 568 298 570
rect 301 568 303 570
rect 306 568 308 570
rect 311 568 313 570
rect 316 568 318 570
rect 333 568 335 570
rect 338 568 340 570
rect 2 566 4 568
rect 7 566 9 568
rect 351 566 353 568
rect 356 566 358 568
rect 20 563 22 565
rect 25 563 27 565
rect 33 564 35 566
rect 42 563 44 565
rect 47 563 49 565
rect 52 563 54 565
rect 57 563 59 565
rect 62 563 64 565
rect 67 563 69 565
rect 72 563 74 565
rect 77 563 79 565
rect 82 563 84 565
rect 87 563 89 565
rect 92 563 94 565
rect 97 563 99 565
rect 102 563 104 565
rect 107 563 109 565
rect 112 563 114 565
rect 117 563 119 565
rect 122 563 124 565
rect 127 563 129 565
rect 132 563 134 565
rect 137 563 139 565
rect 142 563 144 565
rect 147 563 149 565
rect 152 563 154 565
rect 157 563 159 565
rect 162 563 164 565
rect 169 564 171 566
rect 177 563 179 565
rect 182 563 184 565
rect 189 564 191 566
rect 196 563 198 565
rect 201 563 203 565
rect 206 563 208 565
rect 211 563 213 565
rect 216 563 218 565
rect 221 563 223 565
rect 226 563 228 565
rect 231 563 233 565
rect 236 563 238 565
rect 241 563 243 565
rect 246 563 248 565
rect 251 563 253 565
rect 256 563 258 565
rect 261 563 263 565
rect 266 563 268 565
rect 271 563 273 565
rect 276 563 278 565
rect 281 563 283 565
rect 286 563 288 565
rect 291 563 293 565
rect 296 563 298 565
rect 301 563 303 565
rect 306 563 308 565
rect 311 563 313 565
rect 316 563 318 565
rect 325 564 327 566
rect 333 563 335 565
rect 338 563 340 565
rect 2 558 4 560
rect 7 558 9 560
rect 20 558 22 560
rect 25 558 27 560
rect 33 559 35 561
rect 42 558 44 560
rect 47 558 49 560
rect 52 558 54 560
rect 57 558 59 560
rect 62 558 64 560
rect 67 558 69 560
rect 72 558 74 560
rect 77 558 79 560
rect 82 558 84 560
rect 87 558 89 560
rect 92 558 94 560
rect 97 558 99 560
rect 102 558 104 560
rect 107 558 109 560
rect 112 558 114 560
rect 117 558 119 560
rect 122 558 124 560
rect 127 558 129 560
rect 132 558 134 560
rect 137 558 139 560
rect 142 558 144 560
rect 147 558 149 560
rect 152 558 154 560
rect 157 558 159 560
rect 162 558 164 560
rect 169 559 171 561
rect 177 558 179 560
rect 182 558 184 560
rect 189 559 191 561
rect 196 558 198 560
rect 201 558 203 560
rect 206 558 208 560
rect 211 558 213 560
rect 216 558 218 560
rect 221 558 223 560
rect 226 558 228 560
rect 231 558 233 560
rect 236 558 238 560
rect 241 558 243 560
rect 246 558 248 560
rect 251 558 253 560
rect 256 558 258 560
rect 261 558 263 560
rect 266 558 268 560
rect 271 558 273 560
rect 276 558 278 560
rect 281 558 283 560
rect 286 558 288 560
rect 291 558 293 560
rect 296 558 298 560
rect 301 558 303 560
rect 306 558 308 560
rect 311 558 313 560
rect 316 558 318 560
rect 325 559 327 561
rect 333 558 335 560
rect 338 558 340 560
rect 351 558 353 560
rect 356 558 358 560
rect 20 553 22 555
rect 25 553 27 555
rect 33 554 35 556
rect 42 553 44 555
rect 47 553 49 555
rect 52 553 54 555
rect 57 553 59 555
rect 62 553 64 555
rect 67 553 69 555
rect 72 553 74 555
rect 77 553 79 555
rect 82 553 84 555
rect 87 553 89 555
rect 92 553 94 555
rect 97 553 99 555
rect 102 553 104 555
rect 107 553 109 555
rect 112 553 114 555
rect 117 553 119 555
rect 122 553 124 555
rect 127 553 129 555
rect 132 553 134 555
rect 137 553 139 555
rect 142 553 144 555
rect 147 553 149 555
rect 152 553 154 555
rect 157 553 159 555
rect 162 553 164 555
rect 169 554 171 556
rect 177 553 179 555
rect 182 553 184 555
rect 189 554 191 556
rect 196 553 198 555
rect 201 553 203 555
rect 206 553 208 555
rect 211 553 213 555
rect 216 553 218 555
rect 221 553 223 555
rect 226 553 228 555
rect 231 553 233 555
rect 236 553 238 555
rect 241 553 243 555
rect 246 553 248 555
rect 251 553 253 555
rect 256 553 258 555
rect 261 553 263 555
rect 266 553 268 555
rect 271 553 273 555
rect 276 553 278 555
rect 281 553 283 555
rect 286 553 288 555
rect 291 553 293 555
rect 296 553 298 555
rect 301 553 303 555
rect 306 553 308 555
rect 311 553 313 555
rect 316 553 318 555
rect 325 554 327 556
rect 333 553 335 555
rect 338 553 340 555
rect 2 549 4 551
rect 7 549 9 551
rect 20 548 22 550
rect 25 548 27 550
rect 33 549 35 551
rect 42 548 44 550
rect 47 548 49 550
rect 52 548 54 550
rect 57 548 59 550
rect 62 548 64 550
rect 67 548 69 550
rect 72 548 74 550
rect 77 548 79 550
rect 82 548 84 550
rect 87 548 89 550
rect 92 548 94 550
rect 97 548 99 550
rect 102 548 104 550
rect 107 548 109 550
rect 112 548 114 550
rect 117 548 119 550
rect 122 548 124 550
rect 127 548 129 550
rect 132 548 134 550
rect 137 548 139 550
rect 142 548 144 550
rect 147 548 149 550
rect 152 548 154 550
rect 157 548 159 550
rect 162 548 164 550
rect 169 549 171 551
rect 177 548 179 550
rect 182 548 184 550
rect 189 549 191 551
rect 196 548 198 550
rect 201 548 203 550
rect 206 548 208 550
rect 211 548 213 550
rect 216 548 218 550
rect 221 548 223 550
rect 226 548 228 550
rect 231 548 233 550
rect 236 548 238 550
rect 241 548 243 550
rect 246 548 248 550
rect 251 548 253 550
rect 256 548 258 550
rect 261 548 263 550
rect 266 548 268 550
rect 271 548 273 550
rect 276 548 278 550
rect 281 548 283 550
rect 286 548 288 550
rect 291 548 293 550
rect 296 548 298 550
rect 301 548 303 550
rect 306 548 308 550
rect 311 548 313 550
rect 316 548 318 550
rect 325 549 327 551
rect 333 548 335 550
rect 338 548 340 550
rect 351 549 353 551
rect 356 549 358 551
rect 20 543 22 545
rect 25 543 27 545
rect 33 544 35 546
rect 169 544 171 546
rect 177 543 179 545
rect 182 543 184 545
rect 189 544 191 546
rect 325 544 327 546
rect 333 543 335 545
rect 338 543 340 545
rect 2 541 4 543
rect 7 541 9 543
rect 351 541 353 543
rect 356 541 358 543
rect 33 539 35 541
rect 41 538 43 540
rect 51 538 53 540
rect 61 538 63 540
rect 71 538 73 540
rect 81 538 83 540
rect 91 538 93 540
rect 101 538 103 540
rect 111 538 113 540
rect 150 538 152 540
rect 160 538 162 540
rect 169 539 171 541
rect 189 539 191 541
rect 198 538 200 540
rect 208 538 210 540
rect 247 538 249 540
rect 257 538 259 540
rect 267 538 269 540
rect 277 538 279 540
rect 287 538 289 540
rect 297 538 299 540
rect 307 538 309 540
rect 317 538 319 540
rect 325 539 327 541
rect 2 533 4 535
rect 7 533 9 535
rect 33 534 35 536
rect 41 533 43 535
rect 51 533 53 535
rect 61 533 63 535
rect 71 533 73 535
rect 81 533 83 535
rect 91 533 93 535
rect 101 533 103 535
rect 111 533 113 535
rect 150 533 152 535
rect 160 533 162 535
rect 169 534 171 536
rect 189 534 191 536
rect 198 533 200 535
rect 208 533 210 535
rect 247 533 249 535
rect 257 533 259 535
rect 267 533 269 535
rect 277 533 279 535
rect 287 533 289 535
rect 297 533 299 535
rect 307 533 309 535
rect 317 533 319 535
rect 325 534 327 536
rect 351 533 353 535
rect 356 533 358 535
rect 33 529 35 531
rect 41 528 43 530
rect 51 528 53 530
rect 61 528 63 530
rect 71 528 73 530
rect 81 528 83 530
rect 91 528 93 530
rect 101 528 103 530
rect 111 528 113 530
rect 150 528 152 530
rect 160 528 162 530
rect 169 529 171 531
rect 189 529 191 531
rect 198 528 200 530
rect 208 528 210 530
rect 247 528 249 530
rect 257 528 259 530
rect 267 528 269 530
rect 277 528 279 530
rect 287 528 289 530
rect 297 528 299 530
rect 307 528 309 530
rect 317 528 319 530
rect 325 529 327 531
rect 2 525 4 527
rect 7 525 9 527
rect 20 523 22 525
rect 25 523 27 525
rect 33 524 35 526
rect 169 524 171 526
rect 177 523 179 525
rect 182 523 184 525
rect 189 524 191 526
rect 325 524 327 526
rect 351 525 353 527
rect 356 525 358 527
rect 333 523 335 525
rect 338 523 340 525
rect 2 517 4 519
rect 7 517 9 519
rect 20 518 22 520
rect 25 518 27 520
rect 33 519 35 521
rect 42 518 44 520
rect 47 518 49 520
rect 52 518 54 520
rect 57 518 59 520
rect 62 518 64 520
rect 67 518 69 520
rect 72 518 74 520
rect 77 518 79 520
rect 82 518 84 520
rect 87 518 89 520
rect 92 518 94 520
rect 97 518 99 520
rect 102 518 104 520
rect 107 518 109 520
rect 112 518 114 520
rect 117 518 119 520
rect 122 518 124 520
rect 127 518 129 520
rect 132 518 134 520
rect 137 518 139 520
rect 142 518 144 520
rect 147 518 149 520
rect 152 518 154 520
rect 157 518 159 520
rect 162 518 164 520
rect 169 519 171 521
rect 177 518 179 520
rect 182 518 184 520
rect 189 519 191 521
rect 196 518 198 520
rect 201 518 203 520
rect 206 518 208 520
rect 211 518 213 520
rect 216 518 218 520
rect 221 518 223 520
rect 226 518 228 520
rect 231 518 233 520
rect 236 518 238 520
rect 241 518 243 520
rect 246 518 248 520
rect 251 518 253 520
rect 256 518 258 520
rect 261 518 263 520
rect 266 518 268 520
rect 271 518 273 520
rect 276 518 278 520
rect 281 518 283 520
rect 286 518 288 520
rect 291 518 293 520
rect 296 518 298 520
rect 301 518 303 520
rect 306 518 308 520
rect 311 518 313 520
rect 316 518 318 520
rect 325 519 327 521
rect 333 518 335 520
rect 338 518 340 520
rect 351 517 353 519
rect 356 517 358 519
rect 20 513 22 515
rect 25 513 27 515
rect 33 514 35 516
rect 42 513 44 515
rect 47 513 49 515
rect 52 513 54 515
rect 57 513 59 515
rect 62 513 64 515
rect 67 513 69 515
rect 72 513 74 515
rect 77 513 79 515
rect 82 513 84 515
rect 87 513 89 515
rect 92 513 94 515
rect 97 513 99 515
rect 102 513 104 515
rect 107 513 109 515
rect 112 513 114 515
rect 117 513 119 515
rect 122 513 124 515
rect 127 513 129 515
rect 132 513 134 515
rect 137 513 139 515
rect 142 513 144 515
rect 147 513 149 515
rect 152 513 154 515
rect 157 513 159 515
rect 162 513 164 515
rect 169 514 171 516
rect 177 513 179 515
rect 182 513 184 515
rect 189 514 191 516
rect 196 513 198 515
rect 201 513 203 515
rect 206 513 208 515
rect 211 513 213 515
rect 216 513 218 515
rect 221 513 223 515
rect 226 513 228 515
rect 231 513 233 515
rect 236 513 238 515
rect 241 513 243 515
rect 246 513 248 515
rect 251 513 253 515
rect 256 513 258 515
rect 261 513 263 515
rect 266 513 268 515
rect 271 513 273 515
rect 276 513 278 515
rect 281 513 283 515
rect 286 513 288 515
rect 291 513 293 515
rect 296 513 298 515
rect 301 513 303 515
rect 306 513 308 515
rect 311 513 313 515
rect 316 513 318 515
rect 325 514 327 516
rect 333 513 335 515
rect 338 513 340 515
rect 2 509 4 511
rect 7 509 9 511
rect 20 508 22 510
rect 25 508 27 510
rect 33 509 35 511
rect 42 508 44 510
rect 47 508 49 510
rect 52 508 54 510
rect 57 508 59 510
rect 62 508 64 510
rect 67 508 69 510
rect 72 508 74 510
rect 77 508 79 510
rect 82 508 84 510
rect 87 508 89 510
rect 92 508 94 510
rect 97 508 99 510
rect 102 508 104 510
rect 107 508 109 510
rect 112 508 114 510
rect 117 508 119 510
rect 122 508 124 510
rect 127 508 129 510
rect 132 508 134 510
rect 137 508 139 510
rect 142 508 144 510
rect 147 508 149 510
rect 152 508 154 510
rect 157 508 159 510
rect 162 508 164 510
rect 169 509 171 511
rect 177 508 179 510
rect 182 508 184 510
rect 189 509 191 511
rect 196 508 198 510
rect 201 508 203 510
rect 206 508 208 510
rect 211 508 213 510
rect 216 508 218 510
rect 221 508 223 510
rect 226 508 228 510
rect 231 508 233 510
rect 236 508 238 510
rect 241 508 243 510
rect 246 508 248 510
rect 251 508 253 510
rect 256 508 258 510
rect 261 508 263 510
rect 266 508 268 510
rect 271 508 273 510
rect 276 508 278 510
rect 281 508 283 510
rect 286 508 288 510
rect 291 508 293 510
rect 296 508 298 510
rect 301 508 303 510
rect 306 508 308 510
rect 311 508 313 510
rect 316 508 318 510
rect 325 509 327 511
rect 333 508 335 510
rect 338 508 340 510
rect 351 509 353 511
rect 356 509 358 511
rect 20 503 22 505
rect 25 503 27 505
rect 33 504 35 506
rect 42 503 44 505
rect 47 503 49 505
rect 52 503 54 505
rect 57 503 59 505
rect 62 503 64 505
rect 67 503 69 505
rect 72 503 74 505
rect 77 503 79 505
rect 82 503 84 505
rect 87 503 89 505
rect 92 503 94 505
rect 97 503 99 505
rect 102 503 104 505
rect 107 503 109 505
rect 112 503 114 505
rect 117 503 119 505
rect 122 503 124 505
rect 127 503 129 505
rect 132 503 134 505
rect 137 503 139 505
rect 142 503 144 505
rect 147 503 149 505
rect 152 503 154 505
rect 157 503 159 505
rect 162 503 164 505
rect 169 504 171 506
rect 177 503 179 505
rect 182 503 184 505
rect 189 504 191 506
rect 196 503 198 505
rect 201 503 203 505
rect 206 503 208 505
rect 211 503 213 505
rect 216 503 218 505
rect 221 503 223 505
rect 226 503 228 505
rect 231 503 233 505
rect 236 503 238 505
rect 241 503 243 505
rect 246 503 248 505
rect 251 503 253 505
rect 256 503 258 505
rect 261 503 263 505
rect 266 503 268 505
rect 271 503 273 505
rect 276 503 278 505
rect 281 503 283 505
rect 286 503 288 505
rect 291 503 293 505
rect 296 503 298 505
rect 301 503 303 505
rect 306 503 308 505
rect 311 503 313 505
rect 316 503 318 505
rect 325 504 327 506
rect 333 503 335 505
rect 338 503 340 505
rect 2 501 4 503
rect 7 501 9 503
rect 351 501 353 503
rect 356 501 358 503
rect 20 498 22 500
rect 25 498 27 500
rect 33 499 35 501
rect 42 498 44 500
rect 47 498 49 500
rect 52 498 54 500
rect 57 498 59 500
rect 62 498 64 500
rect 67 498 69 500
rect 72 498 74 500
rect 77 498 79 500
rect 82 498 84 500
rect 87 498 89 500
rect 92 498 94 500
rect 97 498 99 500
rect 102 498 104 500
rect 107 498 109 500
rect 112 498 114 500
rect 117 498 119 500
rect 122 498 124 500
rect 127 498 129 500
rect 132 498 134 500
rect 137 498 139 500
rect 142 498 144 500
rect 147 498 149 500
rect 152 498 154 500
rect 157 498 159 500
rect 162 498 164 500
rect 169 499 171 501
rect 177 498 179 500
rect 182 498 184 500
rect 189 499 191 501
rect 196 498 198 500
rect 201 498 203 500
rect 206 498 208 500
rect 211 498 213 500
rect 216 498 218 500
rect 221 498 223 500
rect 226 498 228 500
rect 231 498 233 500
rect 236 498 238 500
rect 241 498 243 500
rect 246 498 248 500
rect 251 498 253 500
rect 256 498 258 500
rect 261 498 263 500
rect 266 498 268 500
rect 271 498 273 500
rect 276 498 278 500
rect 281 498 283 500
rect 286 498 288 500
rect 291 498 293 500
rect 296 498 298 500
rect 301 498 303 500
rect 306 498 308 500
rect 311 498 313 500
rect 316 498 318 500
rect 325 499 327 501
rect 333 498 335 500
rect 338 498 340 500
rect 2 493 4 495
rect 7 493 9 495
rect 20 493 22 495
rect 25 493 27 495
rect 33 494 35 496
rect 42 493 44 495
rect 47 493 49 495
rect 52 493 54 495
rect 57 493 59 495
rect 62 493 64 495
rect 67 493 69 495
rect 72 493 74 495
rect 77 493 79 495
rect 82 493 84 495
rect 87 493 89 495
rect 92 493 94 495
rect 97 493 99 495
rect 102 493 104 495
rect 107 493 109 495
rect 112 493 114 495
rect 117 493 119 495
rect 122 493 124 495
rect 127 493 129 495
rect 132 493 134 495
rect 137 493 139 495
rect 142 493 144 495
rect 147 493 149 495
rect 152 493 154 495
rect 157 493 159 495
rect 162 493 164 495
rect 169 494 171 496
rect 177 493 179 495
rect 182 493 184 495
rect 189 494 191 496
rect 196 493 198 495
rect 201 493 203 495
rect 206 493 208 495
rect 211 493 213 495
rect 216 493 218 495
rect 221 493 223 495
rect 226 493 228 495
rect 231 493 233 495
rect 236 493 238 495
rect 241 493 243 495
rect 246 493 248 495
rect 251 493 253 495
rect 256 493 258 495
rect 261 493 263 495
rect 266 493 268 495
rect 271 493 273 495
rect 276 493 278 495
rect 281 493 283 495
rect 286 493 288 495
rect 291 493 293 495
rect 296 493 298 495
rect 301 493 303 495
rect 306 493 308 495
rect 311 493 313 495
rect 316 493 318 495
rect 325 494 327 496
rect 333 493 335 495
rect 338 493 340 495
rect 351 493 353 495
rect 356 493 358 495
rect 20 488 22 490
rect 25 488 27 490
rect 33 489 35 491
rect 42 488 44 490
rect 47 488 49 490
rect 52 488 54 490
rect 57 488 59 490
rect 62 488 64 490
rect 67 488 69 490
rect 72 488 74 490
rect 77 488 79 490
rect 82 488 84 490
rect 87 488 89 490
rect 92 488 94 490
rect 97 488 99 490
rect 102 488 104 490
rect 107 488 109 490
rect 112 488 114 490
rect 117 488 119 490
rect 122 488 124 490
rect 127 488 129 490
rect 132 488 134 490
rect 137 488 139 490
rect 142 488 144 490
rect 147 488 149 490
rect 152 488 154 490
rect 157 488 159 490
rect 162 488 164 490
rect 169 489 171 491
rect 177 488 179 490
rect 182 488 184 490
rect 189 489 191 491
rect 196 488 198 490
rect 201 488 203 490
rect 206 488 208 490
rect 211 488 213 490
rect 216 488 218 490
rect 221 488 223 490
rect 226 488 228 490
rect 231 488 233 490
rect 236 488 238 490
rect 241 488 243 490
rect 246 488 248 490
rect 251 488 253 490
rect 256 488 258 490
rect 261 488 263 490
rect 266 488 268 490
rect 271 488 273 490
rect 276 488 278 490
rect 281 488 283 490
rect 286 488 288 490
rect 291 488 293 490
rect 296 488 298 490
rect 301 488 303 490
rect 306 488 308 490
rect 311 488 313 490
rect 316 488 318 490
rect 325 489 327 491
rect 333 488 335 490
rect 338 488 340 490
rect 2 485 4 487
rect 7 485 9 487
rect 20 483 22 485
rect 25 483 27 485
rect 33 484 35 486
rect 42 483 44 485
rect 47 483 49 485
rect 52 483 54 485
rect 57 483 59 485
rect 62 483 64 485
rect 67 483 69 485
rect 72 483 74 485
rect 77 483 79 485
rect 82 483 84 485
rect 87 483 89 485
rect 92 483 94 485
rect 97 483 99 485
rect 102 483 104 485
rect 107 483 109 485
rect 112 483 114 485
rect 117 483 119 485
rect 122 483 124 485
rect 127 483 129 485
rect 132 483 134 485
rect 137 483 139 485
rect 142 483 144 485
rect 147 483 149 485
rect 152 483 154 485
rect 157 483 159 485
rect 162 483 164 485
rect 169 484 171 486
rect 177 483 179 485
rect 182 483 184 485
rect 189 484 191 486
rect 196 483 198 485
rect 201 483 203 485
rect 206 483 208 485
rect 211 483 213 485
rect 216 483 218 485
rect 221 483 223 485
rect 226 483 228 485
rect 231 483 233 485
rect 236 483 238 485
rect 241 483 243 485
rect 246 483 248 485
rect 251 483 253 485
rect 256 483 258 485
rect 261 483 263 485
rect 266 483 268 485
rect 271 483 273 485
rect 276 483 278 485
rect 281 483 283 485
rect 286 483 288 485
rect 291 483 293 485
rect 296 483 298 485
rect 301 483 303 485
rect 306 483 308 485
rect 311 483 313 485
rect 316 483 318 485
rect 325 484 327 486
rect 351 485 353 487
rect 356 485 358 487
rect 333 483 335 485
rect 338 483 340 485
rect 2 477 4 479
rect 7 477 9 479
rect 20 478 22 480
rect 25 478 27 480
rect 33 479 35 481
rect 169 479 171 481
rect 177 478 179 480
rect 182 478 184 480
rect 189 479 191 481
rect 325 479 327 481
rect 333 478 335 480
rect 338 478 340 480
rect 351 477 353 479
rect 356 477 358 479
rect 41 473 43 475
rect 51 473 53 475
rect 61 473 63 475
rect 71 473 73 475
rect 81 473 83 475
rect 91 473 93 475
rect 101 473 103 475
rect 111 473 113 475
rect 150 473 152 475
rect 160 473 162 475
rect 198 473 200 475
rect 208 473 210 475
rect 247 473 249 475
rect 257 473 259 475
rect 267 473 269 475
rect 277 473 279 475
rect 287 473 289 475
rect 297 473 299 475
rect 307 473 309 475
rect 317 473 319 475
rect 2 469 4 471
rect 7 469 9 471
rect 41 468 43 470
rect 51 468 53 470
rect 61 468 63 470
rect 71 468 73 470
rect 81 468 83 470
rect 91 468 93 470
rect 101 468 103 470
rect 111 468 113 470
rect 150 468 152 470
rect 160 468 162 470
rect 198 468 200 470
rect 208 468 210 470
rect 247 468 249 470
rect 257 468 259 470
rect 267 468 269 470
rect 277 468 279 470
rect 287 468 289 470
rect 297 468 299 470
rect 307 468 309 470
rect 317 468 319 470
rect 351 469 353 471
rect 356 469 358 471
rect 41 463 43 465
rect 51 463 53 465
rect 61 463 63 465
rect 71 463 73 465
rect 81 463 83 465
rect 91 463 93 465
rect 101 463 103 465
rect 111 463 113 465
rect 150 463 152 465
rect 160 463 162 465
rect 198 463 200 465
rect 208 463 210 465
rect 247 463 249 465
rect 257 463 259 465
rect 267 463 269 465
rect 277 463 279 465
rect 287 463 289 465
rect 297 463 299 465
rect 307 463 309 465
rect 317 463 319 465
rect 2 461 4 463
rect 7 461 9 463
rect 351 461 353 463
rect 356 461 358 463
rect 2 453 4 455
rect 7 453 9 455
rect 351 453 353 455
rect 356 453 358 455
rect 9 445 11 447
rect 17 445 19 447
rect 25 445 27 447
rect 41 445 43 447
rect 49 445 51 447
rect 57 445 59 447
rect 65 445 67 447
rect 73 445 75 447
rect 81 445 83 447
rect 89 445 91 447
rect 97 445 99 447
rect 105 445 107 447
rect 113 445 115 447
rect 150 445 152 447
rect 158 445 160 447
rect 181 445 183 447
rect 198 445 200 447
rect 206 445 208 447
rect 245 445 247 447
rect 253 445 255 447
rect 261 445 263 447
rect 269 445 271 447
rect 277 445 279 447
rect 285 445 287 447
rect 293 445 295 447
rect 301 445 303 447
rect 309 445 311 447
rect 317 445 319 447
rect 333 445 335 447
rect 341 445 343 447
rect 349 445 351 447
rect 9 440 11 442
rect 17 440 19 442
rect 25 440 27 442
rect 41 440 43 442
rect 49 440 51 442
rect 57 440 59 442
rect 65 440 67 442
rect 73 440 75 442
rect 81 440 83 442
rect 89 440 91 442
rect 97 440 99 442
rect 105 440 107 442
rect 113 440 115 442
rect 150 440 152 442
rect 158 440 160 442
rect 181 440 183 442
rect 198 440 200 442
rect 206 440 208 442
rect 245 440 247 442
rect 253 440 255 442
rect 261 440 263 442
rect 269 440 271 442
rect 277 440 279 442
rect 285 440 287 442
rect 293 440 295 442
rect 301 440 303 442
rect 309 440 311 442
rect 317 440 319 442
rect 333 440 335 442
rect 341 440 343 442
rect 349 440 351 442
rect 9 428 11 430
rect 17 428 19 430
rect 25 428 27 430
rect 41 428 43 430
rect 49 428 51 430
rect 57 428 59 430
rect 65 428 67 430
rect 73 428 75 430
rect 81 428 83 430
rect 89 428 91 430
rect 97 428 99 430
rect 105 428 107 430
rect 113 428 115 430
rect 150 428 152 430
rect 158 428 160 430
rect 181 428 183 430
rect 198 428 200 430
rect 206 428 208 430
rect 245 428 247 430
rect 253 428 255 430
rect 261 428 263 430
rect 269 428 271 430
rect 277 428 279 430
rect 285 428 287 430
rect 293 428 295 430
rect 301 428 303 430
rect 309 428 311 430
rect 317 428 319 430
rect 333 428 335 430
rect 341 428 343 430
rect 349 428 351 430
rect 9 423 11 425
rect 17 423 19 425
rect 25 423 27 425
rect 41 423 43 425
rect 49 423 51 425
rect 57 423 59 425
rect 65 423 67 425
rect 73 423 75 425
rect 81 423 83 425
rect 89 423 91 425
rect 97 423 99 425
rect 105 423 107 425
rect 113 423 115 425
rect 150 423 152 425
rect 158 423 160 425
rect 181 423 183 425
rect 198 423 200 425
rect 206 423 208 425
rect 245 423 247 425
rect 253 423 255 425
rect 261 423 263 425
rect 269 423 271 425
rect 277 423 279 425
rect 285 423 287 425
rect 293 423 295 425
rect 301 423 303 425
rect 309 423 311 425
rect 317 423 319 425
rect 333 423 335 425
rect 341 423 343 425
rect 349 423 351 425
rect 9 400 11 402
rect 17 400 19 402
rect 25 400 27 402
rect 41 400 43 402
rect 49 400 51 402
rect 57 400 59 402
rect 65 400 67 402
rect 73 400 75 402
rect 81 400 83 402
rect 89 400 91 402
rect 97 400 99 402
rect 105 400 107 402
rect 113 400 115 402
rect 150 400 152 402
rect 158 400 160 402
rect 181 400 183 402
rect 198 400 200 402
rect 206 400 208 402
rect 245 400 247 402
rect 253 400 255 402
rect 261 400 263 402
rect 269 400 271 402
rect 277 400 279 402
rect 285 400 287 402
rect 293 400 295 402
rect 301 400 303 402
rect 309 400 311 402
rect 317 400 319 402
rect 333 400 335 402
rect 341 400 343 402
rect 349 400 351 402
rect 9 395 11 397
rect 17 395 19 397
rect 25 395 27 397
rect 41 395 43 397
rect 49 395 51 397
rect 57 395 59 397
rect 65 395 67 397
rect 73 395 75 397
rect 81 395 83 397
rect 89 395 91 397
rect 97 395 99 397
rect 105 395 107 397
rect 113 395 115 397
rect 150 395 152 397
rect 158 395 160 397
rect 181 395 183 397
rect 198 395 200 397
rect 206 395 208 397
rect 245 395 247 397
rect 253 395 255 397
rect 261 395 263 397
rect 269 395 271 397
rect 277 395 279 397
rect 285 395 287 397
rect 293 395 295 397
rect 301 395 303 397
rect 309 395 311 397
rect 317 395 319 397
rect 333 395 335 397
rect 341 395 343 397
rect 349 395 351 397
rect 9 383 11 385
rect 17 383 19 385
rect 25 383 27 385
rect 41 383 43 385
rect 49 383 51 385
rect 57 383 59 385
rect 65 383 67 385
rect 73 383 75 385
rect 81 383 83 385
rect 89 383 91 385
rect 97 383 99 385
rect 105 383 107 385
rect 113 383 115 385
rect 150 383 152 385
rect 158 383 160 385
rect 181 383 183 385
rect 198 383 200 385
rect 206 383 208 385
rect 245 383 247 385
rect 253 383 255 385
rect 261 383 263 385
rect 269 383 271 385
rect 277 383 279 385
rect 285 383 287 385
rect 293 383 295 385
rect 301 383 303 385
rect 309 383 311 385
rect 317 383 319 385
rect 333 383 335 385
rect 341 383 343 385
rect 349 383 351 385
rect 357 383 359 385
rect 9 378 11 380
rect 17 378 19 380
rect 25 378 27 380
rect 41 378 43 380
rect 49 378 51 380
rect 57 378 59 380
rect 65 378 67 380
rect 73 378 75 380
rect 81 378 83 380
rect 89 378 91 380
rect 97 378 99 380
rect 105 378 107 380
rect 113 378 115 380
rect 150 378 152 380
rect 158 378 160 380
rect 181 378 183 380
rect 198 378 200 380
rect 206 378 208 380
rect 245 378 247 380
rect 253 378 255 380
rect 261 378 263 380
rect 269 378 271 380
rect 277 378 279 380
rect 285 378 287 380
rect 293 378 295 380
rect 301 378 303 380
rect 309 378 311 380
rect 317 378 319 380
rect 333 378 335 380
rect 341 378 343 380
rect 349 378 351 380
rect 357 378 359 380
rect 2 370 4 372
rect 7 370 9 372
rect 351 370 353 372
rect 356 370 358 372
rect 2 362 4 364
rect 7 362 9 364
rect 351 362 353 364
rect 356 362 358 364
rect 51 360 53 362
rect 61 360 63 362
rect 71 360 73 362
rect 81 360 83 362
rect 91 360 93 362
rect 101 360 103 362
rect 111 360 113 362
rect 154 360 156 362
rect 204 360 206 362
rect 247 360 249 362
rect 257 360 259 362
rect 267 360 269 362
rect 277 360 279 362
rect 287 360 289 362
rect 297 360 299 362
rect 307 360 309 362
rect 2 354 4 356
rect 7 354 9 356
rect 51 355 53 357
rect 61 355 63 357
rect 71 355 73 357
rect 81 355 83 357
rect 91 355 93 357
rect 101 355 103 357
rect 111 355 113 357
rect 154 355 156 357
rect 204 355 206 357
rect 247 355 249 357
rect 257 355 259 357
rect 267 355 269 357
rect 277 355 279 357
rect 287 355 289 357
rect 297 355 299 357
rect 307 355 309 357
rect 351 354 353 356
rect 356 354 358 356
rect 51 350 53 352
rect 61 350 63 352
rect 71 350 73 352
rect 81 350 83 352
rect 91 350 93 352
rect 101 350 103 352
rect 111 350 113 352
rect 154 350 156 352
rect 204 350 206 352
rect 247 350 249 352
rect 257 350 259 352
rect 267 350 269 352
rect 277 350 279 352
rect 287 350 289 352
rect 297 350 299 352
rect 307 350 309 352
rect 2 346 4 348
rect 7 346 9 348
rect 20 345 22 347
rect 25 345 27 347
rect 177 345 179 347
rect 182 345 184 347
rect 333 345 335 347
rect 338 345 340 347
rect 351 346 353 348
rect 356 346 358 348
rect 40 342 42 344
rect 162 342 164 344
rect 196 342 198 344
rect 318 342 320 344
rect 20 340 22 342
rect 25 340 27 342
rect 47 340 49 342
rect 52 340 54 342
rect 57 340 59 342
rect 62 340 64 342
rect 67 340 69 342
rect 72 340 74 342
rect 77 340 79 342
rect 82 340 84 342
rect 87 340 89 342
rect 92 340 94 342
rect 97 340 99 342
rect 102 340 104 342
rect 107 340 109 342
rect 112 340 114 342
rect 117 340 119 342
rect 122 340 124 342
rect 127 340 129 342
rect 132 340 134 342
rect 137 340 139 342
rect 142 340 144 342
rect 147 340 149 342
rect 152 340 154 342
rect 177 340 179 342
rect 182 340 184 342
rect 206 340 208 342
rect 211 340 213 342
rect 216 340 218 342
rect 221 340 223 342
rect 226 340 228 342
rect 231 340 233 342
rect 236 340 238 342
rect 241 340 243 342
rect 246 340 248 342
rect 251 340 253 342
rect 256 340 258 342
rect 261 340 263 342
rect 266 340 268 342
rect 271 340 273 342
rect 276 340 278 342
rect 281 340 283 342
rect 286 340 288 342
rect 291 340 293 342
rect 296 340 298 342
rect 301 340 303 342
rect 306 340 308 342
rect 311 340 313 342
rect 333 340 335 342
rect 338 340 340 342
rect 2 338 4 340
rect 7 338 9 340
rect 40 337 42 339
rect 162 337 164 339
rect 196 337 198 339
rect 318 337 320 339
rect 351 338 353 340
rect 356 338 358 340
rect 20 335 22 337
rect 25 335 27 337
rect 47 335 49 337
rect 52 335 54 337
rect 57 335 59 337
rect 62 335 64 337
rect 67 335 69 337
rect 72 335 74 337
rect 77 335 79 337
rect 82 335 84 337
rect 87 335 89 337
rect 92 335 94 337
rect 97 335 99 337
rect 102 335 104 337
rect 107 335 109 337
rect 112 335 114 337
rect 117 335 119 337
rect 122 335 124 337
rect 127 335 129 337
rect 132 335 134 337
rect 137 335 139 337
rect 142 335 144 337
rect 147 335 149 337
rect 152 335 154 337
rect 177 335 179 337
rect 182 335 184 337
rect 206 335 208 337
rect 211 335 213 337
rect 216 335 218 337
rect 221 335 223 337
rect 226 335 228 337
rect 231 335 233 337
rect 236 335 238 337
rect 241 335 243 337
rect 246 335 248 337
rect 251 335 253 337
rect 256 335 258 337
rect 261 335 263 337
rect 266 335 268 337
rect 271 335 273 337
rect 276 335 278 337
rect 281 335 283 337
rect 286 335 288 337
rect 291 335 293 337
rect 296 335 298 337
rect 301 335 303 337
rect 306 335 308 337
rect 311 335 313 337
rect 333 335 335 337
rect 338 335 340 337
rect 40 332 42 334
rect 162 332 164 334
rect 196 332 198 334
rect 318 332 320 334
rect 2 330 4 332
rect 7 330 9 332
rect 20 330 22 332
rect 25 330 27 332
rect 47 330 49 332
rect 52 330 54 332
rect 57 330 59 332
rect 62 330 64 332
rect 67 330 69 332
rect 72 330 74 332
rect 77 330 79 332
rect 82 330 84 332
rect 87 330 89 332
rect 92 330 94 332
rect 97 330 99 332
rect 102 330 104 332
rect 107 330 109 332
rect 112 330 114 332
rect 117 330 119 332
rect 122 330 124 332
rect 127 330 129 332
rect 132 330 134 332
rect 137 330 139 332
rect 142 330 144 332
rect 147 330 149 332
rect 152 330 154 332
rect 177 330 179 332
rect 182 330 184 332
rect 206 330 208 332
rect 211 330 213 332
rect 216 330 218 332
rect 221 330 223 332
rect 226 330 228 332
rect 231 330 233 332
rect 236 330 238 332
rect 241 330 243 332
rect 246 330 248 332
rect 251 330 253 332
rect 256 330 258 332
rect 261 330 263 332
rect 266 330 268 332
rect 271 330 273 332
rect 276 330 278 332
rect 281 330 283 332
rect 286 330 288 332
rect 291 330 293 332
rect 296 330 298 332
rect 301 330 303 332
rect 306 330 308 332
rect 311 330 313 332
rect 333 330 335 332
rect 338 330 340 332
rect 351 330 353 332
rect 356 330 358 332
rect 40 327 42 329
rect 162 327 164 329
rect 196 327 198 329
rect 318 327 320 329
rect 20 325 22 327
rect 25 325 27 327
rect 47 325 49 327
rect 52 325 54 327
rect 57 325 59 327
rect 62 325 64 327
rect 67 325 69 327
rect 72 325 74 327
rect 77 325 79 327
rect 82 325 84 327
rect 87 325 89 327
rect 92 325 94 327
rect 97 325 99 327
rect 102 325 104 327
rect 107 325 109 327
rect 112 325 114 327
rect 117 325 119 327
rect 122 325 124 327
rect 127 325 129 327
rect 132 325 134 327
rect 137 325 139 327
rect 142 325 144 327
rect 147 325 149 327
rect 152 325 154 327
rect 177 325 179 327
rect 182 325 184 327
rect 206 325 208 327
rect 211 325 213 327
rect 216 325 218 327
rect 221 325 223 327
rect 226 325 228 327
rect 231 325 233 327
rect 236 325 238 327
rect 241 325 243 327
rect 246 325 248 327
rect 251 325 253 327
rect 256 325 258 327
rect 261 325 263 327
rect 266 325 268 327
rect 271 325 273 327
rect 276 325 278 327
rect 281 325 283 327
rect 286 325 288 327
rect 291 325 293 327
rect 296 325 298 327
rect 301 325 303 327
rect 306 325 308 327
rect 311 325 313 327
rect 333 325 335 327
rect 338 325 340 327
rect 2 322 4 324
rect 7 322 9 324
rect 40 322 42 324
rect 162 322 164 324
rect 196 322 198 324
rect 318 322 320 324
rect 351 322 353 324
rect 356 322 358 324
rect 20 320 22 322
rect 25 320 27 322
rect 47 320 49 322
rect 52 320 54 322
rect 57 320 59 322
rect 62 320 64 322
rect 67 320 69 322
rect 72 320 74 322
rect 77 320 79 322
rect 82 320 84 322
rect 87 320 89 322
rect 92 320 94 322
rect 97 320 99 322
rect 102 320 104 322
rect 107 320 109 322
rect 112 320 114 322
rect 117 320 119 322
rect 122 320 124 322
rect 127 320 129 322
rect 132 320 134 322
rect 137 320 139 322
rect 142 320 144 322
rect 147 320 149 322
rect 152 320 154 322
rect 177 320 179 322
rect 182 320 184 322
rect 206 320 208 322
rect 211 320 213 322
rect 216 320 218 322
rect 221 320 223 322
rect 226 320 228 322
rect 231 320 233 322
rect 236 320 238 322
rect 241 320 243 322
rect 246 320 248 322
rect 251 320 253 322
rect 256 320 258 322
rect 261 320 263 322
rect 266 320 268 322
rect 271 320 273 322
rect 276 320 278 322
rect 281 320 283 322
rect 286 320 288 322
rect 291 320 293 322
rect 296 320 298 322
rect 301 320 303 322
rect 306 320 308 322
rect 311 320 313 322
rect 333 320 335 322
rect 338 320 340 322
rect 40 317 42 319
rect 162 317 164 319
rect 196 317 198 319
rect 318 317 320 319
rect 2 314 4 316
rect 7 314 9 316
rect 20 315 22 317
rect 25 315 27 317
rect 47 315 49 317
rect 52 315 54 317
rect 57 315 59 317
rect 62 315 64 317
rect 67 315 69 317
rect 72 315 74 317
rect 77 315 79 317
rect 82 315 84 317
rect 87 315 89 317
rect 92 315 94 317
rect 97 315 99 317
rect 102 315 104 317
rect 107 315 109 317
rect 112 315 114 317
rect 117 315 119 317
rect 122 315 124 317
rect 127 315 129 317
rect 132 315 134 317
rect 137 315 139 317
rect 142 315 144 317
rect 147 315 149 317
rect 152 315 154 317
rect 177 315 179 317
rect 182 315 184 317
rect 206 315 208 317
rect 211 315 213 317
rect 216 315 218 317
rect 221 315 223 317
rect 226 315 228 317
rect 231 315 233 317
rect 236 315 238 317
rect 241 315 243 317
rect 246 315 248 317
rect 251 315 253 317
rect 256 315 258 317
rect 261 315 263 317
rect 266 315 268 317
rect 271 315 273 317
rect 276 315 278 317
rect 281 315 283 317
rect 286 315 288 317
rect 291 315 293 317
rect 296 315 298 317
rect 301 315 303 317
rect 306 315 308 317
rect 311 315 313 317
rect 333 315 335 317
rect 338 315 340 317
rect 351 314 353 316
rect 356 314 358 316
rect 40 312 42 314
rect 162 312 164 314
rect 196 312 198 314
rect 318 312 320 314
rect 20 310 22 312
rect 25 310 27 312
rect 47 310 49 312
rect 52 310 54 312
rect 57 310 59 312
rect 62 310 64 312
rect 67 310 69 312
rect 72 310 74 312
rect 77 310 79 312
rect 82 310 84 312
rect 87 310 89 312
rect 92 310 94 312
rect 97 310 99 312
rect 102 310 104 312
rect 107 310 109 312
rect 112 310 114 312
rect 117 310 119 312
rect 122 310 124 312
rect 127 310 129 312
rect 132 310 134 312
rect 137 310 139 312
rect 142 310 144 312
rect 147 310 149 312
rect 152 310 154 312
rect 177 310 179 312
rect 182 310 184 312
rect 206 310 208 312
rect 211 310 213 312
rect 216 310 218 312
rect 221 310 223 312
rect 226 310 228 312
rect 231 310 233 312
rect 236 310 238 312
rect 241 310 243 312
rect 246 310 248 312
rect 251 310 253 312
rect 256 310 258 312
rect 261 310 263 312
rect 266 310 268 312
rect 271 310 273 312
rect 276 310 278 312
rect 281 310 283 312
rect 286 310 288 312
rect 291 310 293 312
rect 296 310 298 312
rect 301 310 303 312
rect 306 310 308 312
rect 311 310 313 312
rect 333 310 335 312
rect 338 310 340 312
rect 2 306 4 308
rect 7 306 9 308
rect 40 307 42 309
rect 162 307 164 309
rect 196 307 198 309
rect 318 307 320 309
rect 20 305 22 307
rect 25 305 27 307
rect 47 305 49 307
rect 52 305 54 307
rect 57 305 59 307
rect 62 305 64 307
rect 67 305 69 307
rect 72 305 74 307
rect 77 305 79 307
rect 82 305 84 307
rect 87 305 89 307
rect 92 305 94 307
rect 97 305 99 307
rect 102 305 104 307
rect 107 305 109 307
rect 112 305 114 307
rect 117 305 119 307
rect 122 305 124 307
rect 127 305 129 307
rect 132 305 134 307
rect 137 305 139 307
rect 142 305 144 307
rect 147 305 149 307
rect 152 305 154 307
rect 177 305 179 307
rect 182 305 184 307
rect 206 305 208 307
rect 211 305 213 307
rect 216 305 218 307
rect 221 305 223 307
rect 226 305 228 307
rect 231 305 233 307
rect 236 305 238 307
rect 241 305 243 307
rect 246 305 248 307
rect 251 305 253 307
rect 256 305 258 307
rect 261 305 263 307
rect 266 305 268 307
rect 271 305 273 307
rect 276 305 278 307
rect 281 305 283 307
rect 286 305 288 307
rect 291 305 293 307
rect 296 305 298 307
rect 301 305 303 307
rect 306 305 308 307
rect 311 305 313 307
rect 333 305 335 307
rect 338 305 340 307
rect 351 306 353 308
rect 356 306 358 308
rect 40 302 42 304
rect 162 302 164 304
rect 196 302 198 304
rect 318 302 320 304
rect 20 300 22 302
rect 25 300 27 302
rect 177 300 179 302
rect 182 300 184 302
rect 333 300 335 302
rect 338 300 340 302
rect 2 298 4 300
rect 7 298 9 300
rect 40 297 42 299
rect 162 297 164 299
rect 196 297 198 299
rect 318 297 320 299
rect 351 298 353 300
rect 356 298 358 300
rect 51 295 53 297
rect 61 295 63 297
rect 71 295 73 297
rect 81 295 83 297
rect 91 295 93 297
rect 101 295 103 297
rect 111 295 113 297
rect 154 295 156 297
rect 204 295 206 297
rect 247 295 249 297
rect 257 295 259 297
rect 267 295 269 297
rect 277 295 279 297
rect 287 295 289 297
rect 297 295 299 297
rect 307 295 309 297
rect 40 292 42 294
rect 162 292 164 294
rect 196 292 198 294
rect 318 292 320 294
rect 2 290 4 292
rect 7 290 9 292
rect 51 290 53 292
rect 61 290 63 292
rect 71 290 73 292
rect 81 290 83 292
rect 91 290 93 292
rect 101 290 103 292
rect 111 290 113 292
rect 154 290 156 292
rect 204 290 206 292
rect 247 290 249 292
rect 257 290 259 292
rect 267 290 269 292
rect 277 290 279 292
rect 287 290 289 292
rect 297 290 299 292
rect 307 290 309 292
rect 351 290 353 292
rect 356 290 358 292
rect 40 287 42 289
rect 162 287 164 289
rect 196 287 198 289
rect 318 287 320 289
rect 51 285 53 287
rect 61 285 63 287
rect 71 285 73 287
rect 81 285 83 287
rect 91 285 93 287
rect 101 285 103 287
rect 111 285 113 287
rect 154 285 156 287
rect 204 285 206 287
rect 247 285 249 287
rect 257 285 259 287
rect 267 285 269 287
rect 277 285 279 287
rect 287 285 289 287
rect 297 285 299 287
rect 307 285 309 287
rect 2 282 4 284
rect 7 282 9 284
rect 40 282 42 284
rect 162 282 164 284
rect 196 282 198 284
rect 318 282 320 284
rect 351 282 353 284
rect 356 282 358 284
rect 20 280 22 282
rect 25 280 27 282
rect 177 280 179 282
rect 182 280 184 282
rect 333 280 335 282
rect 338 280 340 282
rect 40 277 42 279
rect 162 277 164 279
rect 196 277 198 279
rect 318 277 320 279
rect 2 274 4 276
rect 7 274 9 276
rect 20 275 22 277
rect 25 275 27 277
rect 47 275 49 277
rect 52 275 54 277
rect 57 275 59 277
rect 62 275 64 277
rect 67 275 69 277
rect 72 275 74 277
rect 77 275 79 277
rect 82 275 84 277
rect 87 275 89 277
rect 92 275 94 277
rect 97 275 99 277
rect 102 275 104 277
rect 107 275 109 277
rect 112 275 114 277
rect 117 275 119 277
rect 122 275 124 277
rect 127 275 129 277
rect 132 275 134 277
rect 137 275 139 277
rect 142 275 144 277
rect 147 275 149 277
rect 152 275 154 277
rect 177 275 179 277
rect 182 275 184 277
rect 206 275 208 277
rect 211 275 213 277
rect 216 275 218 277
rect 221 275 223 277
rect 226 275 228 277
rect 231 275 233 277
rect 236 275 238 277
rect 241 275 243 277
rect 246 275 248 277
rect 251 275 253 277
rect 256 275 258 277
rect 261 275 263 277
rect 266 275 268 277
rect 271 275 273 277
rect 276 275 278 277
rect 281 275 283 277
rect 286 275 288 277
rect 291 275 293 277
rect 296 275 298 277
rect 301 275 303 277
rect 306 275 308 277
rect 311 275 313 277
rect 333 275 335 277
rect 338 275 340 277
rect 351 274 353 276
rect 356 274 358 276
rect 40 272 42 274
rect 162 272 164 274
rect 196 272 198 274
rect 318 272 320 274
rect 20 270 22 272
rect 25 270 27 272
rect 47 270 49 272
rect 52 270 54 272
rect 57 270 59 272
rect 62 270 64 272
rect 67 270 69 272
rect 72 270 74 272
rect 77 270 79 272
rect 82 270 84 272
rect 87 270 89 272
rect 92 270 94 272
rect 97 270 99 272
rect 102 270 104 272
rect 107 270 109 272
rect 112 270 114 272
rect 117 270 119 272
rect 122 270 124 272
rect 127 270 129 272
rect 132 270 134 272
rect 137 270 139 272
rect 142 270 144 272
rect 147 270 149 272
rect 152 270 154 272
rect 177 270 179 272
rect 182 270 184 272
rect 206 270 208 272
rect 211 270 213 272
rect 216 270 218 272
rect 221 270 223 272
rect 226 270 228 272
rect 231 270 233 272
rect 236 270 238 272
rect 241 270 243 272
rect 246 270 248 272
rect 251 270 253 272
rect 256 270 258 272
rect 261 270 263 272
rect 266 270 268 272
rect 271 270 273 272
rect 276 270 278 272
rect 281 270 283 272
rect 286 270 288 272
rect 291 270 293 272
rect 296 270 298 272
rect 301 270 303 272
rect 306 270 308 272
rect 311 270 313 272
rect 333 270 335 272
rect 338 270 340 272
rect 2 266 4 268
rect 7 266 9 268
rect 40 267 42 269
rect 162 267 164 269
rect 196 267 198 269
rect 318 267 320 269
rect 20 265 22 267
rect 25 265 27 267
rect 47 265 49 267
rect 52 265 54 267
rect 57 265 59 267
rect 62 265 64 267
rect 67 265 69 267
rect 72 265 74 267
rect 77 265 79 267
rect 82 265 84 267
rect 87 265 89 267
rect 92 265 94 267
rect 97 265 99 267
rect 102 265 104 267
rect 107 265 109 267
rect 112 265 114 267
rect 117 265 119 267
rect 122 265 124 267
rect 127 265 129 267
rect 132 265 134 267
rect 137 265 139 267
rect 142 265 144 267
rect 147 265 149 267
rect 152 265 154 267
rect 177 265 179 267
rect 182 265 184 267
rect 206 265 208 267
rect 211 265 213 267
rect 216 265 218 267
rect 221 265 223 267
rect 226 265 228 267
rect 231 265 233 267
rect 236 265 238 267
rect 241 265 243 267
rect 246 265 248 267
rect 251 265 253 267
rect 256 265 258 267
rect 261 265 263 267
rect 266 265 268 267
rect 271 265 273 267
rect 276 265 278 267
rect 281 265 283 267
rect 286 265 288 267
rect 291 265 293 267
rect 296 265 298 267
rect 301 265 303 267
rect 306 265 308 267
rect 311 265 313 267
rect 333 265 335 267
rect 338 265 340 267
rect 351 266 353 268
rect 356 266 358 268
rect 40 262 42 264
rect 162 262 164 264
rect 20 260 22 262
rect 25 260 27 262
rect 47 260 49 262
rect 52 260 54 262
rect 57 260 59 262
rect 62 260 64 262
rect 67 260 69 262
rect 72 260 74 262
rect 77 260 79 262
rect 82 260 84 262
rect 87 260 89 262
rect 92 260 94 262
rect 97 260 99 262
rect 102 260 104 262
rect 107 260 109 262
rect 112 260 114 262
rect 117 260 119 262
rect 122 260 124 262
rect 127 260 129 262
rect 132 260 134 262
rect 137 260 139 262
rect 142 260 144 262
rect 147 260 149 262
rect 152 260 154 262
rect 177 260 179 262
rect 182 260 184 262
rect 206 260 208 262
rect 211 260 213 262
rect 216 260 218 262
rect 221 260 223 262
rect 226 260 228 262
rect 231 260 233 262
rect 236 260 238 262
rect 241 260 243 262
rect 246 260 248 262
rect 251 260 253 262
rect 256 260 258 262
rect 261 260 263 262
rect 266 260 268 262
rect 271 260 273 262
rect 276 260 278 262
rect 281 260 283 262
rect 286 260 288 262
rect 291 260 293 262
rect 296 260 298 262
rect 301 260 303 262
rect 306 260 308 262
rect 311 260 313 262
rect 333 260 335 262
rect 338 260 340 262
rect 2 258 4 260
rect 7 258 9 260
rect 351 258 353 260
rect 356 258 358 260
rect 20 255 22 257
rect 25 255 27 257
rect 40 256 42 258
rect 47 255 49 257
rect 52 255 54 257
rect 57 255 59 257
rect 62 255 64 257
rect 67 255 69 257
rect 72 255 74 257
rect 77 255 79 257
rect 82 255 84 257
rect 87 255 89 257
rect 92 255 94 257
rect 97 255 99 257
rect 102 255 104 257
rect 107 255 109 257
rect 112 255 114 257
rect 117 255 119 257
rect 122 255 124 257
rect 127 255 129 257
rect 132 255 134 257
rect 137 255 139 257
rect 142 255 144 257
rect 147 255 149 257
rect 152 255 154 257
rect 162 256 164 258
rect 177 255 179 257
rect 182 255 184 257
rect 206 255 208 257
rect 211 255 213 257
rect 216 255 218 257
rect 221 255 223 257
rect 226 255 228 257
rect 231 255 233 257
rect 236 255 238 257
rect 241 255 243 257
rect 246 255 248 257
rect 251 255 253 257
rect 256 255 258 257
rect 261 255 263 257
rect 266 255 268 257
rect 271 255 273 257
rect 276 255 278 257
rect 281 255 283 257
rect 286 255 288 257
rect 291 255 293 257
rect 296 255 298 257
rect 301 255 303 257
rect 306 255 308 257
rect 311 255 313 257
rect 333 255 335 257
rect 338 255 340 257
rect 2 250 4 252
rect 7 250 9 252
rect 20 250 22 252
rect 25 250 27 252
rect 40 251 42 253
rect 47 250 49 252
rect 52 250 54 252
rect 57 250 59 252
rect 62 250 64 252
rect 67 250 69 252
rect 72 250 74 252
rect 77 250 79 252
rect 82 250 84 252
rect 87 250 89 252
rect 92 250 94 252
rect 97 250 99 252
rect 102 250 104 252
rect 107 250 109 252
rect 112 250 114 252
rect 117 250 119 252
rect 122 250 124 252
rect 127 250 129 252
rect 132 250 134 252
rect 137 250 139 252
rect 142 250 144 252
rect 147 250 149 252
rect 152 250 154 252
rect 162 251 164 253
rect 177 250 179 252
rect 182 250 184 252
rect 196 251 198 253
rect 206 250 208 252
rect 211 250 213 252
rect 216 250 218 252
rect 221 250 223 252
rect 226 250 228 252
rect 231 250 233 252
rect 236 250 238 252
rect 241 250 243 252
rect 246 250 248 252
rect 251 250 253 252
rect 256 250 258 252
rect 261 250 263 252
rect 266 250 268 252
rect 271 250 273 252
rect 276 250 278 252
rect 281 250 283 252
rect 286 250 288 252
rect 291 250 293 252
rect 296 250 298 252
rect 301 250 303 252
rect 306 250 308 252
rect 311 250 313 252
rect 318 251 320 253
rect 333 250 335 252
rect 338 250 340 252
rect 351 250 353 252
rect 356 250 358 252
rect 20 245 22 247
rect 25 245 27 247
rect 40 246 42 248
rect 47 245 49 247
rect 52 245 54 247
rect 57 245 59 247
rect 62 245 64 247
rect 67 245 69 247
rect 72 245 74 247
rect 77 245 79 247
rect 82 245 84 247
rect 87 245 89 247
rect 92 245 94 247
rect 97 245 99 247
rect 102 245 104 247
rect 107 245 109 247
rect 112 245 114 247
rect 117 245 119 247
rect 122 245 124 247
rect 127 245 129 247
rect 132 245 134 247
rect 137 245 139 247
rect 142 245 144 247
rect 147 245 149 247
rect 152 245 154 247
rect 162 246 164 248
rect 177 245 179 247
rect 182 245 184 247
rect 196 246 198 248
rect 206 245 208 247
rect 211 245 213 247
rect 216 245 218 247
rect 221 245 223 247
rect 226 245 228 247
rect 231 245 233 247
rect 236 245 238 247
rect 241 245 243 247
rect 246 245 248 247
rect 251 245 253 247
rect 256 245 258 247
rect 261 245 263 247
rect 266 245 268 247
rect 271 245 273 247
rect 276 245 278 247
rect 281 245 283 247
rect 286 245 288 247
rect 291 245 293 247
rect 296 245 298 247
rect 301 245 303 247
rect 306 245 308 247
rect 311 245 313 247
rect 318 246 320 248
rect 333 245 335 247
rect 338 245 340 247
rect 2 241 4 243
rect 7 241 9 243
rect 20 240 22 242
rect 25 240 27 242
rect 40 241 42 243
rect 47 240 49 242
rect 52 240 54 242
rect 57 240 59 242
rect 62 240 64 242
rect 67 240 69 242
rect 72 240 74 242
rect 77 240 79 242
rect 82 240 84 242
rect 87 240 89 242
rect 92 240 94 242
rect 97 240 99 242
rect 102 240 104 242
rect 107 240 109 242
rect 112 240 114 242
rect 117 240 119 242
rect 122 240 124 242
rect 127 240 129 242
rect 132 240 134 242
rect 137 240 139 242
rect 142 240 144 242
rect 147 240 149 242
rect 152 240 154 242
rect 162 241 164 243
rect 177 240 179 242
rect 182 240 184 242
rect 196 241 198 243
rect 206 240 208 242
rect 211 240 213 242
rect 216 240 218 242
rect 221 240 223 242
rect 226 240 228 242
rect 231 240 233 242
rect 236 240 238 242
rect 241 240 243 242
rect 246 240 248 242
rect 251 240 253 242
rect 256 240 258 242
rect 261 240 263 242
rect 266 240 268 242
rect 271 240 273 242
rect 276 240 278 242
rect 281 240 283 242
rect 286 240 288 242
rect 291 240 293 242
rect 296 240 298 242
rect 301 240 303 242
rect 306 240 308 242
rect 311 240 313 242
rect 318 241 320 243
rect 333 240 335 242
rect 338 240 340 242
rect 351 241 353 243
rect 356 241 358 243
rect 20 235 22 237
rect 25 235 27 237
rect 40 236 42 238
rect 162 236 164 238
rect 177 235 179 237
rect 182 235 184 237
rect 196 236 198 238
rect 318 236 320 238
rect 333 235 335 237
rect 338 235 340 237
rect 2 233 4 235
rect 7 233 9 235
rect 351 233 353 235
rect 356 233 358 235
rect 40 231 42 233
rect 51 230 53 232
rect 61 230 63 232
rect 71 230 73 232
rect 81 230 83 232
rect 91 230 93 232
rect 101 230 103 232
rect 111 230 113 232
rect 154 230 156 232
rect 162 231 164 233
rect 196 231 198 233
rect 204 230 206 232
rect 247 230 249 232
rect 257 230 259 232
rect 267 230 269 232
rect 277 230 279 232
rect 287 230 289 232
rect 297 230 299 232
rect 307 230 309 232
rect 318 231 320 233
rect 2 225 4 227
rect 7 225 9 227
rect 51 225 53 227
rect 61 225 63 227
rect 71 225 73 227
rect 81 225 83 227
rect 91 225 93 227
rect 101 225 103 227
rect 111 225 113 227
rect 154 225 156 227
rect 196 226 198 228
rect 204 225 206 227
rect 247 225 249 227
rect 257 225 259 227
rect 267 225 269 227
rect 277 225 279 227
rect 287 225 289 227
rect 297 225 299 227
rect 307 225 309 227
rect 318 226 320 228
rect 351 225 353 227
rect 356 225 358 227
rect 51 220 53 222
rect 61 220 63 222
rect 71 220 73 222
rect 81 220 83 222
rect 91 220 93 222
rect 101 220 103 222
rect 111 220 113 222
rect 154 220 156 222
rect 196 221 198 223
rect 204 220 206 222
rect 247 220 249 222
rect 257 220 259 222
rect 267 220 269 222
rect 277 220 279 222
rect 287 220 289 222
rect 297 220 299 222
rect 307 220 309 222
rect 318 221 320 223
rect 2 217 4 219
rect 7 217 9 219
rect 20 215 22 217
rect 25 215 27 217
rect 40 216 42 218
rect 162 216 164 218
rect 177 215 179 217
rect 182 215 184 217
rect 196 216 198 218
rect 318 216 320 218
rect 351 217 353 219
rect 356 217 358 219
rect 333 215 335 217
rect 338 215 340 217
rect 2 209 4 211
rect 7 209 9 211
rect 20 210 22 212
rect 25 210 27 212
rect 40 211 42 213
rect 47 210 49 212
rect 52 210 54 212
rect 57 210 59 212
rect 62 210 64 212
rect 67 210 69 212
rect 72 210 74 212
rect 77 210 79 212
rect 82 210 84 212
rect 87 210 89 212
rect 92 210 94 212
rect 97 210 99 212
rect 102 210 104 212
rect 107 210 109 212
rect 112 210 114 212
rect 117 210 119 212
rect 122 210 124 212
rect 127 210 129 212
rect 132 210 134 212
rect 137 210 139 212
rect 142 210 144 212
rect 147 210 149 212
rect 152 210 154 212
rect 162 211 164 213
rect 177 210 179 212
rect 182 210 184 212
rect 196 211 198 213
rect 206 210 208 212
rect 211 210 213 212
rect 216 210 218 212
rect 221 210 223 212
rect 226 210 228 212
rect 231 210 233 212
rect 236 210 238 212
rect 241 210 243 212
rect 246 210 248 212
rect 251 210 253 212
rect 256 210 258 212
rect 261 210 263 212
rect 266 210 268 212
rect 271 210 273 212
rect 276 210 278 212
rect 281 210 283 212
rect 286 210 288 212
rect 291 210 293 212
rect 296 210 298 212
rect 301 210 303 212
rect 306 210 308 212
rect 311 210 313 212
rect 318 211 320 213
rect 333 210 335 212
rect 338 210 340 212
rect 351 209 353 211
rect 356 209 358 211
rect 20 205 22 207
rect 25 205 27 207
rect 40 206 42 208
rect 47 205 49 207
rect 52 205 54 207
rect 57 205 59 207
rect 62 205 64 207
rect 67 205 69 207
rect 72 205 74 207
rect 77 205 79 207
rect 82 205 84 207
rect 87 205 89 207
rect 92 205 94 207
rect 97 205 99 207
rect 102 205 104 207
rect 107 205 109 207
rect 112 205 114 207
rect 117 205 119 207
rect 122 205 124 207
rect 127 205 129 207
rect 132 205 134 207
rect 137 205 139 207
rect 142 205 144 207
rect 147 205 149 207
rect 152 205 154 207
rect 162 206 164 208
rect 177 205 179 207
rect 182 205 184 207
rect 196 206 198 208
rect 206 205 208 207
rect 211 205 213 207
rect 216 205 218 207
rect 221 205 223 207
rect 226 205 228 207
rect 231 205 233 207
rect 236 205 238 207
rect 241 205 243 207
rect 246 205 248 207
rect 251 205 253 207
rect 256 205 258 207
rect 261 205 263 207
rect 266 205 268 207
rect 271 205 273 207
rect 276 205 278 207
rect 281 205 283 207
rect 286 205 288 207
rect 291 205 293 207
rect 296 205 298 207
rect 301 205 303 207
rect 306 205 308 207
rect 311 205 313 207
rect 318 206 320 208
rect 333 205 335 207
rect 338 205 340 207
rect 2 201 4 203
rect 7 201 9 203
rect 20 200 22 202
rect 25 200 27 202
rect 40 201 42 203
rect 47 200 49 202
rect 52 200 54 202
rect 57 200 59 202
rect 62 200 64 202
rect 67 200 69 202
rect 72 200 74 202
rect 77 200 79 202
rect 82 200 84 202
rect 87 200 89 202
rect 92 200 94 202
rect 97 200 99 202
rect 102 200 104 202
rect 107 200 109 202
rect 112 200 114 202
rect 117 200 119 202
rect 122 200 124 202
rect 127 200 129 202
rect 132 200 134 202
rect 137 200 139 202
rect 142 200 144 202
rect 147 200 149 202
rect 152 200 154 202
rect 162 201 164 203
rect 177 200 179 202
rect 182 200 184 202
rect 196 201 198 203
rect 206 200 208 202
rect 211 200 213 202
rect 216 200 218 202
rect 221 200 223 202
rect 226 200 228 202
rect 231 200 233 202
rect 236 200 238 202
rect 241 200 243 202
rect 246 200 248 202
rect 251 200 253 202
rect 256 200 258 202
rect 261 200 263 202
rect 266 200 268 202
rect 271 200 273 202
rect 276 200 278 202
rect 281 200 283 202
rect 286 200 288 202
rect 291 200 293 202
rect 296 200 298 202
rect 301 200 303 202
rect 306 200 308 202
rect 311 200 313 202
rect 318 201 320 203
rect 333 200 335 202
rect 338 200 340 202
rect 351 201 353 203
rect 356 201 358 203
rect 20 195 22 197
rect 25 195 27 197
rect 40 196 42 198
rect 47 195 49 197
rect 52 195 54 197
rect 57 195 59 197
rect 62 195 64 197
rect 67 195 69 197
rect 72 195 74 197
rect 77 195 79 197
rect 82 195 84 197
rect 87 195 89 197
rect 92 195 94 197
rect 97 195 99 197
rect 102 195 104 197
rect 107 195 109 197
rect 112 195 114 197
rect 117 195 119 197
rect 122 195 124 197
rect 127 195 129 197
rect 132 195 134 197
rect 137 195 139 197
rect 142 195 144 197
rect 147 195 149 197
rect 152 195 154 197
rect 162 196 164 198
rect 177 195 179 197
rect 182 195 184 197
rect 196 196 198 198
rect 206 195 208 197
rect 211 195 213 197
rect 216 195 218 197
rect 221 195 223 197
rect 226 195 228 197
rect 231 195 233 197
rect 236 195 238 197
rect 241 195 243 197
rect 246 195 248 197
rect 251 195 253 197
rect 256 195 258 197
rect 261 195 263 197
rect 266 195 268 197
rect 271 195 273 197
rect 276 195 278 197
rect 281 195 283 197
rect 286 195 288 197
rect 291 195 293 197
rect 296 195 298 197
rect 301 195 303 197
rect 306 195 308 197
rect 311 195 313 197
rect 318 196 320 198
rect 333 195 335 197
rect 338 195 340 197
rect 2 193 4 195
rect 7 193 9 195
rect 351 193 353 195
rect 356 193 358 195
rect 20 190 22 192
rect 25 190 27 192
rect 40 191 42 193
rect 47 190 49 192
rect 52 190 54 192
rect 57 190 59 192
rect 62 190 64 192
rect 67 190 69 192
rect 72 190 74 192
rect 77 190 79 192
rect 82 190 84 192
rect 87 190 89 192
rect 92 190 94 192
rect 97 190 99 192
rect 102 190 104 192
rect 107 190 109 192
rect 112 190 114 192
rect 117 190 119 192
rect 122 190 124 192
rect 127 190 129 192
rect 132 190 134 192
rect 137 190 139 192
rect 142 190 144 192
rect 147 190 149 192
rect 152 190 154 192
rect 162 191 164 193
rect 177 190 179 192
rect 182 190 184 192
rect 196 191 198 193
rect 206 190 208 192
rect 211 190 213 192
rect 216 190 218 192
rect 221 190 223 192
rect 226 190 228 192
rect 231 190 233 192
rect 236 190 238 192
rect 241 190 243 192
rect 246 190 248 192
rect 251 190 253 192
rect 256 190 258 192
rect 261 190 263 192
rect 266 190 268 192
rect 271 190 273 192
rect 276 190 278 192
rect 281 190 283 192
rect 286 190 288 192
rect 291 190 293 192
rect 296 190 298 192
rect 301 190 303 192
rect 306 190 308 192
rect 311 190 313 192
rect 318 191 320 193
rect 333 190 335 192
rect 338 190 340 192
rect 2 185 4 187
rect 7 185 9 187
rect 20 185 22 187
rect 25 185 27 187
rect 40 186 42 188
rect 47 185 49 187
rect 52 185 54 187
rect 57 185 59 187
rect 62 185 64 187
rect 67 185 69 187
rect 72 185 74 187
rect 77 185 79 187
rect 82 185 84 187
rect 87 185 89 187
rect 92 185 94 187
rect 97 185 99 187
rect 102 185 104 187
rect 107 185 109 187
rect 112 185 114 187
rect 117 185 119 187
rect 122 185 124 187
rect 127 185 129 187
rect 132 185 134 187
rect 137 185 139 187
rect 142 185 144 187
rect 147 185 149 187
rect 152 185 154 187
rect 162 186 164 188
rect 177 185 179 187
rect 182 185 184 187
rect 196 186 198 188
rect 206 185 208 187
rect 211 185 213 187
rect 216 185 218 187
rect 221 185 223 187
rect 226 185 228 187
rect 231 185 233 187
rect 236 185 238 187
rect 241 185 243 187
rect 246 185 248 187
rect 251 185 253 187
rect 256 185 258 187
rect 261 185 263 187
rect 266 185 268 187
rect 271 185 273 187
rect 276 185 278 187
rect 281 185 283 187
rect 286 185 288 187
rect 291 185 293 187
rect 296 185 298 187
rect 301 185 303 187
rect 306 185 308 187
rect 311 185 313 187
rect 318 186 320 188
rect 333 185 335 187
rect 338 185 340 187
rect 351 185 353 187
rect 356 185 358 187
rect 20 180 22 182
rect 25 180 27 182
rect 40 181 42 183
rect 47 180 49 182
rect 52 180 54 182
rect 57 180 59 182
rect 62 180 64 182
rect 67 180 69 182
rect 72 180 74 182
rect 77 180 79 182
rect 82 180 84 182
rect 87 180 89 182
rect 92 180 94 182
rect 97 180 99 182
rect 102 180 104 182
rect 107 180 109 182
rect 112 180 114 182
rect 117 180 119 182
rect 122 180 124 182
rect 127 180 129 182
rect 132 180 134 182
rect 137 180 139 182
rect 142 180 144 182
rect 147 180 149 182
rect 152 180 154 182
rect 162 181 164 183
rect 177 180 179 182
rect 182 180 184 182
rect 196 181 198 183
rect 206 180 208 182
rect 211 180 213 182
rect 216 180 218 182
rect 221 180 223 182
rect 226 180 228 182
rect 231 180 233 182
rect 236 180 238 182
rect 241 180 243 182
rect 246 180 248 182
rect 251 180 253 182
rect 256 180 258 182
rect 261 180 263 182
rect 266 180 268 182
rect 271 180 273 182
rect 276 180 278 182
rect 281 180 283 182
rect 286 180 288 182
rect 291 180 293 182
rect 296 180 298 182
rect 301 180 303 182
rect 306 180 308 182
rect 311 180 313 182
rect 318 181 320 183
rect 333 180 335 182
rect 338 180 340 182
rect 2 177 4 179
rect 7 177 9 179
rect 20 175 22 177
rect 25 175 27 177
rect 40 176 42 178
rect 47 175 49 177
rect 52 175 54 177
rect 57 175 59 177
rect 62 175 64 177
rect 67 175 69 177
rect 72 175 74 177
rect 77 175 79 177
rect 82 175 84 177
rect 87 175 89 177
rect 92 175 94 177
rect 97 175 99 177
rect 102 175 104 177
rect 107 175 109 177
rect 112 175 114 177
rect 117 175 119 177
rect 122 175 124 177
rect 127 175 129 177
rect 132 175 134 177
rect 137 175 139 177
rect 142 175 144 177
rect 147 175 149 177
rect 152 175 154 177
rect 162 176 164 178
rect 177 175 179 177
rect 182 175 184 177
rect 196 176 198 178
rect 206 175 208 177
rect 211 175 213 177
rect 216 175 218 177
rect 221 175 223 177
rect 226 175 228 177
rect 231 175 233 177
rect 236 175 238 177
rect 241 175 243 177
rect 246 175 248 177
rect 251 175 253 177
rect 256 175 258 177
rect 261 175 263 177
rect 266 175 268 177
rect 271 175 273 177
rect 276 175 278 177
rect 281 175 283 177
rect 286 175 288 177
rect 291 175 293 177
rect 296 175 298 177
rect 301 175 303 177
rect 306 175 308 177
rect 311 175 313 177
rect 318 176 320 178
rect 351 177 353 179
rect 356 177 358 179
rect 333 175 335 177
rect 338 175 340 177
rect 2 169 4 171
rect 7 169 9 171
rect 20 170 22 172
rect 25 170 27 172
rect 40 171 42 173
rect 162 171 164 173
rect 177 170 179 172
rect 182 170 184 172
rect 196 171 198 173
rect 318 171 320 173
rect 333 170 335 172
rect 338 170 340 172
rect 351 169 353 171
rect 356 169 358 171
rect 51 165 53 167
rect 61 165 63 167
rect 71 165 73 167
rect 81 165 83 167
rect 91 165 93 167
rect 101 165 103 167
rect 154 165 156 167
rect 204 165 206 167
rect 257 165 259 167
rect 267 165 269 167
rect 277 165 279 167
rect 287 165 289 167
rect 297 165 299 167
rect 307 165 309 167
rect 2 161 4 163
rect 7 161 9 163
rect 51 160 53 162
rect 61 160 63 162
rect 71 160 73 162
rect 81 160 83 162
rect 91 160 93 162
rect 101 160 103 162
rect 154 160 156 162
rect 204 160 206 162
rect 257 160 259 162
rect 267 160 269 162
rect 277 160 279 162
rect 287 160 289 162
rect 297 160 299 162
rect 307 160 309 162
rect 351 161 353 163
rect 356 161 358 163
rect 51 155 53 157
rect 61 155 63 157
rect 71 155 73 157
rect 81 155 83 157
rect 91 155 93 157
rect 101 155 103 157
rect 154 155 156 157
rect 204 155 206 157
rect 257 155 259 157
rect 267 155 269 157
rect 277 155 279 157
rect 287 155 289 157
rect 297 155 299 157
rect 307 155 309 157
rect 2 153 4 155
rect 7 153 9 155
rect 351 153 353 155
rect 356 153 358 155
rect 2 145 4 147
rect 7 145 9 147
rect 351 145 353 147
rect 356 145 358 147
rect 9 137 11 139
rect 17 137 19 139
rect 25 137 27 139
rect 49 137 51 139
rect 57 137 59 139
rect 65 137 67 139
rect 73 137 75 139
rect 81 137 83 139
rect 89 137 91 139
rect 97 137 99 139
rect 105 137 107 139
rect 153 137 155 139
rect 177 137 179 139
rect 205 137 207 139
rect 253 137 255 139
rect 261 137 263 139
rect 269 137 271 139
rect 277 137 279 139
rect 285 137 287 139
rect 293 137 295 139
rect 301 137 303 139
rect 309 137 311 139
rect 333 137 335 139
rect 341 137 343 139
rect 349 137 351 139
rect 9 132 11 134
rect 17 132 19 134
rect 25 132 27 134
rect 49 132 51 134
rect 57 132 59 134
rect 65 132 67 134
rect 73 132 75 134
rect 81 132 83 134
rect 89 132 91 134
rect 97 132 99 134
rect 105 132 107 134
rect 153 132 155 134
rect 177 132 179 134
rect 205 132 207 134
rect 253 132 255 134
rect 261 132 263 134
rect 269 132 271 134
rect 277 132 279 134
rect 285 132 287 134
rect 293 132 295 134
rect 301 132 303 134
rect 309 132 311 134
rect 333 132 335 134
rect 341 132 343 134
rect 349 132 351 134
rect 9 120 11 122
rect 17 120 19 122
rect 25 120 27 122
rect 49 120 51 122
rect 57 120 59 122
rect 65 120 67 122
rect 73 120 75 122
rect 81 120 83 122
rect 89 120 91 122
rect 97 120 99 122
rect 105 120 107 122
rect 113 120 115 122
rect 153 120 155 122
rect 177 120 179 122
rect 205 120 207 122
rect 245 120 247 122
rect 253 120 255 122
rect 261 120 263 122
rect 269 120 271 122
rect 277 120 279 122
rect 285 120 287 122
rect 293 120 295 122
rect 301 120 303 122
rect 309 120 311 122
rect 333 120 335 122
rect 341 120 343 122
rect 349 120 351 122
rect 9 115 11 117
rect 17 115 19 117
rect 25 115 27 117
rect 49 115 51 117
rect 57 115 59 117
rect 65 115 67 117
rect 73 115 75 117
rect 81 115 83 117
rect 89 115 91 117
rect 97 115 99 117
rect 105 115 107 117
rect 113 115 115 117
rect 153 115 155 117
rect 177 115 179 117
rect 205 115 207 117
rect 245 115 247 117
rect 253 115 255 117
rect 261 115 263 117
rect 269 115 271 117
rect 277 115 279 117
rect 285 115 287 117
rect 293 115 295 117
rect 301 115 303 117
rect 309 115 311 117
rect 333 115 335 117
rect 341 115 343 117
rect 349 115 351 117
rect 2 107 4 109
rect 7 107 9 109
rect 351 107 353 109
rect 356 107 358 109
rect 2 102 4 104
rect 7 102 9 104
rect 351 102 353 104
rect 356 102 358 104
rect 2 97 4 99
rect 7 97 9 99
rect 351 97 353 99
rect 356 97 358 99
rect 2 92 4 94
rect 7 92 9 94
rect 351 92 353 94
rect 356 92 358 94
rect 2 87 4 89
rect 7 87 9 89
rect 34 88 36 90
rect 39 88 41 90
rect 44 88 46 90
rect 49 88 51 90
rect 54 88 56 90
rect 59 88 61 90
rect 64 88 66 90
rect 69 88 71 90
rect 289 88 291 90
rect 294 88 296 90
rect 299 88 301 90
rect 304 88 306 90
rect 309 88 311 90
rect 314 88 316 90
rect 319 88 321 90
rect 324 88 326 90
rect 351 87 353 89
rect 356 87 358 89
rect 2 82 4 84
rect 7 82 9 84
rect 351 82 353 84
rect 356 82 358 84
rect 30 80 32 82
rect 35 80 37 82
rect 40 80 42 82
rect 45 80 47 82
rect 50 80 52 82
rect 55 80 57 82
rect 303 80 305 82
rect 308 80 310 82
rect 313 80 315 82
rect 318 80 320 82
rect 323 80 325 82
rect 328 80 330 82
rect 2 77 4 79
rect 7 77 9 79
rect 24 77 26 79
rect 86 78 88 80
rect 91 78 93 80
rect 96 78 98 80
rect 101 78 103 80
rect 106 78 108 80
rect 111 78 113 80
rect 116 78 118 80
rect 121 78 123 80
rect 126 78 128 80
rect 131 78 133 80
rect 136 78 138 80
rect 141 78 143 80
rect 146 78 148 80
rect 151 78 153 80
rect 156 78 158 80
rect 161 78 163 80
rect 166 78 168 80
rect 171 78 173 80
rect 176 78 178 80
rect 181 78 183 80
rect 186 78 188 80
rect 191 78 193 80
rect 196 78 198 80
rect 201 78 203 80
rect 206 78 208 80
rect 211 78 213 80
rect 216 78 218 80
rect 221 78 223 80
rect 226 78 228 80
rect 231 78 233 80
rect 236 78 238 80
rect 241 78 243 80
rect 246 78 248 80
rect 251 78 253 80
rect 256 78 258 80
rect 261 78 263 80
rect 266 78 268 80
rect 271 78 273 80
rect 334 77 336 79
rect 351 77 353 79
rect 356 77 358 79
rect 2 72 4 74
rect 7 72 9 74
rect 24 72 26 74
rect 49 72 51 74
rect 54 72 56 74
rect 59 72 61 74
rect 64 72 66 74
rect 69 72 71 74
rect 86 73 88 75
rect 91 73 93 75
rect 96 73 98 75
rect 101 73 103 75
rect 106 73 108 75
rect 111 73 113 75
rect 116 73 118 75
rect 121 73 123 75
rect 126 73 128 75
rect 131 73 133 75
rect 136 73 138 75
rect 141 73 143 75
rect 146 73 148 75
rect 151 73 153 75
rect 156 73 158 75
rect 161 73 163 75
rect 166 73 168 75
rect 171 73 173 75
rect 176 73 178 75
rect 181 73 183 75
rect 186 73 188 75
rect 191 73 193 75
rect 196 73 198 75
rect 201 73 203 75
rect 206 73 208 75
rect 211 73 213 75
rect 216 73 218 75
rect 221 73 223 75
rect 226 73 228 75
rect 231 73 233 75
rect 236 73 238 75
rect 241 73 243 75
rect 246 73 248 75
rect 251 73 253 75
rect 256 73 258 75
rect 261 73 263 75
rect 266 73 268 75
rect 271 73 273 75
rect 289 72 291 74
rect 294 72 296 74
rect 299 72 301 74
rect 304 72 306 74
rect 309 72 311 74
rect 334 72 336 74
rect 351 72 353 74
rect 356 72 358 74
rect 2 67 4 69
rect 7 67 9 69
rect 24 67 26 69
rect 334 67 336 69
rect 351 67 353 69
rect 356 67 358 69
rect 30 64 32 66
rect 35 64 37 66
rect 40 64 42 66
rect 45 64 47 66
rect 50 64 52 66
rect 55 64 57 66
rect 303 64 305 66
rect 308 64 310 66
rect 313 64 315 66
rect 318 64 320 66
rect 323 64 325 66
rect 328 64 330 66
rect 2 62 4 64
rect 7 62 9 64
rect 24 62 26 64
rect 334 62 336 64
rect 351 62 353 64
rect 356 62 358 64
rect 2 57 4 59
rect 7 57 9 59
rect 24 57 26 59
rect 49 56 51 58
rect 54 56 56 58
rect 59 56 61 58
rect 64 56 66 58
rect 69 56 71 58
rect 289 56 291 58
rect 294 56 296 58
rect 299 56 301 58
rect 304 56 306 58
rect 309 56 311 58
rect 334 57 336 59
rect 351 57 353 59
rect 356 57 358 59
rect 2 52 4 54
rect 7 52 9 54
rect 24 52 26 54
rect 334 52 336 54
rect 351 52 353 54
rect 356 52 358 54
rect 2 47 4 49
rect 7 47 9 49
rect 24 47 26 49
rect 30 48 32 50
rect 35 48 37 50
rect 40 48 42 50
rect 45 48 47 50
rect 50 48 52 50
rect 55 48 57 50
rect 303 48 305 50
rect 308 48 310 50
rect 313 48 315 50
rect 318 48 320 50
rect 323 48 325 50
rect 328 48 330 50
rect 334 47 336 49
rect 351 47 353 49
rect 356 47 358 49
rect 2 42 4 44
rect 7 42 9 44
rect 24 42 26 44
rect 86 43 88 45
rect 91 43 93 45
rect 96 43 98 45
rect 101 43 103 45
rect 106 43 108 45
rect 111 43 113 45
rect 116 43 118 45
rect 121 43 123 45
rect 126 43 128 45
rect 131 43 133 45
rect 136 43 138 45
rect 141 43 143 45
rect 146 43 148 45
rect 151 43 153 45
rect 156 43 158 45
rect 161 43 163 45
rect 166 43 168 45
rect 171 43 173 45
rect 176 43 178 45
rect 181 43 183 45
rect 186 43 188 45
rect 191 43 193 45
rect 196 43 198 45
rect 201 43 203 45
rect 206 43 208 45
rect 211 43 213 45
rect 216 43 218 45
rect 221 43 223 45
rect 226 43 228 45
rect 231 43 233 45
rect 236 43 238 45
rect 241 43 243 45
rect 246 43 248 45
rect 251 43 253 45
rect 256 43 258 45
rect 261 43 263 45
rect 266 43 268 45
rect 271 43 273 45
rect 276 43 278 45
rect 334 42 336 44
rect 351 42 353 44
rect 356 42 358 44
rect 49 40 51 42
rect 54 40 56 42
rect 59 40 61 42
rect 64 40 66 42
rect 69 40 71 42
rect 289 40 291 42
rect 294 40 296 42
rect 299 40 301 42
rect 304 40 306 42
rect 309 40 311 42
rect 2 37 4 39
rect 7 37 9 39
rect 24 37 26 39
rect 86 38 88 40
rect 91 38 93 40
rect 96 38 98 40
rect 101 38 103 40
rect 106 38 108 40
rect 111 38 113 40
rect 116 38 118 40
rect 121 38 123 40
rect 126 38 128 40
rect 131 38 133 40
rect 136 38 138 40
rect 141 38 143 40
rect 146 38 148 40
rect 151 38 153 40
rect 156 38 158 40
rect 161 38 163 40
rect 166 38 168 40
rect 171 38 173 40
rect 176 38 178 40
rect 181 38 183 40
rect 186 38 188 40
rect 191 38 193 40
rect 196 38 198 40
rect 201 38 203 40
rect 206 38 208 40
rect 211 38 213 40
rect 216 38 218 40
rect 221 38 223 40
rect 226 38 228 40
rect 231 38 233 40
rect 236 38 238 40
rect 241 38 243 40
rect 246 38 248 40
rect 251 38 253 40
rect 256 38 258 40
rect 261 38 263 40
rect 266 38 268 40
rect 271 38 273 40
rect 276 38 278 40
rect 334 37 336 39
rect 351 37 353 39
rect 356 37 358 39
rect 2 32 4 34
rect 7 32 9 34
rect 24 32 26 34
rect 30 32 32 34
rect 35 32 37 34
rect 40 32 42 34
rect 45 32 47 34
rect 50 32 52 34
rect 55 32 57 34
rect 303 32 305 34
rect 308 32 310 34
rect 313 32 315 34
rect 318 32 320 34
rect 323 32 325 34
rect 328 32 330 34
rect 334 32 336 34
rect 351 32 353 34
rect 356 32 358 34
rect 2 27 4 29
rect 7 27 9 29
rect 24 27 26 29
rect 334 27 336 29
rect 351 27 353 29
rect 356 27 358 29
rect 49 24 51 26
rect 54 24 56 26
rect 59 24 61 26
rect 64 24 66 26
rect 69 24 71 26
rect 289 24 291 26
rect 294 24 296 26
rect 299 24 301 26
rect 304 24 306 26
rect 309 24 311 26
rect 2 22 4 24
rect 7 22 9 24
rect 24 22 26 24
rect 334 22 336 24
rect 351 22 353 24
rect 356 22 358 24
rect 2 17 4 19
rect 7 17 9 19
rect 24 17 26 19
rect 30 16 32 18
rect 35 16 37 18
rect 40 16 42 18
rect 45 16 47 18
rect 50 16 52 18
rect 55 16 57 18
rect 60 16 62 18
rect 65 16 67 18
rect 293 16 295 18
rect 298 16 300 18
rect 303 16 305 18
rect 308 16 310 18
rect 313 16 315 18
rect 318 16 320 18
rect 323 16 325 18
rect 328 16 330 18
rect 334 17 336 19
rect 351 17 353 19
rect 356 17 358 19
rect 2 12 4 14
rect 7 12 9 14
rect 351 12 353 14
rect 356 12 358 14
rect 7 7 9 9
rect 15 7 17 9
rect 25 7 27 9
rect 33 7 35 9
rect 41 7 43 9
rect 49 7 51 9
rect 57 7 59 9
rect 65 7 67 9
rect 73 7 75 9
rect 81 7 83 9
rect 89 7 91 9
rect 97 7 99 9
rect 105 7 107 9
rect 113 7 115 9
rect 121 7 123 9
rect 129 7 131 9
rect 137 7 139 9
rect 145 7 147 9
rect 153 7 155 9
rect 161 7 163 9
rect 197 7 199 9
rect 205 7 207 9
rect 213 7 215 9
rect 221 7 223 9
rect 229 7 231 9
rect 237 7 239 9
rect 245 7 247 9
rect 253 7 255 9
rect 261 7 263 9
rect 269 7 271 9
rect 277 7 279 9
rect 285 7 287 9
rect 293 7 295 9
rect 301 7 303 9
rect 309 7 311 9
rect 317 7 319 9
rect 325 7 327 9
rect 333 7 335 9
rect 341 7 343 9
rect 351 7 353 9
rect 7 2 9 4
rect 15 2 17 4
rect 25 2 27 4
rect 33 2 35 4
rect 41 2 43 4
rect 49 2 51 4
rect 57 2 59 4
rect 65 2 67 4
rect 73 2 75 4
rect 81 2 83 4
rect 89 2 91 4
rect 97 2 99 4
rect 105 2 107 4
rect 113 2 115 4
rect 121 2 123 4
rect 129 2 131 4
rect 137 2 139 4
rect 145 2 147 4
rect 153 2 155 4
rect 161 2 163 4
rect 197 2 199 4
rect 205 2 207 4
rect 213 2 215 4
rect 221 2 223 4
rect 229 2 231 4
rect 237 2 239 4
rect 245 2 247 4
rect 253 2 255 4
rect 261 2 263 4
rect 269 2 271 4
rect 277 2 279 4
rect 285 2 287 4
rect 293 2 295 4
rect 301 2 303 4
rect 309 2 311 4
rect 317 2 319 4
rect 325 2 327 4
rect 333 2 335 4
rect 341 2 343 4
rect 351 2 353 4
<< metal1 >>
rect 45 767 315 1037
rect 62 757 298 767
rect 72 747 288 757
rect 82 737 278 747
rect 92 727 268 737
rect 102 717 258 727
rect 112 707 248 717
rect 120 704 240 707
rect 0 684 117 695
rect 0 449 11 684
rect 18 656 115 672
rect 18 461 29 656
rect 0 438 29 449
rect 0 421 29 432
rect 32 417 36 653
rect 120 651 143 704
rect 149 684 211 695
rect 168 676 192 680
rect 148 656 164 672
rect 41 612 165 651
rect 39 591 115 607
rect 120 586 143 612
rect 148 591 164 607
rect 41 547 165 586
rect 39 526 115 542
rect 120 521 143 547
rect 148 526 164 542
rect 41 482 165 521
rect 39 461 115 477
rect 39 438 117 449
rect 39 421 117 432
rect 31 408 42 417
rect 0 393 29 404
rect 0 376 29 387
rect 0 141 11 376
rect 18 153 29 364
rect 32 221 36 408
rect 39 393 117 404
rect 39 376 117 387
rect 39 348 115 364
rect 39 299 43 348
rect 120 343 143 482
rect 148 461 164 477
rect 168 457 172 676
rect 175 461 185 672
rect 188 457 192 676
rect 196 656 212 672
rect 217 651 240 704
rect 243 684 360 695
rect 245 656 342 672
rect 195 612 319 651
rect 196 591 212 607
rect 217 586 240 612
rect 245 591 321 607
rect 195 547 319 586
rect 196 526 212 542
rect 217 521 240 547
rect 245 526 321 542
rect 195 482 319 521
rect 196 461 212 477
rect 168 453 192 457
rect 148 438 162 449
rect 148 421 162 432
rect 168 417 172 453
rect 175 438 185 449
rect 175 421 185 432
rect 188 417 192 453
rect 196 438 210 449
rect 196 421 210 432
rect 167 408 193 417
rect 148 393 162 404
rect 148 376 162 387
rect 168 372 172 408
rect 175 393 185 404
rect 175 376 185 387
rect 188 372 192 408
rect 196 393 210 404
rect 196 376 210 387
rect 168 368 192 372
rect 148 348 165 364
rect 46 304 155 343
rect 39 283 115 299
rect 39 234 43 283
rect 120 278 143 304
rect 161 299 165 348
rect 148 283 165 299
rect 46 239 155 278
rect 39 228 115 234
rect 0 130 29 141
rect 0 113 29 124
rect 0 11 11 113
rect 32 109 43 221
rect 49 218 115 228
rect 120 213 143 239
rect 161 234 165 283
rect 148 228 165 234
rect 148 218 157 228
rect 168 221 172 368
rect 46 174 155 213
rect 49 153 115 169
rect 46 130 113 141
rect 46 113 116 124
rect 15 100 108 109
rect 120 100 143 174
rect 147 153 157 169
rect 147 130 157 141
rect 147 113 157 124
rect 161 109 172 221
rect 175 153 185 364
rect 188 256 192 368
rect 195 348 212 364
rect 195 299 199 348
rect 217 343 240 482
rect 245 461 321 477
rect 243 438 321 449
rect 243 421 321 432
rect 324 417 328 653
rect 331 461 342 656
rect 349 449 360 684
rect 331 438 360 449
rect 331 421 360 432
rect 318 408 329 417
rect 243 393 321 404
rect 243 376 321 387
rect 245 348 321 364
rect 205 304 314 343
rect 195 283 212 299
rect 195 264 199 283
rect 217 278 240 304
rect 317 299 321 348
rect 245 283 321 299
rect 176 130 184 141
rect 176 113 184 124
rect 188 109 199 256
rect 205 239 314 278
rect 317 264 321 283
rect 324 256 328 408
rect 331 393 360 404
rect 331 376 360 387
rect 203 218 212 234
rect 217 213 240 239
rect 245 218 311 234
rect 205 174 314 213
rect 203 153 213 169
rect 203 130 213 141
rect 203 113 213 124
rect 152 100 209 109
rect 217 100 240 174
rect 245 153 311 169
rect 248 130 312 141
rect 243 113 312 124
rect 317 109 328 256
rect 331 153 342 364
rect 349 141 360 376
rect 331 130 360 141
rect 331 113 360 124
rect 253 100 345 109
rect 117 97 143 100
rect 111 94 143 97
rect 217 97 243 100
rect 217 94 249 97
rect 105 91 146 94
rect 214 91 255 94
rect 30 87 81 91
rect 99 88 152 91
rect 208 88 261 91
rect 23 79 59 83
rect 23 67 45 79
rect 63 75 81 87
rect 93 85 158 88
rect 202 85 267 88
rect 279 87 330 91
rect 87 82 163 85
rect 197 82 273 85
rect 48 71 81 75
rect 85 71 274 82
rect 279 75 297 87
rect 301 79 337 83
rect 279 71 312 75
rect 23 63 59 67
rect 23 51 45 63
rect 63 59 81 71
rect 48 55 81 59
rect 23 47 59 51
rect 63 47 81 55
rect 279 59 297 71
rect 315 67 337 79
rect 301 63 337 67
rect 279 55 312 59
rect 279 47 297 55
rect 315 51 337 63
rect 301 47 337 51
rect 23 35 45 47
rect 63 43 297 47
rect 48 39 312 43
rect 23 31 59 35
rect 23 19 45 31
rect 63 27 297 39
rect 315 35 337 47
rect 301 31 337 35
rect 48 23 312 27
rect 135 21 225 23
rect 23 11 72 19
rect 147 18 213 21
rect 315 19 337 31
rect 159 15 201 18
rect 0 0 170 11
rect 175 0 187 15
rect 288 11 337 19
rect 349 11 360 113
rect 192 0 360 11
<< metal2 >>
rect 47 769 313 1035
rect 0 684 360 695
rect 0 656 360 672
rect 0 618 360 645
rect 0 591 360 607
rect 0 558 360 585
rect 0 526 360 542
rect 193 525 209 526
rect 0 493 360 520
rect 0 461 360 477
rect 193 460 209 461
rect 0 438 360 449
rect 0 421 360 432
rect 31 408 329 417
rect 0 393 360 404
rect 0 376 360 387
rect 0 348 360 364
rect 0 310 360 337
rect 0 283 360 299
rect 0 250 360 277
rect 0 218 360 234
rect 0 185 360 212
rect 0 153 360 169
rect 0 130 360 141
rect 0 113 360 124
rect 15 100 345 109
rect 0 52 45 78
rect 289 52 360 78
rect 0 0 360 11
<< gv1 >>
rect 59 1021 61 1023
rect 69 1021 71 1023
rect 79 1021 81 1023
rect 89 1021 91 1023
rect 99 1021 101 1023
rect 109 1021 111 1023
rect 119 1021 121 1023
rect 129 1021 131 1023
rect 139 1021 141 1023
rect 149 1021 151 1023
rect 159 1021 161 1023
rect 169 1021 171 1023
rect 179 1021 181 1023
rect 189 1021 191 1023
rect 199 1021 201 1023
rect 209 1021 211 1023
rect 219 1021 221 1023
rect 229 1021 231 1023
rect 239 1021 241 1023
rect 249 1021 251 1023
rect 259 1021 261 1023
rect 269 1021 271 1023
rect 279 1021 281 1023
rect 289 1021 291 1023
rect 299 1021 301 1023
rect 59 1011 61 1013
rect 69 1011 71 1013
rect 79 1011 81 1013
rect 89 1011 91 1013
rect 99 1011 101 1013
rect 109 1011 111 1013
rect 119 1011 121 1013
rect 129 1011 131 1013
rect 139 1011 141 1013
rect 149 1011 151 1013
rect 159 1011 161 1013
rect 169 1011 171 1013
rect 179 1011 181 1013
rect 189 1011 191 1013
rect 199 1011 201 1013
rect 209 1011 211 1013
rect 219 1011 221 1013
rect 229 1011 231 1013
rect 239 1011 241 1013
rect 249 1011 251 1013
rect 259 1011 261 1013
rect 269 1011 271 1013
rect 279 1011 281 1013
rect 289 1011 291 1013
rect 299 1011 301 1013
rect 59 1001 61 1003
rect 69 1001 71 1003
rect 79 1001 81 1003
rect 89 1001 91 1003
rect 99 1001 101 1003
rect 109 1001 111 1003
rect 119 1001 121 1003
rect 129 1001 131 1003
rect 139 1001 141 1003
rect 149 1001 151 1003
rect 159 1001 161 1003
rect 169 1001 171 1003
rect 179 1001 181 1003
rect 189 1001 191 1003
rect 199 1001 201 1003
rect 209 1001 211 1003
rect 219 1001 221 1003
rect 229 1001 231 1003
rect 239 1001 241 1003
rect 249 1001 251 1003
rect 259 1001 261 1003
rect 269 1001 271 1003
rect 279 1001 281 1003
rect 289 1001 291 1003
rect 299 1001 301 1003
rect 59 991 61 993
rect 69 991 71 993
rect 79 991 81 993
rect 89 991 91 993
rect 99 991 101 993
rect 109 991 111 993
rect 119 991 121 993
rect 129 991 131 993
rect 139 991 141 993
rect 149 991 151 993
rect 159 991 161 993
rect 169 991 171 993
rect 179 991 181 993
rect 189 991 191 993
rect 199 991 201 993
rect 209 991 211 993
rect 219 991 221 993
rect 229 991 231 993
rect 239 991 241 993
rect 249 991 251 993
rect 259 991 261 993
rect 269 991 271 993
rect 279 991 281 993
rect 289 991 291 993
rect 299 991 301 993
rect 59 981 61 983
rect 69 981 71 983
rect 79 981 81 983
rect 89 981 91 983
rect 99 981 101 983
rect 109 981 111 983
rect 119 981 121 983
rect 129 981 131 983
rect 139 981 141 983
rect 149 981 151 983
rect 159 981 161 983
rect 169 981 171 983
rect 179 981 181 983
rect 189 981 191 983
rect 199 981 201 983
rect 209 981 211 983
rect 219 981 221 983
rect 229 981 231 983
rect 239 981 241 983
rect 249 981 251 983
rect 259 981 261 983
rect 269 981 271 983
rect 279 981 281 983
rect 289 981 291 983
rect 299 981 301 983
rect 59 971 61 973
rect 69 971 71 973
rect 79 971 81 973
rect 89 971 91 973
rect 99 971 101 973
rect 109 971 111 973
rect 119 971 121 973
rect 129 971 131 973
rect 139 971 141 973
rect 149 971 151 973
rect 159 971 161 973
rect 169 971 171 973
rect 179 971 181 973
rect 189 971 191 973
rect 199 971 201 973
rect 209 971 211 973
rect 219 971 221 973
rect 229 971 231 973
rect 239 971 241 973
rect 249 971 251 973
rect 259 971 261 973
rect 269 971 271 973
rect 279 971 281 973
rect 289 971 291 973
rect 299 971 301 973
rect 59 961 61 963
rect 69 961 71 963
rect 79 961 81 963
rect 89 961 91 963
rect 99 961 101 963
rect 109 961 111 963
rect 119 961 121 963
rect 129 961 131 963
rect 139 961 141 963
rect 149 961 151 963
rect 159 961 161 963
rect 169 961 171 963
rect 179 961 181 963
rect 189 961 191 963
rect 199 961 201 963
rect 209 961 211 963
rect 219 961 221 963
rect 229 961 231 963
rect 239 961 241 963
rect 249 961 251 963
rect 259 961 261 963
rect 269 961 271 963
rect 279 961 281 963
rect 289 961 291 963
rect 299 961 301 963
rect 59 951 61 953
rect 69 951 71 953
rect 79 951 81 953
rect 89 951 91 953
rect 99 951 101 953
rect 109 951 111 953
rect 119 951 121 953
rect 129 951 131 953
rect 139 951 141 953
rect 149 951 151 953
rect 159 951 161 953
rect 169 951 171 953
rect 179 951 181 953
rect 189 951 191 953
rect 199 951 201 953
rect 209 951 211 953
rect 219 951 221 953
rect 229 951 231 953
rect 239 951 241 953
rect 249 951 251 953
rect 259 951 261 953
rect 269 951 271 953
rect 279 951 281 953
rect 289 951 291 953
rect 299 951 301 953
rect 59 941 61 943
rect 69 941 71 943
rect 79 941 81 943
rect 89 941 91 943
rect 99 941 101 943
rect 109 941 111 943
rect 119 941 121 943
rect 129 941 131 943
rect 139 941 141 943
rect 149 941 151 943
rect 159 941 161 943
rect 169 941 171 943
rect 179 941 181 943
rect 189 941 191 943
rect 199 941 201 943
rect 209 941 211 943
rect 219 941 221 943
rect 229 941 231 943
rect 239 941 241 943
rect 249 941 251 943
rect 259 941 261 943
rect 269 941 271 943
rect 279 941 281 943
rect 289 941 291 943
rect 299 941 301 943
rect 59 931 61 933
rect 69 931 71 933
rect 79 931 81 933
rect 89 931 91 933
rect 99 931 101 933
rect 109 931 111 933
rect 119 931 121 933
rect 129 931 131 933
rect 139 931 141 933
rect 149 931 151 933
rect 159 931 161 933
rect 169 931 171 933
rect 179 931 181 933
rect 189 931 191 933
rect 199 931 201 933
rect 209 931 211 933
rect 219 931 221 933
rect 229 931 231 933
rect 239 931 241 933
rect 249 931 251 933
rect 259 931 261 933
rect 269 931 271 933
rect 279 931 281 933
rect 289 931 291 933
rect 299 931 301 933
rect 59 921 61 923
rect 69 921 71 923
rect 79 921 81 923
rect 89 921 91 923
rect 99 921 101 923
rect 109 921 111 923
rect 119 921 121 923
rect 129 921 131 923
rect 139 921 141 923
rect 149 921 151 923
rect 159 921 161 923
rect 169 921 171 923
rect 179 921 181 923
rect 189 921 191 923
rect 199 921 201 923
rect 209 921 211 923
rect 219 921 221 923
rect 229 921 231 923
rect 239 921 241 923
rect 249 921 251 923
rect 259 921 261 923
rect 269 921 271 923
rect 279 921 281 923
rect 289 921 291 923
rect 299 921 301 923
rect 59 911 61 913
rect 69 911 71 913
rect 79 911 81 913
rect 89 911 91 913
rect 99 911 101 913
rect 109 911 111 913
rect 119 911 121 913
rect 129 911 131 913
rect 139 911 141 913
rect 149 911 151 913
rect 159 911 161 913
rect 169 911 171 913
rect 179 911 181 913
rect 189 911 191 913
rect 199 911 201 913
rect 209 911 211 913
rect 219 911 221 913
rect 229 911 231 913
rect 239 911 241 913
rect 249 911 251 913
rect 259 911 261 913
rect 269 911 271 913
rect 279 911 281 913
rect 289 911 291 913
rect 299 911 301 913
rect 59 901 61 903
rect 69 901 71 903
rect 79 901 81 903
rect 89 901 91 903
rect 99 901 101 903
rect 109 901 111 903
rect 119 901 121 903
rect 129 901 131 903
rect 139 901 141 903
rect 149 901 151 903
rect 159 901 161 903
rect 169 901 171 903
rect 179 901 181 903
rect 189 901 191 903
rect 199 901 201 903
rect 209 901 211 903
rect 219 901 221 903
rect 229 901 231 903
rect 239 901 241 903
rect 249 901 251 903
rect 259 901 261 903
rect 269 901 271 903
rect 279 901 281 903
rect 289 901 291 903
rect 299 901 301 903
rect 59 891 61 893
rect 69 891 71 893
rect 79 891 81 893
rect 89 891 91 893
rect 99 891 101 893
rect 109 891 111 893
rect 119 891 121 893
rect 129 891 131 893
rect 139 891 141 893
rect 149 891 151 893
rect 159 891 161 893
rect 169 891 171 893
rect 179 891 181 893
rect 189 891 191 893
rect 199 891 201 893
rect 209 891 211 893
rect 219 891 221 893
rect 229 891 231 893
rect 239 891 241 893
rect 249 891 251 893
rect 259 891 261 893
rect 269 891 271 893
rect 279 891 281 893
rect 289 891 291 893
rect 299 891 301 893
rect 59 881 61 883
rect 69 881 71 883
rect 79 881 81 883
rect 89 881 91 883
rect 99 881 101 883
rect 109 881 111 883
rect 119 881 121 883
rect 129 881 131 883
rect 139 881 141 883
rect 149 881 151 883
rect 159 881 161 883
rect 169 881 171 883
rect 179 881 181 883
rect 189 881 191 883
rect 199 881 201 883
rect 209 881 211 883
rect 219 881 221 883
rect 229 881 231 883
rect 239 881 241 883
rect 249 881 251 883
rect 259 881 261 883
rect 269 881 271 883
rect 279 881 281 883
rect 289 881 291 883
rect 299 881 301 883
rect 59 871 61 873
rect 69 871 71 873
rect 79 871 81 873
rect 89 871 91 873
rect 99 871 101 873
rect 109 871 111 873
rect 119 871 121 873
rect 129 871 131 873
rect 139 871 141 873
rect 149 871 151 873
rect 159 871 161 873
rect 169 871 171 873
rect 179 871 181 873
rect 189 871 191 873
rect 199 871 201 873
rect 209 871 211 873
rect 219 871 221 873
rect 229 871 231 873
rect 239 871 241 873
rect 249 871 251 873
rect 259 871 261 873
rect 269 871 271 873
rect 279 871 281 873
rect 289 871 291 873
rect 299 871 301 873
rect 59 861 61 863
rect 69 861 71 863
rect 79 861 81 863
rect 89 861 91 863
rect 99 861 101 863
rect 109 861 111 863
rect 119 861 121 863
rect 129 861 131 863
rect 139 861 141 863
rect 149 861 151 863
rect 159 861 161 863
rect 169 861 171 863
rect 179 861 181 863
rect 189 861 191 863
rect 199 861 201 863
rect 209 861 211 863
rect 219 861 221 863
rect 229 861 231 863
rect 239 861 241 863
rect 249 861 251 863
rect 259 861 261 863
rect 269 861 271 863
rect 279 861 281 863
rect 289 861 291 863
rect 299 861 301 863
rect 59 851 61 853
rect 69 851 71 853
rect 79 851 81 853
rect 89 851 91 853
rect 99 851 101 853
rect 109 851 111 853
rect 119 851 121 853
rect 129 851 131 853
rect 139 851 141 853
rect 149 851 151 853
rect 159 851 161 853
rect 169 851 171 853
rect 179 851 181 853
rect 189 851 191 853
rect 199 851 201 853
rect 209 851 211 853
rect 219 851 221 853
rect 229 851 231 853
rect 239 851 241 853
rect 249 851 251 853
rect 259 851 261 853
rect 269 851 271 853
rect 279 851 281 853
rect 289 851 291 853
rect 299 851 301 853
rect 59 841 61 843
rect 69 841 71 843
rect 79 841 81 843
rect 89 841 91 843
rect 99 841 101 843
rect 109 841 111 843
rect 119 841 121 843
rect 129 841 131 843
rect 139 841 141 843
rect 149 841 151 843
rect 159 841 161 843
rect 169 841 171 843
rect 179 841 181 843
rect 189 841 191 843
rect 199 841 201 843
rect 209 841 211 843
rect 219 841 221 843
rect 229 841 231 843
rect 239 841 241 843
rect 249 841 251 843
rect 259 841 261 843
rect 269 841 271 843
rect 279 841 281 843
rect 289 841 291 843
rect 299 841 301 843
rect 59 831 61 833
rect 69 831 71 833
rect 79 831 81 833
rect 89 831 91 833
rect 99 831 101 833
rect 109 831 111 833
rect 119 831 121 833
rect 129 831 131 833
rect 139 831 141 833
rect 149 831 151 833
rect 159 831 161 833
rect 169 831 171 833
rect 179 831 181 833
rect 189 831 191 833
rect 199 831 201 833
rect 209 831 211 833
rect 219 831 221 833
rect 229 831 231 833
rect 239 831 241 833
rect 249 831 251 833
rect 259 831 261 833
rect 269 831 271 833
rect 279 831 281 833
rect 289 831 291 833
rect 299 831 301 833
rect 59 821 61 823
rect 69 821 71 823
rect 79 821 81 823
rect 89 821 91 823
rect 99 821 101 823
rect 109 821 111 823
rect 119 821 121 823
rect 129 821 131 823
rect 139 821 141 823
rect 149 821 151 823
rect 159 821 161 823
rect 169 821 171 823
rect 179 821 181 823
rect 189 821 191 823
rect 199 821 201 823
rect 209 821 211 823
rect 219 821 221 823
rect 229 821 231 823
rect 239 821 241 823
rect 249 821 251 823
rect 259 821 261 823
rect 269 821 271 823
rect 279 821 281 823
rect 289 821 291 823
rect 299 821 301 823
rect 59 811 61 813
rect 69 811 71 813
rect 79 811 81 813
rect 89 811 91 813
rect 99 811 101 813
rect 109 811 111 813
rect 119 811 121 813
rect 129 811 131 813
rect 139 811 141 813
rect 149 811 151 813
rect 159 811 161 813
rect 169 811 171 813
rect 179 811 181 813
rect 189 811 191 813
rect 199 811 201 813
rect 209 811 211 813
rect 219 811 221 813
rect 229 811 231 813
rect 239 811 241 813
rect 249 811 251 813
rect 259 811 261 813
rect 269 811 271 813
rect 279 811 281 813
rect 289 811 291 813
rect 299 811 301 813
rect 59 801 61 803
rect 69 801 71 803
rect 79 801 81 803
rect 89 801 91 803
rect 99 801 101 803
rect 109 801 111 803
rect 119 801 121 803
rect 129 801 131 803
rect 139 801 141 803
rect 149 801 151 803
rect 159 801 161 803
rect 169 801 171 803
rect 179 801 181 803
rect 189 801 191 803
rect 199 801 201 803
rect 209 801 211 803
rect 219 801 221 803
rect 229 801 231 803
rect 239 801 241 803
rect 249 801 251 803
rect 259 801 261 803
rect 269 801 271 803
rect 279 801 281 803
rect 289 801 291 803
rect 299 801 301 803
rect 59 791 61 793
rect 69 791 71 793
rect 79 791 81 793
rect 89 791 91 793
rect 99 791 101 793
rect 109 791 111 793
rect 119 791 121 793
rect 129 791 131 793
rect 139 791 141 793
rect 149 791 151 793
rect 159 791 161 793
rect 169 791 171 793
rect 179 791 181 793
rect 189 791 191 793
rect 199 791 201 793
rect 209 791 211 793
rect 219 791 221 793
rect 229 791 231 793
rect 239 791 241 793
rect 249 791 251 793
rect 259 791 261 793
rect 269 791 271 793
rect 279 791 281 793
rect 289 791 291 793
rect 299 791 301 793
rect 59 781 61 783
rect 69 781 71 783
rect 79 781 81 783
rect 89 781 91 783
rect 99 781 101 783
rect 109 781 111 783
rect 119 781 121 783
rect 129 781 131 783
rect 139 781 141 783
rect 149 781 151 783
rect 159 781 161 783
rect 169 781 171 783
rect 179 781 181 783
rect 189 781 191 783
rect 199 781 201 783
rect 209 781 211 783
rect 219 781 221 783
rect 229 781 231 783
rect 239 781 241 783
rect 249 781 251 783
rect 259 781 261 783
rect 269 781 271 783
rect 279 781 281 783
rect 289 781 291 783
rect 299 781 301 783
rect 5 691 7 693
rect 13 691 15 693
rect 21 691 23 693
rect 29 691 31 693
rect 37 691 39 693
rect 45 691 47 693
rect 53 691 55 693
rect 61 691 63 693
rect 69 691 71 693
rect 77 691 79 693
rect 85 691 87 693
rect 93 691 95 693
rect 101 691 103 693
rect 109 691 111 693
rect 155 691 157 693
rect 163 691 165 693
rect 171 691 173 693
rect 179 691 181 693
rect 187 691 189 693
rect 195 691 197 693
rect 203 691 205 693
rect 249 691 251 693
rect 257 691 259 693
rect 265 691 267 693
rect 273 691 275 693
rect 281 691 283 693
rect 289 691 291 693
rect 297 691 299 693
rect 305 691 307 693
rect 313 691 315 693
rect 321 691 323 693
rect 329 691 331 693
rect 337 691 339 693
rect 345 691 347 693
rect 353 691 355 693
rect 5 686 7 688
rect 13 686 15 688
rect 21 686 23 688
rect 29 686 31 688
rect 37 686 39 688
rect 45 686 47 688
rect 53 686 55 688
rect 61 686 63 688
rect 69 686 71 688
rect 77 686 79 688
rect 85 686 87 688
rect 93 686 95 688
rect 101 686 103 688
rect 109 686 111 688
rect 155 686 157 688
rect 163 686 165 688
rect 171 686 173 688
rect 179 686 181 688
rect 187 686 189 688
rect 195 686 197 688
rect 203 686 205 688
rect 249 686 251 688
rect 257 686 259 688
rect 265 686 267 688
rect 273 686 275 688
rect 281 686 283 688
rect 289 686 291 688
rect 297 686 299 688
rect 305 686 307 688
rect 313 686 315 688
rect 321 686 323 688
rect 329 686 331 688
rect 337 686 339 688
rect 345 686 347 688
rect 353 686 355 688
rect 20 668 22 670
rect 25 668 27 670
rect 35 668 37 670
rect 46 668 48 670
rect 56 668 58 670
rect 66 668 68 670
rect 76 668 78 670
rect 86 668 88 670
rect 96 668 98 670
rect 106 668 108 670
rect 155 668 157 670
rect 177 668 179 670
rect 182 668 184 670
rect 203 668 205 670
rect 252 668 254 670
rect 262 668 264 670
rect 272 668 274 670
rect 282 668 284 670
rect 292 668 294 670
rect 302 668 304 670
rect 312 668 314 670
rect 322 668 324 670
rect 332 668 335 670
rect 338 668 340 670
rect 20 663 22 665
rect 25 663 27 665
rect 35 663 37 665
rect 46 663 48 665
rect 56 663 58 665
rect 66 663 68 665
rect 76 663 78 665
rect 86 663 88 665
rect 96 663 98 665
rect 106 663 108 665
rect 155 663 157 665
rect 177 663 179 665
rect 182 663 184 665
rect 203 663 205 665
rect 252 663 254 665
rect 262 663 264 665
rect 272 663 274 665
rect 282 663 284 665
rect 292 663 294 665
rect 302 663 304 665
rect 312 663 314 665
rect 322 663 324 665
rect 333 663 335 665
rect 338 663 340 665
rect 20 658 22 660
rect 25 658 27 660
rect 35 658 37 660
rect 46 658 48 660
rect 56 658 58 660
rect 66 658 68 660
rect 76 658 78 660
rect 86 658 88 660
rect 96 658 98 660
rect 106 658 108 660
rect 155 658 157 660
rect 177 658 179 660
rect 182 658 184 660
rect 203 658 205 660
rect 252 658 254 660
rect 262 658 264 660
rect 272 658 274 660
rect 282 658 284 660
rect 292 658 294 660
rect 302 658 304 660
rect 312 658 314 660
rect 322 658 324 660
rect 333 658 335 660
rect 338 658 340 660
rect 2 642 4 644
rect 7 642 9 644
rect 351 642 353 644
rect 356 642 358 644
rect 2 634 4 636
rect 7 634 9 636
rect 351 634 353 636
rect 356 634 358 636
rect 2 626 4 628
rect 7 626 9 628
rect 351 626 353 628
rect 356 626 358 628
rect 20 603 22 605
rect 25 603 27 605
rect 46 603 48 605
rect 56 603 58 605
rect 66 603 68 605
rect 76 603 78 605
rect 86 603 88 605
rect 96 603 98 605
rect 106 603 108 605
rect 155 603 157 605
rect 177 603 179 605
rect 182 603 184 605
rect 203 603 205 605
rect 252 603 254 605
rect 262 603 264 605
rect 272 603 274 605
rect 282 603 284 605
rect 292 603 294 605
rect 302 603 304 605
rect 312 603 314 605
rect 333 603 335 605
rect 338 603 340 605
rect 20 598 22 600
rect 25 598 27 600
rect 46 598 48 600
rect 56 598 58 600
rect 66 598 68 600
rect 76 598 78 600
rect 86 598 88 600
rect 96 598 98 600
rect 106 598 108 600
rect 155 598 157 600
rect 177 598 179 600
rect 182 598 184 600
rect 203 598 205 600
rect 252 598 254 600
rect 262 598 264 600
rect 272 598 274 600
rect 282 598 284 600
rect 292 598 294 600
rect 302 598 304 600
rect 312 598 314 600
rect 333 598 335 600
rect 338 598 340 600
rect 20 593 22 595
rect 25 593 27 595
rect 46 593 48 595
rect 56 593 58 595
rect 66 593 68 595
rect 76 593 78 595
rect 86 593 88 595
rect 96 593 98 595
rect 106 593 108 595
rect 155 593 157 595
rect 177 593 179 595
rect 182 593 184 595
rect 203 593 205 595
rect 252 593 254 595
rect 262 593 264 595
rect 272 593 274 595
rect 282 593 284 595
rect 292 593 294 595
rect 302 593 304 595
rect 312 593 314 595
rect 333 593 335 595
rect 338 593 340 595
rect 2 578 4 580
rect 7 578 9 580
rect 351 578 353 580
rect 356 578 358 580
rect 2 570 4 572
rect 7 570 9 572
rect 351 570 353 572
rect 356 570 358 572
rect 2 562 4 564
rect 7 562 9 564
rect 351 562 353 564
rect 356 562 358 564
rect 20 538 22 540
rect 25 538 27 540
rect 46 538 48 540
rect 56 538 58 540
rect 66 538 68 540
rect 76 538 78 540
rect 86 538 88 540
rect 96 538 98 540
rect 106 538 108 540
rect 155 538 157 540
rect 177 538 179 540
rect 182 538 184 540
rect 203 538 205 540
rect 252 538 254 540
rect 262 538 264 540
rect 272 538 274 540
rect 282 538 284 540
rect 292 538 294 540
rect 302 538 304 540
rect 312 538 314 540
rect 333 538 335 540
rect 338 538 340 540
rect 20 533 22 535
rect 25 533 27 535
rect 46 533 48 535
rect 56 533 58 535
rect 66 533 68 535
rect 76 533 78 535
rect 86 533 88 535
rect 96 533 98 535
rect 106 533 108 535
rect 155 533 157 535
rect 177 533 179 535
rect 182 533 184 535
rect 203 533 205 535
rect 252 533 254 535
rect 262 533 264 535
rect 272 533 274 535
rect 282 533 284 535
rect 292 533 294 535
rect 302 533 304 535
rect 312 533 314 535
rect 333 533 335 535
rect 338 533 340 535
rect 20 528 22 530
rect 25 528 27 530
rect 46 528 48 530
rect 56 528 58 530
rect 66 528 68 530
rect 76 528 78 530
rect 86 528 88 530
rect 96 528 98 530
rect 106 528 108 530
rect 155 528 157 530
rect 177 528 179 530
rect 182 528 184 530
rect 203 528 205 530
rect 252 528 254 530
rect 262 528 264 530
rect 272 528 274 530
rect 282 528 284 530
rect 292 528 294 530
rect 302 528 304 530
rect 312 528 314 530
rect 333 528 335 530
rect 338 528 340 530
rect 2 513 4 515
rect 7 513 9 515
rect 351 513 353 515
rect 356 513 358 515
rect 2 505 4 507
rect 7 505 9 507
rect 351 505 353 507
rect 356 505 358 507
rect 2 497 4 499
rect 7 497 9 499
rect 351 497 353 499
rect 356 497 358 499
rect 20 473 22 475
rect 25 473 27 475
rect 46 473 48 475
rect 56 473 58 475
rect 66 473 68 475
rect 76 473 78 475
rect 86 473 88 475
rect 96 473 98 475
rect 106 473 108 475
rect 155 473 157 475
rect 177 473 179 475
rect 182 473 184 475
rect 203 473 205 475
rect 252 473 254 475
rect 262 473 264 475
rect 272 473 274 475
rect 282 473 284 475
rect 292 473 294 475
rect 302 473 304 475
rect 312 473 314 475
rect 333 473 335 475
rect 338 473 340 475
rect 20 468 22 470
rect 25 468 27 470
rect 46 468 48 470
rect 56 468 58 470
rect 66 468 68 470
rect 76 468 78 470
rect 86 468 88 470
rect 96 468 98 470
rect 106 468 108 470
rect 155 468 157 470
rect 177 468 179 470
rect 182 468 184 470
rect 203 468 205 470
rect 252 468 254 470
rect 262 468 264 470
rect 272 468 274 470
rect 282 468 284 470
rect 292 468 294 470
rect 302 468 304 470
rect 312 468 314 470
rect 333 468 335 470
rect 338 468 340 470
rect 20 463 22 465
rect 25 463 27 465
rect 46 463 48 465
rect 56 463 58 465
rect 66 463 68 465
rect 76 463 78 465
rect 86 463 88 465
rect 96 463 98 465
rect 106 463 108 465
rect 155 463 157 465
rect 177 463 179 465
rect 182 463 184 465
rect 203 463 205 465
rect 252 463 254 465
rect 262 463 264 465
rect 272 463 274 465
rect 282 463 284 465
rect 292 463 294 465
rect 302 463 304 465
rect 312 463 314 465
rect 333 463 335 465
rect 338 463 340 465
rect 5 445 7 447
rect 13 445 15 447
rect 21 445 23 447
rect 45 445 47 447
rect 53 445 55 447
rect 61 445 63 447
rect 69 445 71 447
rect 77 445 79 447
rect 85 445 87 447
rect 93 445 95 447
rect 101 445 103 447
rect 109 445 111 447
rect 154 445 156 447
rect 177 445 179 447
rect 202 445 204 447
rect 249 445 251 447
rect 257 445 259 447
rect 265 445 267 447
rect 273 445 275 447
rect 281 445 283 447
rect 289 445 291 447
rect 297 445 299 447
rect 305 445 307 447
rect 313 445 315 447
rect 337 445 339 447
rect 345 445 347 447
rect 353 445 355 447
rect 5 440 7 442
rect 13 440 15 442
rect 21 440 23 442
rect 45 440 47 442
rect 53 440 55 442
rect 61 440 63 442
rect 69 440 71 442
rect 77 440 79 442
rect 85 440 87 442
rect 93 440 95 442
rect 101 440 103 442
rect 109 440 111 442
rect 154 440 156 442
rect 177 440 179 442
rect 202 440 204 442
rect 249 440 251 442
rect 257 440 259 442
rect 265 440 267 442
rect 273 440 275 442
rect 281 440 283 442
rect 289 440 291 442
rect 297 440 299 442
rect 305 440 307 442
rect 313 440 315 442
rect 337 440 339 442
rect 345 440 347 442
rect 353 440 355 442
rect 5 428 7 430
rect 13 428 15 430
rect 21 428 23 430
rect 45 428 47 430
rect 53 428 55 430
rect 61 428 63 430
rect 69 428 71 430
rect 77 428 79 430
rect 85 428 87 430
rect 93 428 95 430
rect 101 428 103 430
rect 109 428 111 430
rect 154 428 156 430
rect 177 428 179 430
rect 202 428 204 430
rect 249 428 251 430
rect 257 428 259 430
rect 265 428 267 430
rect 273 428 275 430
rect 281 428 283 430
rect 289 428 291 430
rect 297 428 299 430
rect 305 428 307 430
rect 313 428 315 430
rect 337 428 339 430
rect 345 428 347 430
rect 353 428 355 430
rect 5 423 7 425
rect 13 423 15 425
rect 21 423 23 425
rect 45 423 47 425
rect 53 423 55 425
rect 61 423 63 425
rect 69 423 71 425
rect 77 423 79 425
rect 85 423 87 425
rect 93 423 95 425
rect 101 423 103 425
rect 109 423 111 425
rect 154 423 156 425
rect 177 423 179 425
rect 202 423 204 425
rect 249 423 251 425
rect 257 423 259 425
rect 265 423 267 425
rect 273 423 275 425
rect 281 423 283 425
rect 289 423 291 425
rect 297 423 299 425
rect 305 423 307 425
rect 313 423 315 425
rect 337 423 339 425
rect 345 423 347 425
rect 353 423 355 425
rect 33 414 35 416
rect 38 414 40 416
rect 169 414 171 416
rect 174 414 176 416
rect 179 414 181 416
rect 184 414 186 416
rect 189 414 191 416
rect 320 414 322 416
rect 325 414 327 416
rect 33 409 35 411
rect 38 409 40 411
rect 169 409 171 411
rect 174 409 176 411
rect 179 409 181 411
rect 184 409 186 411
rect 189 409 191 411
rect 320 409 322 411
rect 325 409 327 411
rect 5 400 7 402
rect 13 400 15 402
rect 21 400 23 402
rect 45 400 47 402
rect 53 400 55 402
rect 61 400 63 402
rect 69 400 71 402
rect 77 400 79 402
rect 85 400 87 402
rect 93 400 95 402
rect 101 400 103 402
rect 109 400 111 402
rect 154 400 156 402
rect 177 400 179 402
rect 202 400 204 402
rect 249 400 251 402
rect 257 400 259 402
rect 265 400 267 402
rect 273 400 275 402
rect 281 400 283 402
rect 289 400 291 402
rect 297 400 299 402
rect 305 400 307 402
rect 313 400 315 402
rect 337 400 339 402
rect 345 400 347 402
rect 353 400 355 402
rect 5 395 7 397
rect 13 395 15 397
rect 21 395 23 397
rect 45 395 47 397
rect 53 395 55 397
rect 61 395 63 397
rect 69 395 71 397
rect 77 395 79 397
rect 85 395 87 397
rect 93 395 95 397
rect 101 395 103 397
rect 109 395 111 397
rect 154 395 156 397
rect 177 395 179 397
rect 202 395 204 397
rect 249 395 251 397
rect 257 395 259 397
rect 265 395 267 397
rect 273 395 275 397
rect 281 395 283 397
rect 289 395 291 397
rect 297 395 299 397
rect 305 395 307 397
rect 313 395 315 397
rect 337 395 339 397
rect 345 395 347 397
rect 353 395 355 397
rect 5 383 7 385
rect 13 383 15 385
rect 21 383 23 385
rect 45 383 47 385
rect 53 383 55 385
rect 61 383 63 385
rect 69 383 71 385
rect 77 383 79 385
rect 85 383 87 385
rect 93 383 95 385
rect 101 383 103 385
rect 109 383 111 385
rect 154 383 156 385
rect 177 383 179 385
rect 202 383 204 385
rect 249 383 251 385
rect 257 383 259 385
rect 265 383 267 385
rect 273 383 275 385
rect 281 383 283 385
rect 289 383 291 385
rect 297 383 299 385
rect 305 383 307 385
rect 313 383 315 385
rect 337 383 339 385
rect 345 383 347 385
rect 353 383 355 385
rect 5 378 7 380
rect 13 378 15 380
rect 21 378 23 380
rect 45 378 47 380
rect 53 378 55 380
rect 61 378 63 380
rect 69 378 71 380
rect 77 378 79 380
rect 85 378 87 380
rect 93 378 95 380
rect 101 378 103 380
rect 109 378 111 380
rect 154 378 156 380
rect 177 378 179 380
rect 202 378 204 380
rect 249 378 251 380
rect 257 378 259 380
rect 265 378 267 380
rect 273 378 275 380
rect 281 378 283 380
rect 289 378 291 380
rect 297 378 299 380
rect 305 378 307 380
rect 313 378 315 380
rect 337 378 339 380
rect 345 378 347 380
rect 353 378 355 380
rect 20 360 22 362
rect 25 360 27 362
rect 46 360 48 362
rect 56 360 58 362
rect 66 360 68 362
rect 76 360 78 362
rect 86 360 88 362
rect 96 360 98 362
rect 106 360 108 362
rect 149 360 151 362
rect 154 360 156 362
rect 177 360 179 362
rect 182 360 184 362
rect 204 360 206 362
rect 209 360 211 362
rect 252 360 254 362
rect 262 360 264 362
rect 272 360 274 362
rect 282 360 284 362
rect 292 360 294 362
rect 302 360 304 362
rect 312 360 314 362
rect 333 360 335 362
rect 338 360 340 362
rect 20 355 22 357
rect 25 355 27 357
rect 46 355 48 357
rect 56 355 58 357
rect 66 355 68 357
rect 76 355 78 357
rect 86 355 88 357
rect 96 355 98 357
rect 106 355 108 357
rect 149 355 151 357
rect 154 355 156 357
rect 177 355 179 357
rect 182 355 184 357
rect 204 355 206 357
rect 209 355 211 357
rect 252 355 254 357
rect 262 355 264 357
rect 272 355 274 357
rect 282 355 284 357
rect 292 355 294 357
rect 302 355 304 357
rect 312 355 314 357
rect 333 355 335 357
rect 338 355 340 357
rect 20 350 22 352
rect 25 350 27 352
rect 46 350 48 352
rect 56 350 58 352
rect 66 350 68 352
rect 76 350 78 352
rect 86 350 88 352
rect 96 350 98 352
rect 106 350 108 352
rect 149 350 151 352
rect 154 350 156 352
rect 177 350 179 352
rect 182 350 184 352
rect 204 350 206 352
rect 209 350 211 352
rect 252 350 254 352
rect 262 350 264 352
rect 272 350 274 352
rect 282 350 284 352
rect 292 350 294 352
rect 302 350 304 352
rect 312 350 314 352
rect 333 350 335 352
rect 338 350 340 352
rect 2 334 4 336
rect 7 334 9 336
rect 351 334 353 336
rect 356 334 358 336
rect 2 326 4 328
rect 7 326 9 328
rect 351 326 353 328
rect 356 326 358 328
rect 2 318 4 320
rect 7 318 9 320
rect 351 318 353 320
rect 356 318 358 320
rect 20 295 22 297
rect 25 295 27 297
rect 51 295 53 297
rect 56 295 58 297
rect 61 295 63 297
rect 66 295 68 297
rect 71 295 73 297
rect 76 295 78 297
rect 81 295 83 297
rect 86 295 88 297
rect 91 295 93 297
rect 96 295 98 297
rect 101 295 103 297
rect 106 295 108 297
rect 111 295 113 297
rect 149 295 151 297
rect 154 295 156 297
rect 177 295 179 297
rect 182 295 184 297
rect 204 295 206 297
rect 209 295 211 297
rect 247 295 249 297
rect 252 295 254 297
rect 257 295 259 297
rect 262 295 264 297
rect 267 295 269 297
rect 272 295 274 297
rect 277 295 279 297
rect 282 295 284 297
rect 287 295 289 297
rect 292 295 294 297
rect 297 295 299 297
rect 302 295 304 297
rect 307 295 309 297
rect 333 295 335 297
rect 338 295 340 297
rect 20 290 22 292
rect 25 290 27 292
rect 51 290 53 292
rect 56 290 58 292
rect 61 290 63 292
rect 66 290 68 292
rect 71 290 73 292
rect 76 290 78 292
rect 81 290 83 292
rect 86 290 88 292
rect 91 290 93 292
rect 96 290 98 292
rect 101 290 103 292
rect 106 290 108 292
rect 111 290 113 292
rect 149 290 151 292
rect 154 290 156 292
rect 177 290 179 292
rect 182 290 184 292
rect 204 290 206 292
rect 209 290 211 292
rect 247 290 249 292
rect 252 290 254 292
rect 257 290 259 292
rect 262 290 264 292
rect 267 290 269 292
rect 272 290 274 292
rect 277 290 279 292
rect 282 290 284 292
rect 287 290 289 292
rect 292 290 294 292
rect 297 290 299 292
rect 302 290 304 292
rect 307 290 309 292
rect 333 290 335 292
rect 338 290 340 292
rect 20 285 22 287
rect 25 285 27 287
rect 51 285 53 287
rect 56 285 58 287
rect 61 285 63 287
rect 66 285 68 287
rect 71 285 73 287
rect 76 285 78 287
rect 81 285 83 287
rect 86 285 88 287
rect 91 285 93 287
rect 96 285 98 287
rect 101 285 103 287
rect 106 285 108 287
rect 111 285 113 287
rect 149 285 151 287
rect 154 285 156 287
rect 177 285 179 287
rect 182 285 184 287
rect 204 285 206 287
rect 209 285 211 287
rect 247 285 249 287
rect 252 285 254 287
rect 257 285 259 287
rect 262 285 264 287
rect 267 285 269 287
rect 272 285 274 287
rect 277 285 279 287
rect 282 285 284 287
rect 287 285 289 287
rect 292 285 294 287
rect 297 285 299 287
rect 302 285 304 287
rect 307 285 309 287
rect 333 285 335 287
rect 338 285 340 287
rect 2 270 4 272
rect 7 270 9 272
rect 351 270 353 272
rect 356 270 358 272
rect 2 262 4 264
rect 7 262 9 264
rect 351 262 353 264
rect 356 262 358 264
rect 2 254 4 256
rect 7 254 9 256
rect 351 254 353 256
rect 356 254 358 256
rect 20 230 22 232
rect 25 230 27 232
rect 51 230 53 232
rect 56 230 58 232
rect 61 230 63 232
rect 66 230 68 232
rect 71 230 73 232
rect 76 230 78 232
rect 81 230 83 232
rect 86 230 88 232
rect 91 230 93 232
rect 96 230 98 232
rect 101 230 103 232
rect 106 230 108 232
rect 111 230 113 232
rect 149 230 151 232
rect 154 230 156 232
rect 177 230 179 232
rect 182 230 184 232
rect 204 230 206 232
rect 209 230 211 232
rect 247 230 249 232
rect 252 230 254 232
rect 257 230 259 232
rect 262 230 264 232
rect 267 230 269 232
rect 272 230 274 232
rect 277 230 279 232
rect 282 230 284 232
rect 287 230 289 232
rect 292 230 294 232
rect 297 230 299 232
rect 302 230 304 232
rect 307 230 309 232
rect 333 230 335 232
rect 338 230 340 232
rect 20 225 22 227
rect 25 225 27 227
rect 51 225 53 227
rect 56 225 58 227
rect 61 225 63 227
rect 66 225 68 227
rect 71 225 73 227
rect 76 225 78 227
rect 81 225 83 227
rect 86 225 88 227
rect 91 225 93 227
rect 96 225 98 227
rect 101 225 103 227
rect 106 225 108 227
rect 111 225 113 227
rect 149 225 151 227
rect 154 225 156 227
rect 177 225 179 227
rect 182 225 184 227
rect 204 225 206 227
rect 209 225 211 227
rect 247 225 249 227
rect 252 225 254 227
rect 257 225 259 227
rect 262 225 264 227
rect 267 225 269 227
rect 272 225 274 227
rect 277 225 279 227
rect 282 225 284 227
rect 287 225 289 227
rect 292 225 294 227
rect 297 225 299 227
rect 302 225 304 227
rect 307 225 309 227
rect 333 225 335 227
rect 338 225 340 227
rect 20 220 22 222
rect 25 220 27 222
rect 51 220 53 222
rect 56 220 58 222
rect 61 220 63 222
rect 66 220 68 222
rect 71 220 73 222
rect 76 220 78 222
rect 81 220 83 222
rect 86 220 88 222
rect 91 220 93 222
rect 96 220 98 222
rect 101 220 103 222
rect 106 220 108 222
rect 111 220 113 222
rect 149 220 151 222
rect 154 220 156 222
rect 177 220 179 222
rect 182 220 184 222
rect 204 220 206 222
rect 209 220 211 222
rect 247 220 249 222
rect 252 220 254 222
rect 257 220 259 222
rect 262 220 264 222
rect 267 220 269 222
rect 272 220 274 222
rect 277 220 279 222
rect 282 220 284 222
rect 287 220 289 222
rect 292 220 294 222
rect 297 220 299 222
rect 302 220 304 222
rect 307 220 309 222
rect 333 220 335 222
rect 338 220 340 222
rect 2 205 4 207
rect 7 205 9 207
rect 351 205 353 207
rect 356 205 358 207
rect 2 197 4 199
rect 7 197 9 199
rect 351 197 353 199
rect 356 197 358 199
rect 2 189 4 191
rect 7 189 9 191
rect 351 189 353 191
rect 356 189 358 191
rect 20 165 22 167
rect 25 165 27 167
rect 51 165 53 167
rect 56 165 58 167
rect 61 165 63 167
rect 66 165 68 167
rect 71 165 73 167
rect 76 165 78 167
rect 81 165 83 167
rect 86 165 88 167
rect 91 165 93 167
rect 96 165 98 167
rect 101 165 103 167
rect 106 165 108 167
rect 111 165 113 167
rect 149 165 151 167
rect 154 165 156 167
rect 177 165 179 167
rect 182 165 184 167
rect 204 165 206 167
rect 209 165 211 167
rect 247 165 249 167
rect 252 165 254 167
rect 257 165 259 167
rect 262 165 264 167
rect 267 165 269 167
rect 272 165 274 167
rect 277 165 279 167
rect 282 165 284 167
rect 287 165 289 167
rect 292 165 294 167
rect 297 165 299 167
rect 302 165 304 167
rect 307 165 309 167
rect 333 165 335 167
rect 338 165 340 167
rect 20 160 22 162
rect 25 160 27 162
rect 51 160 53 162
rect 56 160 58 162
rect 61 160 63 162
rect 66 160 68 162
rect 71 160 73 162
rect 76 160 78 162
rect 81 160 83 162
rect 86 160 88 162
rect 91 160 93 162
rect 96 160 98 162
rect 101 160 103 162
rect 106 160 108 162
rect 111 160 113 162
rect 149 160 151 162
rect 154 160 156 162
rect 177 160 179 162
rect 182 160 184 162
rect 204 160 206 162
rect 209 160 211 162
rect 247 160 249 162
rect 252 160 254 162
rect 257 160 259 162
rect 262 160 264 162
rect 267 160 269 162
rect 272 160 274 162
rect 277 160 279 162
rect 282 160 284 162
rect 287 160 289 162
rect 292 160 294 162
rect 297 160 299 162
rect 302 160 304 162
rect 307 160 309 162
rect 333 160 335 162
rect 338 160 340 162
rect 20 155 22 157
rect 25 155 27 157
rect 51 155 53 157
rect 56 155 58 157
rect 61 155 63 157
rect 66 155 68 157
rect 71 155 73 157
rect 76 155 78 157
rect 81 155 83 157
rect 86 155 88 157
rect 91 155 93 157
rect 96 155 98 157
rect 101 155 103 157
rect 106 155 108 157
rect 111 155 113 157
rect 149 155 151 157
rect 154 155 156 157
rect 177 155 179 157
rect 182 155 184 157
rect 204 155 206 157
rect 209 155 211 157
rect 247 155 249 157
rect 252 155 254 157
rect 257 155 259 157
rect 262 155 264 157
rect 267 155 269 157
rect 272 155 274 157
rect 277 155 279 157
rect 282 155 284 157
rect 287 155 289 157
rect 292 155 294 157
rect 297 155 299 157
rect 302 155 304 157
rect 307 155 309 157
rect 333 155 335 157
rect 338 155 340 157
rect 5 137 7 139
rect 13 137 15 139
rect 21 137 23 139
rect 53 137 55 139
rect 61 137 63 139
rect 69 137 71 139
rect 77 137 79 139
rect 85 137 87 139
rect 93 137 95 139
rect 101 137 103 139
rect 109 137 111 139
rect 149 137 151 139
rect 154 137 156 139
rect 179 137 181 139
rect 204 137 206 139
rect 209 137 211 139
rect 249 137 251 139
rect 257 137 259 139
rect 265 137 267 139
rect 273 137 275 139
rect 281 137 283 139
rect 289 137 291 139
rect 297 137 299 139
rect 305 137 307 139
rect 337 137 339 139
rect 345 137 347 139
rect 353 137 355 139
rect 5 132 7 134
rect 13 132 15 134
rect 21 132 23 134
rect 53 132 55 134
rect 61 132 63 134
rect 69 132 71 134
rect 77 132 79 134
rect 85 132 87 134
rect 93 132 95 134
rect 101 132 103 134
rect 109 132 111 134
rect 149 132 151 134
rect 154 132 156 134
rect 179 132 181 134
rect 204 132 206 134
rect 209 132 211 134
rect 249 132 251 134
rect 257 132 259 134
rect 265 132 267 134
rect 273 132 275 134
rect 281 132 283 134
rect 289 132 291 134
rect 297 132 299 134
rect 305 132 307 134
rect 337 132 339 134
rect 345 132 347 134
rect 353 132 355 134
rect 5 120 7 122
rect 13 120 15 122
rect 21 120 23 122
rect 53 120 55 122
rect 61 120 63 122
rect 69 120 71 122
rect 77 120 79 122
rect 85 120 87 122
rect 93 120 95 122
rect 101 120 103 122
rect 109 120 111 122
rect 149 120 151 122
rect 154 120 156 122
rect 179 120 181 122
rect 204 120 206 122
rect 209 120 211 122
rect 249 120 251 122
rect 257 120 259 122
rect 265 120 267 122
rect 273 120 275 122
rect 281 120 283 122
rect 289 120 291 122
rect 297 120 299 122
rect 305 120 307 122
rect 337 120 339 122
rect 345 120 347 122
rect 353 120 355 122
rect 5 115 7 117
rect 13 115 15 117
rect 21 115 23 117
rect 53 115 55 117
rect 61 115 63 117
rect 69 115 71 117
rect 77 115 79 117
rect 85 115 87 117
rect 93 115 95 117
rect 101 115 103 117
rect 109 115 111 117
rect 149 115 151 117
rect 154 115 156 117
rect 179 115 181 117
rect 204 115 206 117
rect 209 115 211 117
rect 249 115 251 117
rect 257 115 259 117
rect 265 115 267 117
rect 273 115 275 117
rect 281 115 283 117
rect 289 115 291 117
rect 297 115 299 117
rect 305 115 307 117
rect 337 115 339 117
rect 345 115 347 117
rect 353 115 355 117
rect 18 106 20 108
rect 23 106 25 108
rect 28 106 30 108
rect 33 106 35 108
rect 38 106 40 108
rect 43 106 45 108
rect 48 106 50 108
rect 53 106 55 108
rect 58 106 60 108
rect 63 106 65 108
rect 68 106 70 108
rect 73 106 75 108
rect 78 106 80 108
rect 83 106 85 108
rect 88 106 90 108
rect 93 106 95 108
rect 98 106 100 108
rect 103 106 105 108
rect 154 106 156 108
rect 159 106 161 108
rect 164 106 166 108
rect 169 106 171 108
rect 174 106 176 108
rect 179 106 181 108
rect 184 106 186 108
rect 189 106 191 108
rect 194 106 196 108
rect 199 106 201 108
rect 204 106 206 108
rect 255 106 257 108
rect 260 106 262 108
rect 265 106 267 108
rect 270 106 272 108
rect 275 106 277 108
rect 280 106 282 108
rect 285 106 287 108
rect 290 106 292 108
rect 295 106 297 108
rect 300 106 302 108
rect 305 106 307 108
rect 310 106 312 108
rect 315 106 317 108
rect 320 106 322 108
rect 325 106 327 108
rect 330 106 332 108
rect 335 106 337 108
rect 340 106 342 108
rect 18 101 20 103
rect 23 101 25 103
rect 28 101 30 103
rect 33 101 35 103
rect 38 101 40 103
rect 43 101 45 103
rect 48 101 50 103
rect 53 101 55 103
rect 58 101 60 103
rect 63 101 65 103
rect 68 101 70 103
rect 73 101 75 103
rect 78 101 80 103
rect 83 101 85 103
rect 88 101 90 103
rect 93 101 95 103
rect 98 101 100 103
rect 103 101 105 103
rect 154 101 156 103
rect 159 101 161 103
rect 164 101 166 103
rect 169 101 171 103
rect 174 101 176 103
rect 179 101 181 103
rect 184 101 186 103
rect 189 101 191 103
rect 194 101 196 103
rect 199 101 201 103
rect 204 101 206 103
rect 255 101 257 103
rect 260 101 262 103
rect 265 101 267 103
rect 270 101 272 103
rect 275 101 277 103
rect 280 101 282 103
rect 285 101 287 103
rect 290 101 292 103
rect 295 101 297 103
rect 300 101 302 103
rect 305 101 307 103
rect 310 101 312 103
rect 315 101 317 103
rect 320 101 322 103
rect 325 101 327 103
rect 330 101 332 103
rect 335 101 337 103
rect 340 101 342 103
rect 2 74 4 76
rect 7 74 9 76
rect 24 74 26 76
rect 29 74 31 76
rect 34 74 36 76
rect 39 74 41 76
rect 319 74 321 76
rect 324 74 326 76
rect 329 74 331 76
rect 334 74 336 76
rect 351 74 353 76
rect 356 74 358 76
rect 2 69 4 71
rect 7 69 9 71
rect 24 69 26 71
rect 29 69 31 71
rect 34 69 36 71
rect 39 69 41 71
rect 319 69 321 71
rect 324 69 326 71
rect 329 69 331 71
rect 334 69 336 71
rect 351 69 353 71
rect 356 69 358 71
rect 2 64 4 66
rect 7 64 9 66
rect 24 64 26 66
rect 29 64 31 66
rect 34 64 36 66
rect 39 64 41 66
rect 319 64 321 66
rect 324 64 326 66
rect 329 64 331 66
rect 334 64 336 66
rect 351 64 353 66
rect 356 64 358 66
rect 2 59 4 61
rect 7 59 9 61
rect 24 59 26 61
rect 29 59 31 61
rect 34 59 36 61
rect 39 59 41 61
rect 319 59 321 61
rect 324 59 326 61
rect 329 59 331 61
rect 334 59 336 61
rect 351 59 353 61
rect 356 59 358 61
rect 2 54 4 56
rect 7 54 9 56
rect 24 54 26 56
rect 29 54 31 56
rect 34 54 36 56
rect 39 54 41 56
rect 319 54 321 56
rect 324 54 326 56
rect 329 54 331 56
rect 334 54 336 56
rect 351 54 353 56
rect 356 54 358 56
rect 3 7 5 9
rect 11 7 13 9
rect 21 7 23 9
rect 29 7 31 9
rect 37 7 39 9
rect 45 7 47 9
rect 53 7 55 9
rect 61 7 63 9
rect 69 7 71 9
rect 77 7 79 9
rect 85 7 87 9
rect 93 7 95 9
rect 101 7 103 9
rect 109 7 111 9
rect 117 7 119 9
rect 125 7 127 9
rect 133 7 135 9
rect 141 7 143 9
rect 149 7 151 9
rect 157 7 159 9
rect 165 7 167 9
rect 193 7 195 9
rect 201 7 203 9
rect 209 7 211 9
rect 217 7 219 9
rect 225 7 227 9
rect 233 7 235 9
rect 241 7 243 9
rect 249 7 251 9
rect 257 7 259 9
rect 265 7 267 9
rect 273 7 275 9
rect 281 7 283 9
rect 289 7 291 9
rect 297 7 299 9
rect 305 7 307 9
rect 313 7 315 9
rect 321 7 323 9
rect 329 7 331 9
rect 337 7 339 9
rect 345 7 347 9
rect 355 7 357 9
rect 3 2 5 4
rect 11 2 13 4
rect 21 2 23 4
rect 29 2 31 4
rect 37 2 39 4
rect 45 2 47 4
rect 53 2 55 4
rect 61 2 63 4
rect 69 2 71 4
rect 77 2 79 4
rect 85 2 87 4
rect 93 2 95 4
rect 101 2 103 4
rect 109 2 111 4
rect 117 2 119 4
rect 125 2 127 4
rect 133 2 135 4
rect 141 2 143 4
rect 149 2 151 4
rect 157 2 159 4
rect 165 2 167 4
rect 193 2 195 4
rect 201 2 203 4
rect 209 2 211 4
rect 217 2 219 4
rect 225 2 227 4
rect 233 2 235 4
rect 241 2 243 4
rect 249 2 251 4
rect 257 2 259 4
rect 265 2 267 4
rect 273 2 275 4
rect 281 2 283 4
rect 289 2 291 4
rect 297 2 299 4
rect 305 2 307 4
rect 313 2 315 4
rect 321 2 323 4
rect 329 2 331 4
rect 337 2 339 4
rect 345 2 347 4
rect 355 2 357 4
<< metal3 >>
rect 51 1027 309 1031
rect 51 777 55 1027
rect 305 777 309 1027
rect 51 773 309 777
rect 23 0 39 695
rect 55 0 71 695
rect 87 0 103 695
rect 119 0 135 695
rect 151 0 167 695
rect 193 0 209 695
rect 225 0 241 695
rect 257 0 273 695
rect 289 0 305 695
rect 321 0 337 695
<< gv2 >>
rect 64 1016 66 1018
rect 74 1016 76 1018
rect 84 1016 86 1018
rect 94 1016 96 1018
rect 104 1016 106 1018
rect 114 1016 116 1018
rect 124 1016 126 1018
rect 134 1016 136 1018
rect 144 1016 146 1018
rect 154 1016 156 1018
rect 164 1016 166 1018
rect 174 1016 176 1018
rect 184 1016 186 1018
rect 194 1016 196 1018
rect 204 1016 206 1018
rect 214 1016 216 1018
rect 224 1016 226 1018
rect 234 1016 236 1018
rect 244 1016 246 1018
rect 254 1016 256 1018
rect 264 1016 266 1018
rect 274 1016 276 1018
rect 284 1016 286 1018
rect 294 1016 296 1018
rect 64 1006 66 1008
rect 74 1006 76 1008
rect 84 1006 86 1008
rect 94 1006 96 1008
rect 104 1006 106 1008
rect 114 1006 116 1008
rect 124 1006 126 1008
rect 134 1006 136 1008
rect 144 1006 146 1008
rect 154 1006 156 1008
rect 164 1006 166 1008
rect 174 1006 176 1008
rect 184 1006 186 1008
rect 194 1006 196 1008
rect 204 1006 206 1008
rect 214 1006 216 1008
rect 224 1006 226 1008
rect 234 1006 236 1008
rect 244 1006 246 1008
rect 254 1006 256 1008
rect 264 1006 266 1008
rect 274 1006 276 1008
rect 284 1006 286 1008
rect 294 1006 296 1008
rect 64 996 66 998
rect 74 996 76 998
rect 84 996 86 998
rect 94 996 96 998
rect 104 996 106 998
rect 114 996 116 998
rect 124 996 126 998
rect 134 996 136 998
rect 144 996 146 998
rect 154 996 156 998
rect 164 996 166 998
rect 174 996 176 998
rect 184 996 186 998
rect 194 996 196 998
rect 204 996 206 998
rect 214 996 216 998
rect 224 996 226 998
rect 234 996 236 998
rect 244 996 246 998
rect 254 996 256 998
rect 264 996 266 998
rect 274 996 276 998
rect 284 996 286 998
rect 294 996 296 998
rect 64 986 66 988
rect 74 986 76 988
rect 84 986 86 988
rect 94 986 96 988
rect 104 986 106 988
rect 114 986 116 988
rect 124 986 126 988
rect 134 986 136 988
rect 144 986 146 988
rect 154 986 156 988
rect 164 986 166 988
rect 174 986 176 988
rect 184 986 186 988
rect 194 986 196 988
rect 204 986 206 988
rect 214 986 216 988
rect 224 986 226 988
rect 234 986 236 988
rect 244 986 246 988
rect 254 986 256 988
rect 264 986 266 988
rect 274 986 276 988
rect 284 986 286 988
rect 294 986 296 988
rect 64 976 66 978
rect 74 976 76 978
rect 84 976 86 978
rect 94 976 96 978
rect 104 976 106 978
rect 114 976 116 978
rect 124 976 126 978
rect 134 976 136 978
rect 144 976 146 978
rect 154 976 156 978
rect 164 976 166 978
rect 174 976 176 978
rect 184 976 186 978
rect 194 976 196 978
rect 204 976 206 978
rect 214 976 216 978
rect 224 976 226 978
rect 234 976 236 978
rect 244 976 246 978
rect 254 976 256 978
rect 264 976 266 978
rect 274 976 276 978
rect 284 976 286 978
rect 294 976 296 978
rect 64 966 66 968
rect 74 966 76 968
rect 84 966 86 968
rect 94 966 96 968
rect 104 966 106 968
rect 114 966 116 968
rect 124 966 126 968
rect 134 966 136 968
rect 144 966 146 968
rect 154 966 156 968
rect 164 966 166 968
rect 174 966 176 968
rect 184 966 186 968
rect 194 966 196 968
rect 204 966 206 968
rect 214 966 216 968
rect 224 966 226 968
rect 234 966 236 968
rect 244 966 246 968
rect 254 966 256 968
rect 264 966 266 968
rect 274 966 276 968
rect 284 966 286 968
rect 294 966 296 968
rect 64 956 66 958
rect 74 956 76 958
rect 84 956 86 958
rect 94 956 96 958
rect 104 956 106 958
rect 114 956 116 958
rect 124 956 126 958
rect 134 956 136 958
rect 144 956 146 958
rect 154 956 156 958
rect 164 956 166 958
rect 174 956 176 958
rect 184 956 186 958
rect 194 956 196 958
rect 204 956 206 958
rect 214 956 216 958
rect 224 956 226 958
rect 234 956 236 958
rect 244 956 246 958
rect 254 956 256 958
rect 264 956 266 958
rect 274 956 276 958
rect 284 956 286 958
rect 294 956 296 958
rect 64 946 66 948
rect 74 946 76 948
rect 84 946 86 948
rect 94 946 96 948
rect 104 946 106 948
rect 114 946 116 948
rect 124 946 126 948
rect 134 946 136 948
rect 144 946 146 948
rect 154 946 156 948
rect 164 946 166 948
rect 174 946 176 948
rect 184 946 186 948
rect 194 946 196 948
rect 204 946 206 948
rect 214 946 216 948
rect 224 946 226 948
rect 234 946 236 948
rect 244 946 246 948
rect 254 946 256 948
rect 264 946 266 948
rect 274 946 276 948
rect 284 946 286 948
rect 294 946 296 948
rect 64 936 66 938
rect 74 936 76 938
rect 84 936 86 938
rect 94 936 96 938
rect 104 936 106 938
rect 114 936 116 938
rect 124 936 126 938
rect 134 936 136 938
rect 144 936 146 938
rect 154 936 156 938
rect 164 936 166 938
rect 174 936 176 938
rect 184 936 186 938
rect 194 936 196 938
rect 204 936 206 938
rect 214 936 216 938
rect 224 936 226 938
rect 234 936 236 938
rect 244 936 246 938
rect 254 936 256 938
rect 264 936 266 938
rect 274 936 276 938
rect 284 936 286 938
rect 294 936 296 938
rect 64 926 66 928
rect 74 926 76 928
rect 84 926 86 928
rect 94 926 96 928
rect 104 926 106 928
rect 114 926 116 928
rect 124 926 126 928
rect 134 926 136 928
rect 144 926 146 928
rect 154 926 156 928
rect 164 926 166 928
rect 174 926 176 928
rect 184 926 186 928
rect 194 926 196 928
rect 204 926 206 928
rect 214 926 216 928
rect 224 926 226 928
rect 234 926 236 928
rect 244 926 246 928
rect 254 926 256 928
rect 264 926 266 928
rect 274 926 276 928
rect 284 926 286 928
rect 294 926 296 928
rect 64 916 66 918
rect 74 916 76 918
rect 84 916 86 918
rect 94 916 96 918
rect 104 916 106 918
rect 114 916 116 918
rect 124 916 126 918
rect 134 916 136 918
rect 144 916 146 918
rect 154 916 156 918
rect 164 916 166 918
rect 174 916 176 918
rect 184 916 186 918
rect 194 916 196 918
rect 204 916 206 918
rect 214 916 216 918
rect 224 916 226 918
rect 234 916 236 918
rect 244 916 246 918
rect 254 916 256 918
rect 264 916 266 918
rect 274 916 276 918
rect 284 916 286 918
rect 294 916 296 918
rect 64 906 66 908
rect 74 906 76 908
rect 84 906 86 908
rect 94 906 96 908
rect 104 906 106 908
rect 114 906 116 908
rect 124 906 126 908
rect 134 906 136 908
rect 144 906 146 908
rect 154 906 156 908
rect 164 906 166 908
rect 174 906 176 908
rect 184 906 186 908
rect 194 906 196 908
rect 204 906 206 908
rect 214 906 216 908
rect 224 906 226 908
rect 234 906 236 908
rect 244 906 246 908
rect 254 906 256 908
rect 264 906 266 908
rect 274 906 276 908
rect 284 906 286 908
rect 294 906 296 908
rect 64 896 66 898
rect 74 896 76 898
rect 84 896 86 898
rect 94 896 96 898
rect 104 896 106 898
rect 114 896 116 898
rect 124 896 126 898
rect 134 896 136 898
rect 144 896 146 898
rect 154 896 156 898
rect 164 896 166 898
rect 174 896 176 898
rect 184 896 186 898
rect 194 896 196 898
rect 204 896 206 898
rect 214 896 216 898
rect 224 896 226 898
rect 234 896 236 898
rect 244 896 246 898
rect 254 896 256 898
rect 264 896 266 898
rect 274 896 276 898
rect 284 896 286 898
rect 294 896 296 898
rect 64 886 66 888
rect 74 886 76 888
rect 84 886 86 888
rect 94 886 96 888
rect 104 886 106 888
rect 114 886 116 888
rect 124 886 126 888
rect 134 886 136 888
rect 144 886 146 888
rect 154 886 156 888
rect 164 886 166 888
rect 174 886 176 888
rect 184 886 186 888
rect 194 886 196 888
rect 204 886 206 888
rect 214 886 216 888
rect 224 886 226 888
rect 234 886 236 888
rect 244 886 246 888
rect 254 886 256 888
rect 264 886 266 888
rect 274 886 276 888
rect 284 886 286 888
rect 294 886 296 888
rect 64 876 66 878
rect 74 876 76 878
rect 84 876 86 878
rect 94 876 96 878
rect 104 876 106 878
rect 114 876 116 878
rect 124 876 126 878
rect 134 876 136 878
rect 144 876 146 878
rect 154 876 156 878
rect 164 876 166 878
rect 174 876 176 878
rect 184 876 186 878
rect 194 876 196 878
rect 204 876 206 878
rect 214 876 216 878
rect 224 876 226 878
rect 234 876 236 878
rect 244 876 246 878
rect 254 876 256 878
rect 264 876 266 878
rect 274 876 276 878
rect 284 876 286 878
rect 294 876 296 878
rect 64 866 66 868
rect 74 866 76 868
rect 84 866 86 868
rect 94 866 96 868
rect 104 866 106 868
rect 114 866 116 868
rect 124 866 126 868
rect 134 866 136 868
rect 144 866 146 868
rect 154 866 156 868
rect 164 866 166 868
rect 174 866 176 868
rect 184 866 186 868
rect 194 866 196 868
rect 204 866 206 868
rect 214 866 216 868
rect 224 866 226 868
rect 234 866 236 868
rect 244 866 246 868
rect 254 866 256 868
rect 264 866 266 868
rect 274 866 276 868
rect 284 866 286 868
rect 294 866 296 868
rect 64 856 66 858
rect 74 856 76 858
rect 84 856 86 858
rect 94 856 96 858
rect 104 856 106 858
rect 114 856 116 858
rect 124 856 126 858
rect 134 856 136 858
rect 144 856 146 858
rect 154 856 156 858
rect 164 856 166 858
rect 174 856 176 858
rect 184 856 186 858
rect 194 856 196 858
rect 204 856 206 858
rect 214 856 216 858
rect 224 856 226 858
rect 234 856 236 858
rect 244 856 246 858
rect 254 856 256 858
rect 264 856 266 858
rect 274 856 276 858
rect 284 856 286 858
rect 294 856 296 858
rect 64 846 66 848
rect 74 846 76 848
rect 84 846 86 848
rect 94 846 96 848
rect 104 846 106 848
rect 114 846 116 848
rect 124 846 126 848
rect 134 846 136 848
rect 144 846 146 848
rect 154 846 156 848
rect 164 846 166 848
rect 174 846 176 848
rect 184 846 186 848
rect 194 846 196 848
rect 204 846 206 848
rect 214 846 216 848
rect 224 846 226 848
rect 234 846 236 848
rect 244 846 246 848
rect 254 846 256 848
rect 264 846 266 848
rect 274 846 276 848
rect 284 846 286 848
rect 294 846 296 848
rect 64 836 66 838
rect 74 836 76 838
rect 84 836 86 838
rect 94 836 96 838
rect 104 836 106 838
rect 114 836 116 838
rect 124 836 126 838
rect 134 836 136 838
rect 144 836 146 838
rect 154 836 156 838
rect 164 836 166 838
rect 174 836 176 838
rect 184 836 186 838
rect 194 836 196 838
rect 204 836 206 838
rect 214 836 216 838
rect 224 836 226 838
rect 234 836 236 838
rect 244 836 246 838
rect 254 836 256 838
rect 264 836 266 838
rect 274 836 276 838
rect 284 836 286 838
rect 294 836 296 838
rect 64 826 66 828
rect 74 826 76 828
rect 84 826 86 828
rect 94 826 96 828
rect 104 826 106 828
rect 114 826 116 828
rect 124 826 126 828
rect 134 826 136 828
rect 144 826 146 828
rect 154 826 156 828
rect 164 826 166 828
rect 174 826 176 828
rect 184 826 186 828
rect 194 826 196 828
rect 204 826 206 828
rect 214 826 216 828
rect 224 826 226 828
rect 234 826 236 828
rect 244 826 246 828
rect 254 826 256 828
rect 264 826 266 828
rect 274 826 276 828
rect 284 826 286 828
rect 294 826 296 828
rect 64 816 66 818
rect 74 816 76 818
rect 84 816 86 818
rect 94 816 96 818
rect 104 816 106 818
rect 114 816 116 818
rect 124 816 126 818
rect 134 816 136 818
rect 144 816 146 818
rect 154 816 156 818
rect 164 816 166 818
rect 174 816 176 818
rect 184 816 186 818
rect 194 816 196 818
rect 204 816 206 818
rect 214 816 216 818
rect 224 816 226 818
rect 234 816 236 818
rect 244 816 246 818
rect 254 816 256 818
rect 264 816 266 818
rect 274 816 276 818
rect 284 816 286 818
rect 294 816 296 818
rect 64 806 66 808
rect 74 806 76 808
rect 84 806 86 808
rect 94 806 96 808
rect 104 806 106 808
rect 114 806 116 808
rect 124 806 126 808
rect 134 806 136 808
rect 144 806 146 808
rect 154 806 156 808
rect 164 806 166 808
rect 174 806 176 808
rect 184 806 186 808
rect 194 806 196 808
rect 204 806 206 808
rect 214 806 216 808
rect 224 806 226 808
rect 234 806 236 808
rect 244 806 246 808
rect 254 806 256 808
rect 264 806 266 808
rect 274 806 276 808
rect 284 806 286 808
rect 294 806 296 808
rect 64 796 66 798
rect 74 796 76 798
rect 84 796 86 798
rect 94 796 96 798
rect 104 796 106 798
rect 114 796 116 798
rect 124 796 126 798
rect 134 796 136 798
rect 144 796 146 798
rect 154 796 156 798
rect 164 796 166 798
rect 174 796 176 798
rect 184 796 186 798
rect 194 796 196 798
rect 204 796 206 798
rect 214 796 216 798
rect 224 796 226 798
rect 234 796 236 798
rect 244 796 246 798
rect 254 796 256 798
rect 264 796 266 798
rect 274 796 276 798
rect 284 796 286 798
rect 294 796 296 798
rect 64 786 66 788
rect 74 786 76 788
rect 84 786 86 788
rect 94 786 96 788
rect 104 786 106 788
rect 114 786 116 788
rect 124 786 126 788
rect 134 786 136 788
rect 144 786 146 788
rect 154 786 156 788
rect 164 786 166 788
rect 174 786 176 788
rect 184 786 186 788
rect 194 786 196 788
rect 204 786 206 788
rect 214 786 216 788
rect 224 786 226 788
rect 234 786 236 788
rect 244 786 246 788
rect 254 786 256 788
rect 264 786 266 788
rect 274 786 276 788
rect 284 786 286 788
rect 294 786 296 788
rect 25 691 27 693
rect 30 691 32 693
rect 35 691 37 693
rect 89 691 91 693
rect 94 691 96 693
rect 99 691 101 693
rect 153 691 155 693
rect 158 691 160 693
rect 163 691 165 693
rect 227 691 229 693
rect 232 691 234 693
rect 237 691 239 693
rect 291 691 293 693
rect 296 691 298 693
rect 301 691 303 693
rect 25 686 27 688
rect 30 686 32 688
rect 35 686 37 688
rect 89 686 91 688
rect 94 686 96 688
rect 99 686 101 688
rect 153 686 155 688
rect 158 686 160 688
rect 163 686 165 688
rect 227 686 229 688
rect 232 686 234 688
rect 237 686 239 688
rect 291 686 293 688
rect 296 686 298 688
rect 301 686 303 688
rect 57 668 59 670
rect 62 668 64 670
rect 67 668 69 670
rect 121 668 123 670
rect 126 668 128 670
rect 131 668 133 670
rect 195 668 197 670
rect 200 668 202 670
rect 205 668 207 670
rect 259 668 261 670
rect 264 668 266 670
rect 269 668 271 670
rect 323 668 325 670
rect 328 668 330 670
rect 333 668 335 670
rect 57 663 59 665
rect 62 663 64 665
rect 67 663 69 665
rect 121 663 123 665
rect 126 663 128 665
rect 131 663 133 665
rect 195 663 197 665
rect 200 663 202 665
rect 205 663 207 665
rect 259 663 261 665
rect 264 663 266 665
rect 269 663 271 665
rect 323 663 325 665
rect 328 663 330 665
rect 333 663 335 665
rect 57 658 59 660
rect 62 658 64 660
rect 67 658 69 660
rect 121 658 123 660
rect 126 658 128 660
rect 131 658 133 660
rect 195 658 197 660
rect 200 658 202 660
rect 205 658 207 660
rect 259 658 261 660
rect 264 658 266 660
rect 269 658 271 660
rect 323 658 325 660
rect 328 658 330 660
rect 333 658 335 660
rect 25 640 27 642
rect 30 640 32 642
rect 35 640 37 642
rect 89 640 91 642
rect 94 640 96 642
rect 99 640 101 642
rect 153 640 155 642
rect 158 640 160 642
rect 163 640 165 642
rect 227 640 229 642
rect 232 640 234 642
rect 237 640 239 642
rect 291 640 293 642
rect 296 640 298 642
rect 301 640 303 642
rect 25 635 27 637
rect 30 635 32 637
rect 35 635 37 637
rect 89 635 91 637
rect 94 635 96 637
rect 99 635 101 637
rect 153 635 155 637
rect 158 635 160 637
rect 163 635 165 637
rect 227 635 229 637
rect 232 635 234 637
rect 237 635 239 637
rect 291 635 293 637
rect 296 635 298 637
rect 301 635 303 637
rect 25 630 27 632
rect 30 630 32 632
rect 35 630 37 632
rect 89 630 91 632
rect 94 630 96 632
rect 99 630 101 632
rect 153 630 155 632
rect 158 630 160 632
rect 163 630 165 632
rect 227 630 229 632
rect 232 630 234 632
rect 237 630 239 632
rect 291 630 293 632
rect 296 630 298 632
rect 301 630 303 632
rect 25 625 27 627
rect 30 625 32 627
rect 35 625 37 627
rect 89 625 91 627
rect 94 625 96 627
rect 99 625 101 627
rect 153 625 155 627
rect 158 625 160 627
rect 163 625 165 627
rect 227 625 229 627
rect 232 625 234 627
rect 237 625 239 627
rect 291 625 293 627
rect 296 625 298 627
rect 301 625 303 627
rect 25 620 27 622
rect 30 620 32 622
rect 35 620 37 622
rect 89 620 91 622
rect 94 620 96 622
rect 99 620 101 622
rect 153 620 155 622
rect 158 620 160 622
rect 163 620 165 622
rect 227 620 229 622
rect 232 620 234 622
rect 237 620 239 622
rect 291 620 293 622
rect 296 620 298 622
rect 301 620 303 622
rect 57 603 59 605
rect 62 603 64 605
rect 67 603 69 605
rect 121 603 123 605
rect 126 603 128 605
rect 131 603 133 605
rect 195 603 197 605
rect 200 603 202 605
rect 205 603 207 605
rect 259 603 261 605
rect 264 603 266 605
rect 269 603 271 605
rect 323 603 325 605
rect 328 603 330 605
rect 333 603 335 605
rect 57 598 59 600
rect 62 598 64 600
rect 67 598 69 600
rect 121 598 123 600
rect 126 598 128 600
rect 131 598 133 600
rect 195 598 197 600
rect 200 598 202 600
rect 205 598 207 600
rect 259 598 261 600
rect 264 598 266 600
rect 269 598 271 600
rect 323 598 325 600
rect 328 598 330 600
rect 333 598 335 600
rect 57 593 59 595
rect 62 593 64 595
rect 67 593 69 595
rect 121 593 123 595
rect 126 593 128 595
rect 131 593 133 595
rect 195 593 197 595
rect 200 593 202 595
rect 205 593 207 595
rect 259 593 261 595
rect 264 593 266 595
rect 269 593 271 595
rect 323 593 325 595
rect 328 593 330 595
rect 333 593 335 595
rect 25 580 27 582
rect 30 580 32 582
rect 35 580 37 582
rect 89 580 91 582
rect 94 580 96 582
rect 99 580 101 582
rect 153 580 155 582
rect 158 580 160 582
rect 163 580 165 582
rect 227 580 229 582
rect 232 580 234 582
rect 237 580 239 582
rect 291 580 293 582
rect 296 580 298 582
rect 301 580 303 582
rect 25 575 27 577
rect 30 575 32 577
rect 35 575 37 577
rect 89 575 91 577
rect 94 575 96 577
rect 99 575 101 577
rect 153 575 155 577
rect 158 575 160 577
rect 163 575 165 577
rect 227 575 229 577
rect 232 575 234 577
rect 237 575 239 577
rect 291 575 293 577
rect 296 575 298 577
rect 301 575 303 577
rect 25 570 27 572
rect 30 570 32 572
rect 35 570 37 572
rect 89 570 91 572
rect 94 570 96 572
rect 99 570 101 572
rect 153 570 155 572
rect 158 570 160 572
rect 163 570 165 572
rect 227 570 229 572
rect 232 570 234 572
rect 237 570 239 572
rect 291 570 293 572
rect 296 570 298 572
rect 301 570 303 572
rect 25 565 27 567
rect 30 565 32 567
rect 35 565 37 567
rect 89 565 91 567
rect 94 565 96 567
rect 99 565 101 567
rect 153 565 155 567
rect 158 565 160 567
rect 163 565 165 567
rect 227 565 229 567
rect 232 565 234 567
rect 237 565 239 567
rect 291 565 293 567
rect 296 565 298 567
rect 301 565 303 567
rect 25 560 27 562
rect 30 560 32 562
rect 35 560 37 562
rect 89 560 91 562
rect 94 560 96 562
rect 99 560 101 562
rect 153 560 155 562
rect 158 560 160 562
rect 163 560 165 562
rect 227 560 229 562
rect 232 560 234 562
rect 237 560 239 562
rect 291 560 293 562
rect 296 560 298 562
rect 301 560 303 562
rect 57 538 59 540
rect 62 538 64 540
rect 67 538 69 540
rect 121 538 123 540
rect 126 538 128 540
rect 131 538 133 540
rect 195 537 197 539
rect 200 537 202 539
rect 205 537 207 539
rect 259 538 261 540
rect 264 538 266 540
rect 269 538 271 540
rect 323 538 325 540
rect 328 538 330 540
rect 333 538 335 540
rect 57 533 59 535
rect 62 533 64 535
rect 67 533 69 535
rect 121 533 123 535
rect 126 533 128 535
rect 131 533 133 535
rect 195 532 197 534
rect 200 532 202 534
rect 205 532 207 534
rect 259 533 261 535
rect 264 533 266 535
rect 269 533 271 535
rect 323 533 325 535
rect 328 533 330 535
rect 333 533 335 535
rect 57 528 59 530
rect 62 528 64 530
rect 67 528 69 530
rect 121 528 123 530
rect 126 528 128 530
rect 131 528 133 530
rect 195 527 197 529
rect 200 527 202 529
rect 205 527 207 529
rect 259 528 261 530
rect 264 528 266 530
rect 269 528 271 530
rect 323 528 325 530
rect 328 528 330 530
rect 333 528 335 530
rect 25 515 27 517
rect 30 515 32 517
rect 35 515 37 517
rect 89 515 91 517
rect 94 515 96 517
rect 99 515 101 517
rect 153 515 155 517
rect 158 515 160 517
rect 163 515 165 517
rect 227 515 229 517
rect 232 515 234 517
rect 237 515 239 517
rect 291 515 293 517
rect 296 515 298 517
rect 301 515 303 517
rect 25 510 27 512
rect 30 510 32 512
rect 35 510 37 512
rect 89 510 91 512
rect 94 510 96 512
rect 99 510 101 512
rect 153 510 155 512
rect 158 510 160 512
rect 163 510 165 512
rect 227 510 229 512
rect 232 510 234 512
rect 237 510 239 512
rect 291 510 293 512
rect 296 510 298 512
rect 301 510 303 512
rect 25 505 27 507
rect 30 505 32 507
rect 35 505 37 507
rect 89 505 91 507
rect 94 505 96 507
rect 99 505 101 507
rect 153 505 155 507
rect 158 505 160 507
rect 163 505 165 507
rect 227 505 229 507
rect 232 505 234 507
rect 237 505 239 507
rect 291 505 293 507
rect 296 505 298 507
rect 301 505 303 507
rect 25 500 27 502
rect 30 500 32 502
rect 35 500 37 502
rect 89 500 91 502
rect 94 500 96 502
rect 99 500 101 502
rect 153 500 155 502
rect 158 500 160 502
rect 163 500 165 502
rect 227 500 229 502
rect 232 500 234 502
rect 237 500 239 502
rect 291 500 293 502
rect 296 500 298 502
rect 301 500 303 502
rect 25 495 27 497
rect 30 495 32 497
rect 35 495 37 497
rect 89 495 91 497
rect 94 495 96 497
rect 99 495 101 497
rect 153 495 155 497
rect 158 495 160 497
rect 163 495 165 497
rect 227 495 229 497
rect 232 495 234 497
rect 237 495 239 497
rect 291 495 293 497
rect 296 495 298 497
rect 301 495 303 497
rect 57 473 59 475
rect 62 473 64 475
rect 67 473 69 475
rect 121 473 123 475
rect 126 473 128 475
rect 131 473 133 475
rect 195 472 197 474
rect 200 472 202 474
rect 205 472 207 474
rect 259 473 261 475
rect 264 473 266 475
rect 269 473 271 475
rect 323 473 325 475
rect 328 473 330 475
rect 333 473 335 475
rect 57 468 59 470
rect 62 468 64 470
rect 67 468 69 470
rect 121 468 123 470
rect 126 468 128 470
rect 131 468 133 470
rect 195 467 197 469
rect 200 467 202 469
rect 205 467 207 469
rect 259 468 261 470
rect 264 468 266 470
rect 269 468 271 470
rect 323 468 325 470
rect 328 468 330 470
rect 333 468 335 470
rect 57 463 59 465
rect 62 463 64 465
rect 67 463 69 465
rect 121 463 123 465
rect 126 463 128 465
rect 131 463 133 465
rect 195 462 197 464
rect 200 462 202 464
rect 205 462 207 464
rect 259 463 261 465
rect 264 463 266 465
rect 269 463 271 465
rect 323 463 325 465
rect 328 463 330 465
rect 333 463 335 465
rect 25 445 27 447
rect 30 445 32 447
rect 35 445 37 447
rect 89 445 91 447
rect 94 445 96 447
rect 99 445 101 447
rect 153 445 155 447
rect 158 445 160 447
rect 163 445 165 447
rect 227 445 229 447
rect 232 445 234 447
rect 237 445 239 447
rect 291 445 293 447
rect 296 445 298 447
rect 301 445 303 447
rect 25 440 27 442
rect 30 440 32 442
rect 35 440 37 442
rect 89 440 91 442
rect 94 440 96 442
rect 99 440 101 442
rect 153 440 155 442
rect 158 440 160 442
rect 163 440 165 442
rect 227 440 229 442
rect 232 440 234 442
rect 237 440 239 442
rect 291 440 293 442
rect 296 440 298 442
rect 301 440 303 442
rect 57 428 59 430
rect 62 428 64 430
rect 67 428 69 430
rect 121 428 123 430
rect 126 428 128 430
rect 131 428 133 430
rect 195 428 197 430
rect 200 428 202 430
rect 205 428 207 430
rect 259 428 261 430
rect 264 428 266 430
rect 269 428 271 430
rect 323 428 325 430
rect 328 428 330 430
rect 333 428 335 430
rect 57 423 59 425
rect 62 423 64 425
rect 67 423 69 425
rect 121 423 123 425
rect 126 423 128 425
rect 131 423 133 425
rect 195 423 197 425
rect 200 423 202 425
rect 205 423 207 425
rect 259 423 261 425
rect 264 423 266 425
rect 269 423 271 425
rect 323 423 325 425
rect 328 423 330 425
rect 333 423 335 425
rect 25 400 27 402
rect 30 400 32 402
rect 35 400 37 402
rect 89 400 91 402
rect 94 400 96 402
rect 99 400 101 402
rect 153 400 155 402
rect 158 400 160 402
rect 163 400 165 402
rect 227 400 229 402
rect 232 400 234 402
rect 237 400 239 402
rect 291 400 293 402
rect 296 400 298 402
rect 301 400 303 402
rect 25 395 27 397
rect 30 395 32 397
rect 35 395 37 397
rect 89 395 91 397
rect 94 395 96 397
rect 99 395 101 397
rect 153 395 155 397
rect 158 395 160 397
rect 163 395 165 397
rect 227 395 229 397
rect 232 395 234 397
rect 237 395 239 397
rect 291 395 293 397
rect 296 395 298 397
rect 301 395 303 397
rect 57 383 59 385
rect 62 383 64 385
rect 67 383 69 385
rect 121 383 123 385
rect 126 383 128 385
rect 131 383 133 385
rect 195 383 197 385
rect 200 383 202 385
rect 205 383 207 385
rect 259 383 261 385
rect 264 383 266 385
rect 269 383 271 385
rect 323 383 325 385
rect 328 383 330 385
rect 333 383 335 385
rect 57 378 59 380
rect 62 378 64 380
rect 67 378 69 380
rect 121 378 123 380
rect 126 378 128 380
rect 131 378 133 380
rect 195 378 197 380
rect 200 378 202 380
rect 205 378 207 380
rect 259 378 261 380
rect 264 378 266 380
rect 269 378 271 380
rect 323 378 325 380
rect 328 378 330 380
rect 333 378 335 380
rect 25 360 27 362
rect 30 360 32 362
rect 35 360 37 362
rect 89 360 91 362
rect 94 360 96 362
rect 99 360 101 362
rect 153 360 155 362
rect 158 360 160 362
rect 163 360 165 362
rect 227 360 229 362
rect 232 360 234 362
rect 237 360 239 362
rect 291 360 293 362
rect 296 360 298 362
rect 301 360 303 362
rect 25 355 27 357
rect 30 355 32 357
rect 35 355 37 357
rect 89 355 91 357
rect 94 355 96 357
rect 99 355 101 357
rect 153 355 155 357
rect 158 355 160 357
rect 163 355 165 357
rect 227 355 229 357
rect 232 355 234 357
rect 237 355 239 357
rect 291 355 293 357
rect 296 355 298 357
rect 301 355 303 357
rect 25 350 27 352
rect 30 350 32 352
rect 35 350 37 352
rect 89 350 91 352
rect 94 350 96 352
rect 99 350 101 352
rect 153 350 155 352
rect 158 350 160 352
rect 163 350 165 352
rect 227 350 229 352
rect 232 350 234 352
rect 237 350 239 352
rect 291 350 293 352
rect 296 350 298 352
rect 301 350 303 352
rect 57 332 59 334
rect 62 332 64 334
rect 67 332 69 334
rect 121 332 123 334
rect 126 332 128 334
rect 131 332 133 334
rect 195 332 197 334
rect 200 332 202 334
rect 205 332 207 334
rect 259 332 261 334
rect 264 332 266 334
rect 269 332 271 334
rect 323 332 325 334
rect 328 332 330 334
rect 333 332 335 334
rect 57 327 59 329
rect 62 327 64 329
rect 67 327 69 329
rect 121 327 123 329
rect 126 327 128 329
rect 131 327 133 329
rect 195 327 197 329
rect 200 327 202 329
rect 205 327 207 329
rect 259 327 261 329
rect 264 327 266 329
rect 269 327 271 329
rect 323 327 325 329
rect 328 327 330 329
rect 333 327 335 329
rect 57 322 59 324
rect 62 322 64 324
rect 67 322 69 324
rect 121 322 123 324
rect 126 322 128 324
rect 131 322 133 324
rect 195 322 197 324
rect 200 322 202 324
rect 205 322 207 324
rect 259 322 261 324
rect 264 322 266 324
rect 269 322 271 324
rect 323 322 325 324
rect 328 322 330 324
rect 333 322 335 324
rect 57 317 59 319
rect 62 317 64 319
rect 67 317 69 319
rect 121 317 123 319
rect 126 317 128 319
rect 131 317 133 319
rect 195 317 197 319
rect 200 317 202 319
rect 205 317 207 319
rect 259 317 261 319
rect 264 317 266 319
rect 269 317 271 319
rect 323 317 325 319
rect 328 317 330 319
rect 333 317 335 319
rect 57 312 59 314
rect 62 312 64 314
rect 67 312 69 314
rect 121 312 123 314
rect 126 312 128 314
rect 131 312 133 314
rect 195 312 197 314
rect 200 312 202 314
rect 205 312 207 314
rect 259 312 261 314
rect 264 312 266 314
rect 269 312 271 314
rect 323 312 325 314
rect 328 312 330 314
rect 333 312 335 314
rect 25 295 27 297
rect 30 295 32 297
rect 35 295 37 297
rect 89 295 91 297
rect 94 295 96 297
rect 99 295 101 297
rect 153 295 155 297
rect 158 295 160 297
rect 163 295 165 297
rect 227 295 229 297
rect 232 295 234 297
rect 237 295 239 297
rect 291 295 293 297
rect 296 295 298 297
rect 301 295 303 297
rect 25 290 27 292
rect 30 290 32 292
rect 35 290 37 292
rect 89 290 91 292
rect 94 290 96 292
rect 99 290 101 292
rect 153 290 155 292
rect 158 290 160 292
rect 163 290 165 292
rect 227 290 229 292
rect 232 290 234 292
rect 237 290 239 292
rect 291 290 293 292
rect 296 290 298 292
rect 301 290 303 292
rect 25 285 27 287
rect 30 285 32 287
rect 35 285 37 287
rect 89 285 91 287
rect 94 285 96 287
rect 99 285 101 287
rect 153 285 155 287
rect 158 285 160 287
rect 163 285 165 287
rect 227 285 229 287
rect 232 285 234 287
rect 237 285 239 287
rect 291 285 293 287
rect 296 285 298 287
rect 301 285 303 287
rect 57 272 59 274
rect 62 272 64 274
rect 67 272 69 274
rect 121 272 123 274
rect 126 272 128 274
rect 131 272 133 274
rect 195 272 197 274
rect 200 272 202 274
rect 205 272 207 274
rect 259 272 261 274
rect 264 272 266 274
rect 269 272 271 274
rect 323 272 325 274
rect 328 272 330 274
rect 333 272 335 274
rect 57 267 59 269
rect 62 267 64 269
rect 67 267 69 269
rect 121 267 123 269
rect 126 267 128 269
rect 131 267 133 269
rect 195 267 197 269
rect 200 267 202 269
rect 205 267 207 269
rect 259 267 261 269
rect 264 267 266 269
rect 269 267 271 269
rect 323 267 325 269
rect 328 267 330 269
rect 333 267 335 269
rect 57 262 59 264
rect 62 262 64 264
rect 67 262 69 264
rect 121 262 123 264
rect 126 262 128 264
rect 131 262 133 264
rect 195 262 197 264
rect 200 262 202 264
rect 205 262 207 264
rect 259 262 261 264
rect 264 262 266 264
rect 269 262 271 264
rect 323 262 325 264
rect 328 262 330 264
rect 333 262 335 264
rect 57 257 59 259
rect 62 257 64 259
rect 67 257 69 259
rect 121 257 123 259
rect 126 257 128 259
rect 131 257 133 259
rect 195 257 197 259
rect 200 257 202 259
rect 205 257 207 259
rect 259 257 261 259
rect 264 257 266 259
rect 269 257 271 259
rect 323 257 325 259
rect 328 257 330 259
rect 333 257 335 259
rect 57 252 59 254
rect 62 252 64 254
rect 67 252 69 254
rect 121 252 123 254
rect 126 252 128 254
rect 131 252 133 254
rect 195 252 197 254
rect 200 252 202 254
rect 205 252 207 254
rect 259 252 261 254
rect 264 252 266 254
rect 269 252 271 254
rect 323 252 325 254
rect 328 252 330 254
rect 333 252 335 254
rect 25 230 27 232
rect 30 230 32 232
rect 35 230 37 232
rect 89 230 91 232
rect 94 230 96 232
rect 99 230 101 232
rect 153 230 155 232
rect 158 230 160 232
rect 163 230 165 232
rect 227 230 229 232
rect 232 230 234 232
rect 237 230 239 232
rect 291 230 293 232
rect 296 230 298 232
rect 301 230 303 232
rect 25 225 27 227
rect 30 225 32 227
rect 35 225 37 227
rect 89 225 91 227
rect 94 225 96 227
rect 99 225 101 227
rect 153 225 155 227
rect 158 225 160 227
rect 163 225 165 227
rect 227 225 229 227
rect 232 225 234 227
rect 237 225 239 227
rect 291 225 293 227
rect 296 225 298 227
rect 301 225 303 227
rect 25 220 27 222
rect 30 220 32 222
rect 35 220 37 222
rect 89 220 91 222
rect 94 220 96 222
rect 99 220 101 222
rect 153 220 155 222
rect 158 220 160 222
rect 163 220 165 222
rect 227 220 229 222
rect 232 220 234 222
rect 237 220 239 222
rect 291 220 293 222
rect 296 220 298 222
rect 301 220 303 222
rect 57 207 59 209
rect 62 207 64 209
rect 67 207 69 209
rect 121 207 123 209
rect 126 207 128 209
rect 131 207 133 209
rect 195 207 197 209
rect 200 207 202 209
rect 205 207 207 209
rect 259 207 261 209
rect 264 207 266 209
rect 269 207 271 209
rect 323 207 325 209
rect 328 207 330 209
rect 333 207 335 209
rect 57 202 59 204
rect 62 202 64 204
rect 67 202 69 204
rect 121 202 123 204
rect 126 202 128 204
rect 131 202 133 204
rect 195 202 197 204
rect 200 202 202 204
rect 205 202 207 204
rect 259 202 261 204
rect 264 202 266 204
rect 269 202 271 204
rect 323 202 325 204
rect 328 202 330 204
rect 333 202 335 204
rect 57 197 59 199
rect 62 197 64 199
rect 67 197 69 199
rect 121 197 123 199
rect 126 197 128 199
rect 131 197 133 199
rect 195 197 197 199
rect 200 197 202 199
rect 205 197 207 199
rect 259 197 261 199
rect 264 197 266 199
rect 269 197 271 199
rect 323 197 325 199
rect 328 197 330 199
rect 333 197 335 199
rect 57 192 59 194
rect 62 192 64 194
rect 67 192 69 194
rect 121 192 123 194
rect 126 192 128 194
rect 131 192 133 194
rect 195 192 197 194
rect 200 192 202 194
rect 205 192 207 194
rect 259 192 261 194
rect 264 192 266 194
rect 269 192 271 194
rect 323 192 325 194
rect 328 192 330 194
rect 333 192 335 194
rect 57 187 59 189
rect 62 187 64 189
rect 67 187 69 189
rect 121 187 123 189
rect 126 187 128 189
rect 131 187 133 189
rect 195 187 197 189
rect 200 187 202 189
rect 205 187 207 189
rect 259 187 261 189
rect 264 187 266 189
rect 269 187 271 189
rect 323 187 325 189
rect 328 187 330 189
rect 333 187 335 189
rect 25 165 27 167
rect 30 165 32 167
rect 35 165 37 167
rect 89 165 91 167
rect 94 165 96 167
rect 99 165 101 167
rect 153 165 155 167
rect 158 165 160 167
rect 163 165 165 167
rect 227 165 229 167
rect 232 165 234 167
rect 237 165 239 167
rect 291 165 293 167
rect 296 165 298 167
rect 301 165 303 167
rect 25 160 27 162
rect 30 160 32 162
rect 35 160 37 162
rect 89 160 91 162
rect 94 160 96 162
rect 99 160 101 162
rect 153 160 155 162
rect 158 160 160 162
rect 163 160 165 162
rect 227 160 229 162
rect 232 160 234 162
rect 237 160 239 162
rect 291 160 293 162
rect 296 160 298 162
rect 301 160 303 162
rect 25 155 27 157
rect 30 155 32 157
rect 35 155 37 157
rect 89 155 91 157
rect 94 155 96 157
rect 99 155 101 157
rect 153 155 155 157
rect 158 155 160 157
rect 163 155 165 157
rect 227 155 229 157
rect 232 155 234 157
rect 237 155 239 157
rect 291 155 293 157
rect 296 155 298 157
rect 301 155 303 157
rect 57 137 59 139
rect 62 137 64 139
rect 67 137 69 139
rect 121 137 123 139
rect 126 137 128 139
rect 131 137 133 139
rect 195 137 197 139
rect 200 137 202 139
rect 205 137 207 139
rect 259 137 261 139
rect 264 137 266 139
rect 269 137 271 139
rect 323 137 325 139
rect 328 137 330 139
rect 333 137 335 139
rect 57 132 59 134
rect 62 132 64 134
rect 67 132 69 134
rect 121 132 123 134
rect 126 132 128 134
rect 131 132 133 134
rect 195 132 197 134
rect 200 132 202 134
rect 205 132 207 134
rect 259 132 261 134
rect 264 132 266 134
rect 269 132 271 134
rect 323 132 325 134
rect 328 132 330 134
rect 333 132 335 134
rect 25 120 27 122
rect 30 120 32 122
rect 35 120 37 122
rect 89 120 91 122
rect 94 120 96 122
rect 99 120 101 122
rect 153 120 155 122
rect 158 120 160 122
rect 163 120 165 122
rect 227 120 229 122
rect 232 120 234 122
rect 237 120 239 122
rect 291 120 293 122
rect 296 120 298 122
rect 301 120 303 122
rect 25 115 27 117
rect 30 115 32 117
rect 35 115 37 117
rect 89 115 91 117
rect 94 115 96 117
rect 99 115 101 117
rect 153 115 155 117
rect 158 115 160 117
rect 163 115 165 117
rect 227 115 229 117
rect 232 115 234 117
rect 237 115 239 117
rect 291 115 293 117
rect 296 115 298 117
rect 301 115 303 117
rect 25 74 27 76
rect 30 74 32 76
rect 35 74 37 76
rect 291 74 293 76
rect 296 74 298 76
rect 301 74 303 76
rect 25 69 27 71
rect 30 69 32 71
rect 35 69 37 71
rect 291 69 293 71
rect 296 69 298 71
rect 301 69 303 71
rect 25 64 27 66
rect 30 64 32 66
rect 35 64 37 66
rect 291 64 293 66
rect 296 64 298 66
rect 301 64 303 66
rect 25 59 27 61
rect 30 59 32 61
rect 35 59 37 61
rect 291 59 293 61
rect 296 59 298 61
rect 301 59 303 61
rect 25 54 27 56
rect 30 54 32 56
rect 35 54 37 56
rect 291 54 293 56
rect 296 54 298 56
rect 301 54 303 56
rect 25 7 27 9
rect 30 7 32 9
rect 35 7 37 9
rect 89 7 91 9
rect 94 7 96 9
rect 99 7 101 9
rect 153 7 155 9
rect 158 7 160 9
rect 163 7 165 9
rect 227 7 229 9
rect 232 7 234 9
rect 237 7 239 9
rect 291 7 293 9
rect 296 7 298 9
rect 301 7 303 9
rect 25 2 27 4
rect 30 2 32 4
rect 35 2 37 4
rect 89 2 91 4
rect 94 2 96 4
rect 99 2 101 4
rect 153 2 155 4
rect 158 2 160 4
rect 163 2 165 4
rect 227 2 229 4
rect 232 2 234 4
rect 237 2 239 4
rect 291 2 293 4
rect 296 2 298 4
rect 301 2 303 4
<< pad >>
rect 55 777 305 1027
<< pseudo_rnwell >>
rect 80 47 81 71
rect 279 47 280 71
<< rnwell >>
rect 81 47 279 71
<< labels >>
rlabel rnwell s 168 57 168 57 2 r0_body
rlabel metal1 s 145 711 145 711 2 pad
port 1 ne
rlabel metal1 s 178 4 178 4 2 xpad
port 2 ne
rlabel metal1 s 77 103 77 103 2 a
port 3 ne
rlabel nwell s -2 131 -2 131 2 vdd
rlabel metal2 s 336 466 336 466 2 vdd
port 4 ne
rlabel metal2 s 284 5 284 5 2 vss
port 5 ne
<< end >>
