`celldefine
module and2_b (z, a, b);
  output z;
  input  a;
  input  b;

  and G1 (z, a, b);
endmodule
`endcelldefine
