magic
tech scmos
timestamp 1545344122
<< metal1 >>
rect 18 76 24 79
rect 18 41 24 45
rect 18 0 24 3
use inv_b  0 mag
timestamp 1544839573
transform 1 0 0 0 1 0
box 0 0 24 81
use dlyrc_7ns  1 mag
timestamp 1545342674
transform 1 0 -7 0 1 0
box 31 0 148 79
<< labels >>
rlabel metal1 s 8 29 8 29 2 a
<< end >>
