magic
tech amic5n
magscale 1 2
timestamp 1624397900
<< nwell >>
rect -260 1100 1160 2990
<< ntransistor >>
rect 450 190 570 800
<< ptransistor >>
rect 450 1410 570 2690
<< nselect >>
rect -20 0 920 860
<< pselect >>
rect -15 1340 920 2880
<< ndiffusion >>
rect 210 740 450 800
rect 210 640 270 740
rect 370 640 450 740
rect 210 350 450 640
rect 210 250 270 350
rect 370 250 450 350
rect 210 190 450 250
rect 570 740 810 800
rect 570 640 650 740
rect 750 640 810 740
rect 570 350 810 640
rect 570 250 650 350
rect 750 250 810 350
rect 570 190 810 250
<< pdiffusion >>
rect 210 2630 450 2690
rect 210 2530 270 2630
rect 370 2530 450 2630
rect 210 2430 450 2530
rect 210 2330 270 2430
rect 370 2330 450 2430
rect 210 2230 450 2330
rect 210 2130 270 2230
rect 370 2130 450 2230
rect 210 2030 450 2130
rect 210 1930 270 2030
rect 370 1930 450 2030
rect 210 1830 450 1930
rect 210 1730 270 1830
rect 370 1730 450 1830
rect 210 1630 450 1730
rect 210 1530 270 1630
rect 370 1530 450 1630
rect 210 1410 450 1530
rect 570 2630 810 2690
rect 570 2530 650 2630
rect 750 2530 810 2630
rect 570 2370 810 2530
rect 570 2270 650 2370
rect 750 2270 810 2370
rect 570 2170 810 2270
rect 570 2070 650 2170
rect 750 2070 810 2170
rect 570 1970 810 2070
rect 570 1870 650 1970
rect 750 1870 810 1970
rect 570 1770 810 1870
rect 570 1670 650 1770
rect 750 1670 810 1770
rect 570 1410 810 1670
<< ndcontact >>
rect 270 640 370 740
rect 270 250 370 350
rect 650 640 750 740
rect 650 250 750 350
<< pdcontact >>
rect 270 2530 370 2630
rect 270 2330 370 2430
rect 270 2130 370 2230
rect 270 1930 370 2030
rect 270 1730 370 1830
rect 270 1530 370 1630
rect 650 2530 750 2630
rect 650 2270 750 2370
rect 650 2070 750 2170
rect 650 1870 750 1970
rect 650 1670 750 1770
<< polysilicon >>
rect 450 2690 570 2820
rect 450 1370 570 1410
rect 230 1330 570 1370
rect 230 1230 270 1330
rect 370 1230 570 1330
rect 230 1190 570 1230
rect 450 800 570 1190
rect 450 60 570 190
<< polycontact >>
rect 270 1230 370 1330
<< metal1 >>
rect 0 2790 900 2970
rect 230 2630 410 2790
rect 230 2530 270 2630
rect 370 2530 410 2630
rect 230 2430 410 2530
rect 230 2330 270 2430
rect 370 2330 410 2430
rect 230 2230 410 2330
rect 230 2130 270 2230
rect 370 2130 410 2230
rect 230 2030 410 2130
rect 230 1930 270 2030
rect 370 1930 410 2030
rect 230 1830 410 1930
rect 230 1730 270 1830
rect 370 1730 410 1830
rect 230 1630 410 1730
rect 230 1530 270 1630
rect 370 1530 410 1630
rect 230 1490 410 1530
rect 610 2630 840 2670
rect 610 2530 650 2630
rect 750 2530 840 2630
rect 610 2370 840 2530
rect 610 2270 650 2370
rect 750 2270 840 2370
rect 610 2170 840 2270
rect 610 2070 650 2170
rect 750 2070 840 2170
rect 610 1970 840 2070
rect 610 1870 650 1970
rect 750 1870 840 1970
rect 610 1770 840 1870
rect 610 1670 650 1770
rect 750 1670 840 1770
rect 610 1510 840 1670
rect 230 1330 790 1370
rect 230 1230 270 1330
rect 370 1230 790 1330
rect 230 1190 790 1230
rect 230 740 410 780
rect 230 640 270 740
rect 370 640 410 740
rect 230 350 410 640
rect 230 250 270 350
rect 370 250 410 350
rect 230 90 410 250
rect 610 740 790 1190
rect 610 640 650 740
rect 750 640 790 740
rect 610 350 790 640
rect 610 250 650 350
rect 750 250 790 350
rect 610 210 790 250
rect 0 -90 900 90
<< bb >>
rect 650 1470 750 1570
<< labels >>
flabel metal1 s 190 2830 190 2830 2 FreeSans 800 0 0 0 vdd
port 1 ne
flabel metal1 s 10 10 10 10 2 FreeSans 800 0 0 0 vss
port 2 ne
flabel metal1 s 670 1570 670 1570 2 FreeSans 800 0 0 0 z
port 0 ne
flabel nwell 70 1115 70 1115 2 FreeSans 800 0 0 0 vdd
<< properties >>
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
