`celldefine
module tie0_b (z);
  output z;

  assign z = 1'b0;
endmodule
`endcelldefine
