magic
tech amic5n
timestamp 1608317706
<< poly2capcontact >>
rect 875 515 1405 625
<< poly2cap >>
rect 810 240 1470 900
<< psubstratepdiff >>
rect 1890 390 2250 690
<< polysilicon >>
rect 660 60 1620 1050
<< psubstratepcontact >>
rect 2045 515 2095 565
<< polycontact >>
rect 695 95 745 145
<< polycontact >>
rect 845 95 895 145
<< polycontact >>
rect 995 95 1045 145
<< polycontact >>
rect 1145 95 1195 145
<< polycontact >>
rect 1295 95 1345 145
<< polycontact >>
rect 1445 95 1495 145
<< metal1 >>
rect 1260 630 1410 810
rect 2010 180 2130 600
rect 660 0 1620 180
rect 1890 0 2250 180
<< labels >>
flabel metal1 s 1350 720 1350 720 2 FreeSans 400 0 0 0 n2x
port 2 ne
flabel metal1  2070 60 2070 60 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 1080 30 1080 30 2 FreeSans 400 0 0 0 n2
port 5 ne
<< checkpaint >>
rect -10 -10 2260 1060
<< end >>
