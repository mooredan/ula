magic
tech amic5n
timestamp 1606782623
<< error_p >>
rect -3800 -190 -3780 -150
rect -3930 -210 -3780 -190
rect -3740 -250 -3720 -190
<< nwell >>
rect -4220 640 -3620 2100
rect 570 760 1290 2320
<< ntransistor >>
rect -3950 -100 -3890 450
rect 900 10 960 580
rect -3950 -460 -3890 -300
<< ptransistor >>
rect -3950 790 -3890 1940
rect 900 940 960 2140
<< nselect >>
rect -4100 -130 -3460 530
rect 690 -50 1170 640
rect -4100 -540 -3730 -270
<< pselect >>
rect -4100 760 -3740 1970
rect 690 880 1170 2200
<< ndiffusion >>
rect 750 545 900 580
rect 750 495 785 545
rect 835 495 900 545
rect -4070 420 -3950 450
rect -4070 370 -4040 420
rect -3990 370 -3950 420
rect -4070 -100 -3950 370
rect -3890 420 -3770 450
rect -3890 370 -3850 420
rect -3800 370 -3770 420
rect -3890 -20 -3770 370
rect -3890 -70 -3850 -20
rect -3800 -70 -3770 -20
rect -3890 -100 -3770 -70
rect -3670 420 -3510 470
rect -3670 370 -3640 420
rect -3590 370 -3510 420
rect -3670 -100 -3510 370
rect 750 395 900 495
rect 750 345 785 395
rect 835 345 900 395
rect 750 245 900 345
rect 750 195 785 245
rect 835 195 900 245
rect 750 95 900 195
rect 750 45 785 95
rect 835 45 900 95
rect 750 10 900 45
rect 960 545 1110 580
rect 960 495 1025 545
rect 1075 495 1110 545
rect 960 335 1110 495
rect 960 285 1025 335
rect 1075 285 1110 335
rect 960 155 1110 285
rect 960 105 1025 155
rect 1075 105 1110 155
rect 960 10 1110 105
rect -4070 -330 -3950 -300
rect -4070 -380 -4040 -330
rect -3990 -380 -3950 -330
rect -4070 -460 -3950 -380
rect -3890 -330 -3770 -300
rect -3890 -380 -3850 -330
rect -3800 -380 -3770 -330
rect -3890 -460 -3770 -380
<< pdiffusion >>
rect 750 2105 900 2140
rect 750 2055 785 2105
rect 835 2055 900 2105
rect -4070 1910 -3950 1940
rect -4070 1860 -4040 1910
rect -3990 1860 -3950 1910
rect -4070 790 -3950 1860
rect -3890 1910 -3770 1940
rect -3890 1860 -3850 1910
rect -3800 1860 -3770 1910
rect -3890 790 -3770 1860
rect 750 1925 900 2055
rect 750 1875 785 1925
rect 835 1875 900 1925
rect 750 1775 900 1875
rect 750 1725 785 1775
rect 835 1725 900 1775
rect 750 1625 900 1725
rect 750 1575 785 1625
rect 835 1575 900 1625
rect 750 1475 900 1575
rect 750 1425 785 1475
rect 835 1425 900 1475
rect 750 1325 900 1425
rect 750 1275 785 1325
rect 835 1275 900 1325
rect 750 1175 900 1275
rect 750 1125 785 1175
rect 835 1125 900 1175
rect 750 1025 900 1125
rect 750 975 785 1025
rect 835 975 900 1025
rect 750 940 900 975
rect 960 2045 1110 2140
rect 960 1995 1025 2045
rect 1075 1995 1110 2045
rect 960 1895 1110 1995
rect 960 1845 1025 1895
rect 1075 1845 1110 1895
rect 960 1715 1110 1845
rect 960 1665 1025 1715
rect 1075 1665 1110 1715
rect 960 1535 1110 1665
rect 960 1485 1025 1535
rect 1075 1485 1110 1535
rect 960 1355 1110 1485
rect 960 1305 1025 1355
rect 1075 1305 1110 1355
rect 960 1175 1110 1305
rect 960 1125 1025 1175
rect 1075 1125 1110 1175
rect 960 1025 1110 1125
rect 960 975 1025 1025
rect 1075 975 1110 1025
rect 960 940 1110 975
<< ndcontact >>
rect 785 495 835 545
rect -4040 370 -3990 420
rect -3850 370 -3800 420
rect -3850 -70 -3800 -20
rect -3640 370 -3590 420
rect 785 345 835 395
rect 785 195 835 245
rect 785 45 835 95
rect 1025 495 1075 545
rect 1025 285 1075 335
rect 1025 105 1075 155
rect -4040 -380 -3990 -330
rect -3850 -380 -3800 -330
<< pdcontact >>
rect 785 2055 835 2105
rect -4040 1860 -3990 1910
rect -3850 1860 -3800 1910
rect 785 1875 835 1925
rect 785 1725 835 1775
rect 785 1575 835 1625
rect 785 1425 835 1475
rect 785 1275 835 1325
rect 785 1125 835 1175
rect 785 975 835 1025
rect 1025 1995 1075 2045
rect 1025 1845 1075 1895
rect 1025 1665 1075 1715
rect 1025 1485 1075 1535
rect 1025 1305 1075 1355
rect 1025 1125 1075 1175
rect 1025 975 1075 1025
<< polysilicon >>
rect -3950 2070 -3890 2290
rect 900 2140 960 2205
rect -3950 1940 -3890 2010
rect 900 850 960 940
rect -3950 645 -3890 790
rect 750 785 960 850
rect 750 735 815 785
rect 865 735 960 785
rect 750 670 960 735
rect -4060 625 -3890 645
rect -4060 575 -4040 625
rect -3990 575 -3890 625
rect 900 580 960 670
rect -4060 555 -3890 575
rect -3950 450 -3890 555
rect 900 -55 960 10
rect -3950 -170 -3890 -100
rect -3950 -300 -3890 -230
rect -3950 -530 -3890 -460
<< polycontact >>
rect 815 735 865 785
rect -4040 575 -3990 625
<< metal1 >>
rect 690 2170 1170 2260
rect 750 2105 870 2170
rect 750 2055 785 2105
rect 835 2055 870 2105
rect -4060 1990 -3780 2050
rect -4060 1910 -3970 1990
rect -4060 1860 -4040 1910
rect -3990 1860 -3970 1910
rect -4060 870 -3970 1860
rect -3870 1910 -3780 1930
rect -3870 1860 -3850 1910
rect -3800 1860 -3780 1910
rect -4060 625 -3970 645
rect -4060 575 -4040 625
rect -3990 575 -3970 625
rect -4060 555 -3970 575
rect -4060 420 -3970 440
rect -4060 370 -4040 420
rect -3990 370 -3970 420
rect -4060 -150 -3970 370
rect -3870 420 -3780 1860
rect 750 1925 870 2055
rect 750 1875 785 1925
rect 835 1875 870 1925
rect 750 1775 870 1875
rect 750 1725 785 1775
rect 835 1725 870 1775
rect 750 1625 870 1725
rect 750 1575 785 1625
rect 835 1575 870 1625
rect 750 1475 870 1575
rect 750 1425 785 1475
rect 835 1425 870 1475
rect 750 1325 870 1425
rect 750 1275 785 1325
rect 835 1275 870 1325
rect 750 1175 870 1275
rect 750 1125 785 1175
rect 835 1125 870 1175
rect 750 1025 870 1125
rect 750 975 785 1025
rect 835 975 870 1025
rect 750 940 870 975
rect 990 2045 1110 2080
rect 990 1995 1025 2045
rect 1075 1995 1110 2045
rect 990 1895 1110 1995
rect 990 1845 1025 1895
rect 1075 1845 1110 1895
rect 990 1715 1110 1845
rect 990 1665 1025 1715
rect 1075 1665 1110 1715
rect 990 1535 1110 1665
rect 990 1485 1025 1535
rect 1075 1485 1110 1535
rect 990 1355 1110 1485
rect 990 1305 1025 1355
rect 1075 1305 1110 1355
rect 990 1175 1110 1305
rect 990 1125 1025 1175
rect 1075 1125 1110 1175
rect 990 1025 1110 1125
rect 990 975 1025 1025
rect 1075 975 1110 1025
rect 780 785 900 820
rect 780 735 815 785
rect 865 735 900 785
rect 780 700 900 735
rect 750 545 870 580
rect 750 495 785 545
rect 835 495 870 545
rect -3870 370 -3850 420
rect -3800 370 -3780 420
rect -3870 -20 -3780 370
rect -3660 420 -3570 440
rect -3660 370 -3640 420
rect -3590 370 -3570 420
rect -3660 350 -3570 370
rect 750 395 870 495
rect 750 345 785 395
rect 835 345 870 395
rect 750 245 870 345
rect 750 195 785 245
rect 835 195 870 245
rect 750 95 870 195
rect 750 45 785 95
rect 835 45 870 95
rect 990 545 1110 975
rect 990 495 1025 545
rect 1075 495 1110 545
rect 990 335 1110 495
rect 990 285 1025 335
rect 1075 285 1110 335
rect 990 155 1110 285
rect 990 105 1025 155
rect 1075 105 1110 155
rect 990 70 1110 105
rect 750 -20 870 45
rect -3870 -70 -3850 -20
rect -3800 -70 -3780 -20
rect -3870 -90 -3780 -70
rect 690 -110 1170 -20
rect -4060 -210 -3780 -150
rect -3740 -250 -3590 -190
rect -4060 -330 -3970 -310
rect -4060 -380 -4040 -330
rect -3990 -380 -3970 -330
rect -4060 -400 -3970 -380
rect -3870 -330 -3780 -250
rect -3870 -380 -3850 -330
rect -3800 -380 -3780 -330
rect -3870 -400 -3780 -380
rect -2320 -785 -2230 -645
rect -2320 -835 -2300 -785
rect -2250 -835 -2230 -785
rect -2320 -945 -2230 -835
rect -2320 -995 -2300 -945
rect -2250 -995 -2230 -945
rect -2320 -1075 -2230 -995
rect -2170 -785 -2080 -655
rect -2170 -835 -2150 -785
rect -2100 -835 -2080 -785
rect -2170 -945 -2080 -835
rect -2170 -995 -2150 -945
rect -2100 -995 -2080 -945
rect -2170 -1055 -2080 -995
<< via1 >>
rect -2300 -835 -2250 -785
rect -2300 -995 -2250 -945
rect -2150 -835 -2100 -785
rect -2150 -995 -2100 -945
<< metal2 >>
rect -2960 2635 330 2725
rect -2960 2475 330 2565
rect -2960 2315 330 2405
rect -2960 2155 330 2245
rect -4200 1995 -3040 2085
rect -2960 1995 330 2085
rect -2960 1835 330 1925
rect -2960 1675 330 1765
rect -2960 1515 330 1605
rect -2960 1355 330 1445
rect -2960 1195 330 1285
rect -2960 1035 330 1125
rect -2960 875 330 965
rect -3090 715 330 805
rect -3090 555 330 645
rect -2960 395 330 485
rect -2960 235 330 325
rect -2960 75 330 165
rect -2960 -85 330 5
rect -4200 -245 -3040 -155
rect -2960 -245 330 -155
rect -2960 -405 330 -315
rect -2960 -565 330 -475
rect -2910 -785 -1830 -765
rect -2910 -835 -2815 -785
rect -2765 -835 -2655 -785
rect -2605 -835 -2300 -785
rect -2250 -835 -2150 -785
rect -2100 -835 -1830 -785
rect -2910 -855 -1830 -835
rect -2910 -945 -1830 -925
rect -2910 -995 -2815 -945
rect -2765 -995 -2655 -945
rect -2605 -995 -2300 -945
rect -2250 -995 -2150 -945
rect -2100 -995 -1830 -945
rect -2910 -1015 -1830 -995
<< via2 >>
rect -2815 -835 -2765 -785
rect -2655 -835 -2605 -785
rect -2815 -995 -2765 -945
rect -2655 -995 -2605 -945
<< metal3 >>
rect -2830 -765 -2750 -695
rect -2670 -765 -2590 -695
rect -2835 -785 -2745 -765
rect -2835 -835 -2815 -785
rect -2765 -835 -2745 -785
rect -2835 -855 -2745 -835
rect -2675 -785 -2585 -765
rect -2675 -835 -2655 -785
rect -2605 -835 -2585 -785
rect -2675 -855 -2585 -835
rect -2830 -925 -2750 -855
rect -2670 -925 -2590 -855
rect -2835 -945 -2745 -925
rect -2835 -995 -2815 -945
rect -2765 -995 -2745 -945
rect -2835 -1015 -2745 -995
rect -2675 -945 -2585 -925
rect -2675 -995 -2655 -945
rect -2605 -995 -2585 -945
rect -2675 -1015 -2585 -995
rect -2830 -1075 -2750 -1015
rect -2670 -1075 -2590 -1015
<< labels >>
flabel nwell 690 820 690 820 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 720 -80 720 -80 2 FreeSans 400 0 0 0 vss
port 4 ne
flabel metal1 s 720 2200 720 2200 2 FreeSans 400 0 0 0 vdd
port 3 ne
flabel metal1 s 1050 700 1050 700 2 FreeSans 400 0 0 0 z
port 1 ne
flabel metal1 s 840 760 840 760 2 FreeSans 400 0 0 0 a
port 2 ne
<< end >>
