magic
tech amic5n
timestamp 1622307144
<< nwell >>
rect -130 550 730 1495
<< ntransistor >>
rect 165 275 225 400
rect 375 95 435 400
<< ptransistor >>
rect 165 800 225 985
rect 375 700 435 1345
<< nselect >>
rect -10 0 610 430
<< pselect >>
rect -10 670 610 1440
<< ndiffusion >>
rect 45 365 165 400
rect 45 315 75 365
rect 125 315 165 365
rect 45 275 165 315
rect 225 370 375 400
rect 225 320 285 370
rect 335 320 375 370
rect 225 275 375 320
rect 255 175 375 275
rect 255 125 285 175
rect 335 125 375 175
rect 255 95 375 125
rect 435 370 555 400
rect 435 320 475 370
rect 525 320 555 370
rect 435 175 555 320
rect 435 125 475 175
rect 525 125 555 175
rect 435 95 555 125
<< pdiffusion >>
rect 255 1315 375 1345
rect 255 1265 285 1315
rect 335 1265 375 1315
rect 255 1215 375 1265
rect 255 1165 285 1215
rect 335 1165 375 1215
rect 255 1115 375 1165
rect 255 1065 285 1115
rect 335 1065 375 1115
rect 255 1015 375 1065
rect 255 985 285 1015
rect 45 915 165 985
rect 45 865 75 915
rect 125 865 165 915
rect 45 800 165 865
rect 225 965 285 985
rect 335 965 375 1015
rect 225 915 375 965
rect 225 865 285 915
rect 335 865 375 915
rect 225 815 375 865
rect 225 800 285 815
rect 255 765 285 800
rect 335 765 375 815
rect 255 700 375 765
rect 435 1315 555 1345
rect 435 1265 475 1315
rect 525 1265 555 1315
rect 435 1180 555 1265
rect 435 1130 475 1180
rect 525 1130 555 1180
rect 435 1080 555 1130
rect 435 1030 475 1080
rect 525 1030 555 1080
rect 435 980 555 1030
rect 435 930 475 980
rect 525 930 555 980
rect 435 880 555 930
rect 435 830 475 880
rect 525 830 555 880
rect 435 780 555 830
rect 435 730 475 780
rect 525 730 555 780
rect 435 700 555 730
<< ndcontact >>
rect 75 315 125 365
rect 285 320 335 370
rect 285 125 335 175
rect 475 320 525 370
rect 475 125 525 175
<< pdcontact >>
rect 285 1265 335 1315
rect 285 1165 335 1215
rect 285 1065 335 1115
rect 75 865 125 915
rect 285 965 335 1015
rect 285 865 335 915
rect 285 765 335 815
rect 475 1265 525 1315
rect 475 1130 525 1180
rect 475 1030 525 1080
rect 475 930 525 980
rect 475 830 525 880
rect 475 730 525 780
<< polysilicon >>
rect 375 1345 435 1410
rect 105 1145 225 1165
rect 105 1095 125 1145
rect 175 1095 225 1145
rect 105 1075 225 1095
rect 165 985 225 1075
rect 165 755 225 800
rect 125 695 225 755
rect 125 480 185 695
rect 375 630 435 700
rect 265 610 435 630
rect 265 560 285 610
rect 335 560 435 610
rect 265 540 435 560
rect 125 420 225 480
rect 165 400 225 420
rect 375 400 435 540
rect 165 210 225 275
rect 375 30 435 95
<< polycontact >>
rect 125 1095 175 1145
rect 285 560 335 610
<< metal1 >>
rect 0 1395 600 1485
rect 265 1315 355 1395
rect 265 1265 285 1315
rect 335 1265 355 1315
rect 265 1215 355 1265
rect 265 1165 285 1215
rect 335 1165 355 1215
rect 30 1145 195 1165
rect 30 1095 125 1145
rect 175 1095 195 1145
rect 30 1075 195 1095
rect 265 1115 355 1165
rect 265 1065 285 1115
rect 335 1065 355 1115
rect 265 1015 355 1065
rect 265 965 285 1015
rect 335 965 355 1015
rect 55 915 145 945
rect 55 865 75 915
rect 125 865 145 915
rect 55 630 145 865
rect 265 915 355 965
rect 265 865 285 915
rect 335 865 355 915
rect 265 815 355 865
rect 265 765 285 815
rect 335 765 355 815
rect 265 745 355 765
rect 455 1315 545 1335
rect 455 1265 475 1315
rect 525 1265 545 1315
rect 455 1180 545 1265
rect 455 1130 475 1180
rect 525 1130 545 1180
rect 455 1080 545 1130
rect 455 1030 475 1080
rect 525 1030 545 1080
rect 455 980 545 1030
rect 455 930 475 980
rect 525 930 545 980
rect 455 880 545 930
rect 455 830 475 880
rect 525 830 545 880
rect 455 780 545 830
rect 455 730 475 780
rect 525 730 545 780
rect 455 685 545 730
rect 55 610 355 630
rect 55 560 285 610
rect 335 560 355 610
rect 55 540 355 560
rect 55 365 145 540
rect 455 435 570 685
rect 55 315 75 365
rect 125 315 145 365
rect 55 285 145 315
rect 265 370 355 390
rect 265 320 285 370
rect 335 320 355 370
rect 265 175 355 320
rect 265 125 285 175
rect 335 125 355 175
rect 265 45 355 125
rect 455 370 545 435
rect 455 320 475 370
rect 525 320 545 370
rect 455 175 545 320
rect 455 125 475 175
rect 525 125 545 175
rect 455 105 545 125
rect 0 -45 600 45
<< labels >>
flabel metal1 s 255 -25 255 -25 2 FreeSans 400 0 0 0 vss
port 12 ne
flabel metal1 s 245 1415 245 1415 2 FreeSans 400 0 0 0 vdd
port 11 ne
flabel nwell 545 600 545 600 2 FreeSans 400 0 0 0 vdd
flabel metal1 s 485 470 485 470 2 FreeSans 400 0 0 0 z
port 20 ne
flabel metal1 s 125 1085 125 1085 2 FreeSans 400 0 0 0 a
port 7 ne
<< end >>
