magic
tech amic5n
timestamp 1608317708
<< checkpaint >>
rect -10 -10 10 10
<< end >>
