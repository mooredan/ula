magic
tech scmos
magscale 1 2
timestamp 1570494029
<< error_p >>
rect 20 1320 22 1322
rect 578 1320 580 1322
rect 18 1318 20 1320
rect 580 1318 582 1320
rect 80 1296 90 1298
rect 78 1294 90 1296
rect 510 1296 520 1298
rect 510 1294 522 1296
rect 80 1290 82 1294
rect 518 1290 520 1294
rect 80 1286 90 1290
rect 78 1284 90 1286
rect 510 1286 520 1290
rect 510 1284 522 1286
rect 80 1282 82 1284
rect 518 1282 520 1284
rect 82 1280 84 1282
rect 516 1280 518 1282
rect 50 1279 52 1280
rect 548 1279 550 1280
rect 48 1277 50 1278
rect 550 1277 552 1278
rect 50 1259 52 1260
rect 548 1259 550 1260
rect 48 1257 50 1258
rect 550 1257 552 1258
rect 96 1242 98 1244
rect 502 1242 504 1244
rect 94 1240 96 1242
rect 504 1240 506 1242
rect 50 1239 52 1240
rect 548 1239 550 1240
rect 48 1237 50 1238
rect 550 1237 552 1238
rect 50 1219 52 1220
rect 548 1219 550 1220
rect 48 1217 50 1218
rect 550 1217 552 1218
rect 50 1199 52 1200
rect 548 1199 550 1200
rect 48 1197 50 1198
rect 550 1197 552 1198
rect 94 1180 96 1182
rect 504 1180 506 1182
rect 50 1179 52 1180
rect 96 1178 98 1180
rect 502 1178 504 1180
rect 548 1179 550 1180
rect 48 1177 50 1178
rect 550 1177 552 1178
rect 50 1159 52 1160
rect 548 1159 550 1160
rect 48 1157 50 1158
rect 550 1157 552 1158
rect 50 1139 52 1140
rect 548 1139 550 1140
rect 48 1137 50 1138
rect 550 1137 552 1138
rect 50 1119 52 1120
rect 548 1119 550 1120
rect 48 1117 50 1118
rect 550 1117 552 1118
rect 96 1114 98 1116
rect 502 1114 504 1116
rect 94 1112 96 1114
rect 504 1112 506 1114
rect 50 1099 52 1100
rect 548 1099 550 1100
rect 48 1097 50 1098
rect 550 1097 552 1098
rect 50 1079 52 1080
rect 548 1079 550 1080
rect 48 1077 50 1078
rect 550 1077 552 1078
rect 50 1059 52 1060
rect 548 1059 550 1060
rect 48 1057 50 1058
rect 550 1057 552 1058
rect 94 1052 96 1054
rect 504 1052 506 1054
rect 96 1050 98 1052
rect 502 1050 504 1052
rect 50 1039 52 1040
rect 548 1039 550 1040
rect 48 1037 50 1038
rect 550 1037 552 1038
rect 50 1019 52 1020
rect 548 1019 550 1020
rect 48 1017 50 1018
rect 550 1017 552 1018
rect 50 999 52 1000
rect 548 999 550 1000
rect 48 997 50 998
rect 550 997 552 998
rect 96 984 98 986
rect 502 984 504 986
rect 94 982 96 984
rect 504 982 506 984
rect 50 979 52 980
rect 548 979 550 980
rect 48 977 50 978
rect 550 977 552 978
rect 50 959 52 960
rect 548 959 550 960
rect 48 957 50 958
rect 550 957 552 958
rect 50 939 52 940
rect 548 939 550 940
rect 48 937 50 938
rect 550 937 552 938
rect 94 922 96 924
rect 504 922 506 924
rect 96 920 98 922
rect 502 920 504 922
rect 50 919 52 920
rect 548 919 550 920
rect 48 917 50 918
rect 550 917 552 918
rect 50 899 52 900
rect 548 899 550 900
rect 48 897 50 898
rect 550 897 552 898
rect 62 873 64 875
rect 536 873 538 875
rect 60 871 62 873
rect 538 871 540 873
rect 32 828 34 830
rect 62 828 64 830
rect 92 828 94 830
rect 122 828 124 830
rect 152 828 154 830
rect 182 828 184 830
rect 212 828 214 830
rect 386 828 388 830
rect 416 828 418 830
rect 446 828 448 830
rect 476 828 478 830
rect 506 828 508 830
rect 536 828 538 830
rect 566 828 568 830
rect 34 826 36 828
rect 40 826 42 828
rect 64 826 66 828
rect 70 826 72 828
rect 94 826 96 828
rect 100 826 102 828
rect 124 826 126 828
rect 130 826 132 828
rect 154 826 156 828
rect 160 826 162 828
rect 184 826 186 828
rect 190 826 192 828
rect 214 826 216 828
rect 220 826 222 828
rect 378 826 380 828
rect 384 826 386 828
rect 408 826 410 828
rect 414 826 416 828
rect 438 826 440 828
rect 444 826 446 828
rect 468 826 470 828
rect 474 826 476 828
rect 498 826 500 828
rect 504 826 506 828
rect 528 826 530 828
rect 534 826 536 828
rect 558 826 560 828
rect 564 826 566 828
rect 42 824 44 826
rect 72 824 74 826
rect 102 824 104 826
rect 132 824 134 826
rect 162 824 164 826
rect 192 824 194 826
rect 222 824 224 826
rect 376 824 378 826
rect 406 824 408 826
rect 436 824 438 826
rect 466 824 468 826
rect 496 824 498 826
rect 526 824 528 826
rect 556 824 558 826
rect 42 818 44 820
rect 72 818 74 820
rect 102 818 104 820
rect 132 818 134 820
rect 162 818 164 820
rect 192 818 194 820
rect 222 818 224 820
rect 376 818 378 820
rect 406 818 408 820
rect 436 818 438 820
rect 466 818 468 820
rect 496 818 498 820
rect 526 818 528 820
rect 556 818 558 820
rect 34 816 36 818
rect 40 816 42 818
rect 64 816 66 818
rect 70 816 72 818
rect 94 816 96 818
rect 100 816 102 818
rect 124 816 126 818
rect 130 816 132 818
rect 154 816 156 818
rect 160 816 162 818
rect 184 816 186 818
rect 190 816 192 818
rect 214 816 216 818
rect 220 816 222 818
rect 378 816 380 818
rect 384 816 386 818
rect 408 816 410 818
rect 414 816 416 818
rect 438 816 440 818
rect 444 816 446 818
rect 468 816 470 818
rect 474 816 476 818
rect 498 816 500 818
rect 504 816 506 818
rect 528 816 530 818
rect 534 816 536 818
rect 558 816 560 818
rect 564 816 566 818
rect 32 814 34 816
rect 62 814 64 816
rect 92 814 94 816
rect 122 814 124 816
rect 152 814 154 816
rect 182 814 184 816
rect 212 814 214 816
rect 386 814 388 816
rect 416 814 418 816
rect 446 814 448 816
rect 476 814 478 816
rect 506 814 508 816
rect 536 814 538 816
rect 566 814 568 816
rect 32 808 34 810
rect 62 808 64 810
rect 92 808 94 810
rect 122 808 124 810
rect 152 808 154 810
rect 182 808 184 810
rect 212 808 214 810
rect 386 808 388 810
rect 416 808 418 810
rect 446 808 448 810
rect 476 808 478 810
rect 506 808 508 810
rect 536 808 538 810
rect 566 808 568 810
rect 34 806 36 808
rect 40 806 42 808
rect 64 806 66 808
rect 70 806 72 808
rect 94 806 96 808
rect 100 806 102 808
rect 124 806 126 808
rect 130 806 132 808
rect 154 806 156 808
rect 160 806 162 808
rect 184 806 186 808
rect 190 806 192 808
rect 214 806 216 808
rect 220 806 222 808
rect 378 806 380 808
rect 384 806 386 808
rect 408 806 410 808
rect 414 806 416 808
rect 438 806 440 808
rect 444 806 446 808
rect 468 806 470 808
rect 474 806 476 808
rect 498 806 500 808
rect 504 806 506 808
rect 528 806 530 808
rect 534 806 536 808
rect 558 806 560 808
rect 564 806 566 808
rect 42 804 44 806
rect 72 804 74 806
rect 102 804 104 806
rect 132 804 134 806
rect 162 804 164 806
rect 192 804 194 806
rect 222 804 224 806
rect 376 804 378 806
rect 406 804 408 806
rect 436 804 438 806
rect 466 804 468 806
rect 496 804 498 806
rect 526 804 528 806
rect 556 804 558 806
rect 42 798 44 800
rect 72 798 74 800
rect 102 798 104 800
rect 132 798 134 800
rect 162 798 164 800
rect 192 798 194 800
rect 222 798 224 800
rect 376 798 378 800
rect 406 798 408 800
rect 436 798 438 800
rect 466 798 468 800
rect 496 798 498 800
rect 526 798 528 800
rect 556 798 558 800
rect 34 796 36 798
rect 40 796 42 798
rect 64 796 66 798
rect 70 796 72 798
rect 94 796 96 798
rect 100 796 102 798
rect 124 796 126 798
rect 130 796 132 798
rect 154 796 156 798
rect 160 796 162 798
rect 184 796 186 798
rect 190 796 192 798
rect 214 796 216 798
rect 220 796 222 798
rect 378 796 380 798
rect 384 796 386 798
rect 408 796 410 798
rect 414 796 416 798
rect 438 796 440 798
rect 444 796 446 798
rect 468 796 470 798
rect 474 796 476 798
rect 498 796 500 798
rect 504 796 506 798
rect 528 796 530 798
rect 534 796 536 798
rect 558 796 560 798
rect 564 796 566 798
rect 32 794 34 796
rect 62 794 64 796
rect 92 794 94 796
rect 122 794 124 796
rect 152 794 154 796
rect 182 794 184 796
rect 212 794 214 796
rect 386 794 388 796
rect 416 794 418 796
rect 446 794 448 796
rect 476 794 478 796
rect 506 794 508 796
rect 536 794 538 796
rect 566 794 568 796
rect 32 788 34 790
rect 62 788 64 790
rect 92 788 94 790
rect 122 788 124 790
rect 152 788 154 790
rect 182 788 184 790
rect 212 788 214 790
rect 386 788 388 790
rect 416 788 418 790
rect 446 788 448 790
rect 476 788 478 790
rect 506 788 508 790
rect 536 788 538 790
rect 566 788 568 790
rect 34 786 36 788
rect 40 786 42 788
rect 64 786 66 788
rect 70 786 72 788
rect 94 786 96 788
rect 100 786 102 788
rect 124 786 126 788
rect 130 786 132 788
rect 154 786 156 788
rect 160 786 162 788
rect 184 786 186 788
rect 190 786 192 788
rect 214 786 216 788
rect 220 786 222 788
rect 378 786 380 788
rect 384 786 386 788
rect 408 786 410 788
rect 414 786 416 788
rect 438 786 440 788
rect 444 786 446 788
rect 468 786 470 788
rect 474 786 476 788
rect 498 786 500 788
rect 504 786 506 788
rect 528 786 530 788
rect 534 786 536 788
rect 558 786 560 788
rect 564 786 566 788
rect 42 784 44 786
rect 72 784 74 786
rect 102 784 104 786
rect 132 784 134 786
rect 162 784 164 786
rect 192 784 194 786
rect 222 784 224 786
rect 376 784 378 786
rect 406 784 408 786
rect 436 784 438 786
rect 466 784 468 786
rect 496 784 498 786
rect 526 784 528 786
rect 556 784 558 786
rect 42 778 44 780
rect 72 778 74 780
rect 526 778 528 780
rect 556 778 558 780
rect 34 776 36 778
rect 40 776 42 778
rect 64 776 66 778
rect 70 776 72 778
rect 94 776 96 778
rect 110 776 112 778
rect 124 776 126 778
rect 140 776 142 778
rect 154 776 156 778
rect 170 776 172 778
rect 184 776 186 778
rect 200 776 202 778
rect 214 776 216 778
rect 230 776 232 778
rect 244 776 246 778
rect 260 776 262 778
rect 274 776 276 778
rect 280 776 282 778
rect 318 776 320 778
rect 324 776 326 778
rect 338 776 340 778
rect 354 776 356 778
rect 368 776 370 778
rect 384 776 386 778
rect 398 776 400 778
rect 414 776 416 778
rect 428 776 430 778
rect 444 776 446 778
rect 458 776 460 778
rect 474 776 476 778
rect 488 776 490 778
rect 504 776 506 778
rect 528 776 530 778
rect 534 776 536 778
rect 558 776 560 778
rect 564 776 566 778
rect 32 774 34 776
rect 62 774 64 776
rect 92 774 94 776
rect 112 774 114 776
rect 122 774 124 776
rect 142 774 144 776
rect 152 774 154 776
rect 172 774 174 776
rect 182 774 184 776
rect 202 774 204 776
rect 212 774 214 776
rect 232 774 234 776
rect 242 774 244 776
rect 262 774 264 776
rect 272 774 274 776
rect 282 774 284 776
rect 316 774 318 776
rect 326 774 328 776
rect 336 774 338 776
rect 356 774 358 776
rect 366 774 368 776
rect 386 774 388 776
rect 396 774 398 776
rect 416 774 418 776
rect 426 774 428 776
rect 446 774 448 776
rect 456 774 458 776
rect 476 774 478 776
rect 486 774 488 776
rect 506 774 508 776
rect 536 774 538 776
rect 566 774 568 776
rect 32 768 34 770
rect 62 768 64 770
rect 92 768 94 770
rect 112 768 114 770
rect 122 768 124 770
rect 142 768 144 770
rect 152 768 154 770
rect 172 768 174 770
rect 182 768 184 770
rect 202 768 204 770
rect 212 768 214 770
rect 232 768 234 770
rect 242 768 244 770
rect 262 768 264 770
rect 272 768 274 770
rect 282 768 284 770
rect 316 768 318 770
rect 326 768 328 770
rect 336 768 338 770
rect 356 768 358 770
rect 366 768 368 770
rect 386 768 388 770
rect 396 768 398 770
rect 416 768 418 770
rect 426 768 428 770
rect 446 768 448 770
rect 456 768 458 770
rect 476 768 478 770
rect 486 768 488 770
rect 506 768 508 770
rect 536 768 538 770
rect 566 768 568 770
rect 34 766 36 768
rect 40 766 42 768
rect 64 766 66 768
rect 70 766 72 768
rect 94 766 96 768
rect 110 766 112 768
rect 124 766 126 768
rect 140 766 142 768
rect 154 766 156 768
rect 170 766 172 768
rect 184 766 186 768
rect 200 766 202 768
rect 214 766 216 768
rect 230 766 232 768
rect 244 766 246 768
rect 260 766 262 768
rect 274 766 276 768
rect 280 766 282 768
rect 318 766 320 768
rect 324 766 326 768
rect 338 766 340 768
rect 354 766 356 768
rect 368 766 370 768
rect 384 766 386 768
rect 398 766 400 768
rect 414 766 416 768
rect 428 766 430 768
rect 444 766 446 768
rect 458 766 460 768
rect 474 766 476 768
rect 488 766 490 768
rect 504 766 506 768
rect 528 766 530 768
rect 534 766 536 768
rect 558 766 560 768
rect 564 766 566 768
rect 42 764 44 766
rect 72 764 74 766
rect 526 764 528 766
rect 556 764 558 766
rect 42 758 44 760
rect 72 758 74 760
rect 102 758 104 760
rect 132 758 134 760
rect 162 758 164 760
rect 192 758 194 760
rect 222 758 224 760
rect 376 758 378 760
rect 406 758 408 760
rect 436 758 438 760
rect 466 758 468 760
rect 496 758 498 760
rect 526 758 528 760
rect 556 758 558 760
rect 34 756 36 758
rect 40 756 42 758
rect 64 756 66 758
rect 70 756 72 758
rect 94 756 96 758
rect 100 756 102 758
rect 124 756 126 758
rect 130 756 132 758
rect 154 756 156 758
rect 160 756 162 758
rect 184 756 186 758
rect 190 756 192 758
rect 214 756 216 758
rect 220 756 222 758
rect 378 756 380 758
rect 384 756 386 758
rect 408 756 410 758
rect 414 756 416 758
rect 438 756 440 758
rect 444 756 446 758
rect 468 756 470 758
rect 474 756 476 758
rect 498 756 500 758
rect 504 756 506 758
rect 528 756 530 758
rect 534 756 536 758
rect 558 756 560 758
rect 564 756 566 758
rect 32 754 34 756
rect 62 754 64 756
rect 92 754 94 756
rect 122 754 124 756
rect 152 754 154 756
rect 182 754 184 756
rect 212 754 214 756
rect 386 754 388 756
rect 416 754 418 756
rect 446 754 448 756
rect 476 754 478 756
rect 506 754 508 756
rect 536 754 538 756
rect 566 754 568 756
rect 32 748 34 750
rect 62 748 64 750
rect 92 748 94 750
rect 122 748 124 750
rect 152 748 154 750
rect 182 748 184 750
rect 212 748 214 750
rect 386 748 388 750
rect 416 748 418 750
rect 446 748 448 750
rect 476 748 478 750
rect 506 748 508 750
rect 536 748 538 750
rect 566 748 568 750
rect 34 746 36 748
rect 40 746 42 748
rect 64 746 66 748
rect 70 746 72 748
rect 94 746 96 748
rect 100 746 102 748
rect 124 746 126 748
rect 130 746 132 748
rect 154 746 156 748
rect 160 746 162 748
rect 184 746 186 748
rect 190 746 192 748
rect 214 746 216 748
rect 220 746 222 748
rect 378 746 380 748
rect 384 746 386 748
rect 408 746 410 748
rect 414 746 416 748
rect 438 746 440 748
rect 444 746 446 748
rect 468 746 470 748
rect 474 746 476 748
rect 498 746 500 748
rect 504 746 506 748
rect 528 746 530 748
rect 534 746 536 748
rect 558 746 560 748
rect 564 746 566 748
rect 42 744 44 746
rect 72 744 74 746
rect 102 744 104 746
rect 132 744 134 746
rect 162 744 164 746
rect 192 744 194 746
rect 222 744 224 746
rect 376 744 378 746
rect 406 744 408 746
rect 436 744 438 746
rect 466 744 468 746
rect 496 744 498 746
rect 526 744 528 746
rect 556 744 558 746
rect 222 738 224 740
rect 376 738 378 740
rect 220 736 222 738
rect 378 736 380 738
rect 220 726 222 728
rect 378 726 380 728
rect 222 724 224 726
rect 376 724 378 726
rect 42 718 44 720
rect 72 718 74 720
rect 102 718 104 720
rect 132 718 134 720
rect 162 718 164 720
rect 192 718 194 720
rect 222 718 224 720
rect 376 718 378 720
rect 406 718 408 720
rect 436 718 438 720
rect 466 718 468 720
rect 496 718 498 720
rect 526 718 528 720
rect 556 718 558 720
rect 34 716 36 718
rect 40 716 42 718
rect 64 716 66 718
rect 70 716 72 718
rect 94 716 96 718
rect 100 716 102 718
rect 124 716 126 718
rect 130 716 132 718
rect 154 716 156 718
rect 160 716 162 718
rect 184 716 186 718
rect 190 716 192 718
rect 214 716 216 718
rect 220 716 222 718
rect 378 716 380 718
rect 384 716 386 718
rect 408 716 410 718
rect 414 716 416 718
rect 438 716 440 718
rect 444 716 446 718
rect 468 716 470 718
rect 474 716 476 718
rect 498 716 500 718
rect 504 716 506 718
rect 528 716 530 718
rect 534 716 536 718
rect 558 716 560 718
rect 564 716 566 718
rect 32 714 34 716
rect 62 714 64 716
rect 92 714 94 716
rect 122 714 124 716
rect 152 714 154 716
rect 182 714 184 716
rect 212 714 214 716
rect 386 714 388 716
rect 416 714 418 716
rect 446 714 448 716
rect 476 714 478 716
rect 506 714 508 716
rect 536 714 538 716
rect 566 714 568 716
rect 32 708 34 710
rect 62 708 64 710
rect 92 708 94 710
rect 122 708 124 710
rect 152 708 154 710
rect 182 708 184 710
rect 212 708 214 710
rect 386 708 388 710
rect 416 708 418 710
rect 446 708 448 710
rect 476 708 478 710
rect 506 708 508 710
rect 536 708 538 710
rect 566 708 568 710
rect 34 706 36 708
rect 40 706 42 708
rect 64 706 66 708
rect 70 706 72 708
rect 94 706 96 708
rect 100 706 102 708
rect 124 706 126 708
rect 130 706 132 708
rect 154 706 156 708
rect 160 706 162 708
rect 184 706 186 708
rect 190 706 192 708
rect 214 706 216 708
rect 220 706 222 708
rect 378 706 380 708
rect 384 706 386 708
rect 408 706 410 708
rect 414 706 416 708
rect 438 706 440 708
rect 444 706 446 708
rect 468 706 470 708
rect 474 706 476 708
rect 498 706 500 708
rect 504 706 506 708
rect 528 706 530 708
rect 534 706 536 708
rect 558 706 560 708
rect 564 706 566 708
rect 42 704 44 706
rect 72 704 74 706
rect 102 704 104 706
rect 132 704 134 706
rect 162 704 164 706
rect 192 704 194 706
rect 222 704 224 706
rect 376 704 378 706
rect 406 704 408 706
rect 436 704 438 706
rect 466 704 468 706
rect 496 704 498 706
rect 526 704 528 706
rect 556 704 558 706
rect 42 698 44 700
rect 72 698 74 700
rect 102 698 104 700
rect 132 698 134 700
rect 162 698 164 700
rect 192 698 194 700
rect 222 698 224 700
rect 376 698 378 700
rect 406 698 408 700
rect 436 698 438 700
rect 466 698 468 700
rect 496 698 498 700
rect 526 698 528 700
rect 556 698 558 700
rect 34 696 36 698
rect 40 696 42 698
rect 64 696 66 698
rect 70 696 72 698
rect 94 696 96 698
rect 100 696 102 698
rect 124 696 126 698
rect 130 696 132 698
rect 154 696 156 698
rect 160 696 162 698
rect 184 696 186 698
rect 190 696 192 698
rect 214 696 216 698
rect 220 696 222 698
rect 378 696 380 698
rect 384 696 386 698
rect 408 696 410 698
rect 414 696 416 698
rect 438 696 440 698
rect 444 696 446 698
rect 468 696 470 698
rect 474 696 476 698
rect 498 696 500 698
rect 504 696 506 698
rect 528 696 530 698
rect 534 696 536 698
rect 558 696 560 698
rect 564 696 566 698
rect 32 694 34 696
rect 62 694 64 696
rect 92 694 94 696
rect 122 694 124 696
rect 152 694 154 696
rect 182 694 184 696
rect 212 694 214 696
rect 386 694 388 696
rect 416 694 418 696
rect 446 694 448 696
rect 476 694 478 696
rect 506 694 508 696
rect 536 694 538 696
rect 566 694 568 696
rect 32 644 34 646
rect 62 644 64 646
rect 92 644 94 646
rect 122 644 124 646
rect 152 644 154 646
rect 182 644 184 646
rect 416 644 418 646
rect 446 644 448 646
rect 476 644 478 646
rect 506 644 508 646
rect 536 644 538 646
rect 566 644 568 646
rect 34 642 36 644
rect 40 642 42 644
rect 64 642 66 644
rect 70 642 72 644
rect 94 642 96 644
rect 100 642 102 644
rect 124 642 126 644
rect 130 642 132 644
rect 154 642 156 644
rect 160 642 162 644
rect 184 642 186 644
rect 414 642 416 644
rect 438 642 440 644
rect 444 642 446 644
rect 468 642 470 644
rect 474 642 476 644
rect 498 642 500 644
rect 504 642 506 644
rect 528 642 530 644
rect 534 642 536 644
rect 558 642 560 644
rect 564 642 566 644
rect 42 640 44 642
rect 72 640 74 642
rect 102 640 104 642
rect 132 640 134 642
rect 162 640 164 642
rect 436 640 438 642
rect 466 640 468 642
rect 496 640 498 642
rect 526 640 528 642
rect 556 640 558 642
rect 42 634 44 636
rect 72 634 74 636
rect 102 634 104 636
rect 132 634 134 636
rect 162 634 164 636
rect 436 634 438 636
rect 466 634 468 636
rect 496 634 498 636
rect 526 634 528 636
rect 556 634 558 636
rect 34 632 36 634
rect 40 632 42 634
rect 64 632 66 634
rect 70 632 72 634
rect 94 632 96 634
rect 100 632 102 634
rect 124 632 126 634
rect 130 632 132 634
rect 154 632 156 634
rect 160 632 162 634
rect 184 632 186 634
rect 414 632 416 634
rect 438 632 440 634
rect 444 632 446 634
rect 468 632 470 634
rect 474 632 476 634
rect 498 632 500 634
rect 504 632 506 634
rect 528 632 530 634
rect 534 632 536 634
rect 558 632 560 634
rect 564 632 566 634
rect 32 630 34 632
rect 62 630 64 632
rect 92 630 94 632
rect 122 630 124 632
rect 152 630 154 632
rect 182 630 184 632
rect 416 630 418 632
rect 446 630 448 632
rect 476 630 478 632
rect 506 630 508 632
rect 536 630 538 632
rect 566 630 568 632
rect 32 624 34 626
rect 62 624 64 626
rect 92 624 94 626
rect 122 624 124 626
rect 152 624 154 626
rect 182 624 184 626
rect 416 624 418 626
rect 446 624 448 626
rect 476 624 478 626
rect 506 624 508 626
rect 536 624 538 626
rect 566 624 568 626
rect 34 622 36 624
rect 40 622 42 624
rect 64 622 66 624
rect 70 622 72 624
rect 94 622 96 624
rect 100 622 102 624
rect 124 622 126 624
rect 130 622 132 624
rect 154 622 156 624
rect 160 622 162 624
rect 184 622 186 624
rect 414 622 416 624
rect 438 622 440 624
rect 444 622 446 624
rect 468 622 470 624
rect 474 622 476 624
rect 498 622 500 624
rect 504 622 506 624
rect 528 622 530 624
rect 534 622 536 624
rect 558 622 560 624
rect 564 622 566 624
rect 42 620 44 622
rect 72 620 74 622
rect 102 620 104 622
rect 132 620 134 622
rect 162 620 164 622
rect 436 620 438 622
rect 466 620 468 622
rect 496 620 498 622
rect 526 620 528 622
rect 556 620 558 622
rect 42 594 44 596
rect 72 594 74 596
rect 102 594 104 596
rect 132 594 134 596
rect 162 594 164 596
rect 436 594 438 596
rect 466 594 468 596
rect 496 594 498 596
rect 526 594 528 596
rect 556 594 558 596
rect 34 592 36 594
rect 40 592 42 594
rect 64 592 66 594
rect 70 592 72 594
rect 94 592 96 594
rect 100 592 102 594
rect 124 592 126 594
rect 130 592 132 594
rect 154 592 156 594
rect 160 592 162 594
rect 184 592 186 594
rect 414 592 416 594
rect 438 592 440 594
rect 444 592 446 594
rect 468 592 470 594
rect 474 592 476 594
rect 498 592 500 594
rect 504 592 506 594
rect 528 592 530 594
rect 534 592 536 594
rect 558 592 560 594
rect 564 592 566 594
rect 32 590 34 592
rect 62 590 64 592
rect 92 590 94 592
rect 122 590 124 592
rect 152 590 154 592
rect 182 590 184 592
rect 416 590 418 592
rect 446 590 448 592
rect 476 590 478 592
rect 506 590 508 592
rect 536 590 538 592
rect 566 590 568 592
rect 32 584 34 586
rect 62 584 64 586
rect 92 584 94 586
rect 506 584 508 586
rect 536 584 538 586
rect 566 584 568 586
rect 34 582 36 584
rect 40 582 42 584
rect 64 582 66 584
rect 70 582 72 584
rect 94 582 96 584
rect 100 582 102 584
rect 114 582 116 584
rect 130 582 132 584
rect 144 582 146 584
rect 160 582 162 584
rect 174 582 176 584
rect 424 582 426 584
rect 438 582 440 584
rect 454 582 456 584
rect 468 582 470 584
rect 484 582 486 584
rect 498 582 500 584
rect 504 582 506 584
rect 528 582 530 584
rect 534 582 536 584
rect 558 582 560 584
rect 564 582 566 584
rect 42 580 44 582
rect 72 580 74 582
rect 102 580 104 582
rect 112 580 114 582
rect 132 580 134 582
rect 142 580 144 582
rect 162 580 164 582
rect 172 580 174 582
rect 426 580 428 582
rect 436 580 438 582
rect 456 580 458 582
rect 466 580 468 582
rect 486 580 488 582
rect 496 580 498 582
rect 526 580 528 582
rect 556 580 558 582
rect 42 574 44 576
rect 72 574 74 576
rect 102 574 104 576
rect 112 574 114 576
rect 132 574 134 576
rect 142 574 144 576
rect 162 574 164 576
rect 172 574 174 576
rect 426 574 428 576
rect 436 574 438 576
rect 456 574 458 576
rect 466 574 468 576
rect 486 574 488 576
rect 496 574 498 576
rect 526 574 528 576
rect 556 574 558 576
rect 34 572 36 574
rect 40 572 42 574
rect 64 572 66 574
rect 70 572 72 574
rect 94 572 96 574
rect 100 572 102 574
rect 114 572 116 574
rect 130 572 132 574
rect 144 572 146 574
rect 160 572 162 574
rect 174 572 176 574
rect 424 572 426 574
rect 438 572 440 574
rect 454 572 456 574
rect 468 572 470 574
rect 484 572 486 574
rect 498 572 500 574
rect 504 572 506 574
rect 528 572 530 574
rect 534 572 536 574
rect 558 572 560 574
rect 564 572 566 574
rect 32 570 34 572
rect 62 570 64 572
rect 92 570 94 572
rect 506 570 508 572
rect 536 570 538 572
rect 566 570 568 572
rect 32 564 34 566
rect 62 564 64 566
rect 92 564 94 566
rect 122 564 124 566
rect 152 564 154 566
rect 182 564 184 566
rect 416 564 418 566
rect 446 564 448 566
rect 476 564 478 566
rect 506 564 508 566
rect 536 564 538 566
rect 566 564 568 566
rect 34 562 36 564
rect 40 562 42 564
rect 64 562 66 564
rect 70 562 72 564
rect 94 562 96 564
rect 100 562 102 564
rect 124 562 126 564
rect 130 562 132 564
rect 154 562 156 564
rect 160 562 162 564
rect 184 562 186 564
rect 414 562 416 564
rect 438 562 440 564
rect 444 562 446 564
rect 468 562 470 564
rect 474 562 476 564
rect 498 562 500 564
rect 504 562 506 564
rect 528 562 530 564
rect 534 562 536 564
rect 558 562 560 564
rect 564 562 566 564
rect 42 560 44 562
rect 72 560 74 562
rect 102 560 104 562
rect 132 560 134 562
rect 162 560 164 562
rect 436 560 438 562
rect 466 560 468 562
rect 496 560 498 562
rect 526 560 528 562
rect 556 560 558 562
rect 42 554 44 556
rect 72 554 74 556
rect 102 554 104 556
rect 132 554 134 556
rect 162 554 164 556
rect 436 554 438 556
rect 466 554 468 556
rect 496 554 498 556
rect 526 554 528 556
rect 556 554 558 556
rect 34 552 36 554
rect 40 552 42 554
rect 64 552 66 554
rect 70 552 72 554
rect 94 552 96 554
rect 100 552 102 554
rect 124 552 126 554
rect 130 552 132 554
rect 154 552 156 554
rect 160 552 162 554
rect 184 552 186 554
rect 414 552 416 554
rect 438 552 440 554
rect 444 552 446 554
rect 468 552 470 554
rect 474 552 476 554
rect 498 552 500 554
rect 504 552 506 554
rect 528 552 530 554
rect 534 552 536 554
rect 558 552 560 554
rect 564 552 566 554
rect 32 550 34 552
rect 62 550 64 552
rect 92 550 94 552
rect 122 550 124 552
rect 152 550 154 552
rect 182 550 184 552
rect 416 550 418 552
rect 446 550 448 552
rect 476 550 478 552
rect 506 550 508 552
rect 536 550 538 552
rect 566 550 568 552
rect 32 544 34 546
rect 62 544 64 546
rect 92 544 94 546
rect 122 544 124 546
rect 152 544 154 546
rect 182 544 184 546
rect 416 544 418 546
rect 446 544 448 546
rect 476 544 478 546
rect 506 544 508 546
rect 536 544 538 546
rect 566 544 568 546
rect 34 542 36 544
rect 40 542 42 544
rect 64 542 66 544
rect 70 542 72 544
rect 94 542 96 544
rect 100 542 102 544
rect 124 542 126 544
rect 130 542 132 544
rect 154 542 156 544
rect 160 542 162 544
rect 184 542 186 544
rect 414 542 416 544
rect 438 542 440 544
rect 444 542 446 544
rect 468 542 470 544
rect 474 542 476 544
rect 498 542 500 544
rect 504 542 506 544
rect 528 542 530 544
rect 534 542 536 544
rect 558 542 560 544
rect 564 542 566 544
rect 42 540 44 542
rect 72 540 74 542
rect 102 540 104 542
rect 132 540 134 542
rect 162 540 164 542
rect 436 540 438 542
rect 466 540 468 542
rect 496 540 498 542
rect 526 540 528 542
rect 556 540 558 542
rect 42 534 44 536
rect 72 534 74 536
rect 102 534 104 536
rect 132 534 134 536
rect 162 534 164 536
rect 436 534 438 536
rect 466 534 468 536
rect 496 534 498 536
rect 526 534 528 536
rect 556 534 558 536
rect 34 532 36 534
rect 40 532 42 534
rect 64 532 66 534
rect 70 532 72 534
rect 94 532 96 534
rect 100 532 102 534
rect 124 532 126 534
rect 130 532 132 534
rect 154 532 156 534
rect 160 532 162 534
rect 184 532 186 534
rect 414 532 416 534
rect 438 532 440 534
rect 444 532 446 534
rect 468 532 470 534
rect 474 532 476 534
rect 498 532 500 534
rect 504 532 506 534
rect 528 532 530 534
rect 534 532 536 534
rect 558 532 560 534
rect 564 532 566 534
rect 32 530 34 532
rect 62 530 64 532
rect 92 530 94 532
rect 122 530 124 532
rect 152 530 154 532
rect 182 530 184 532
rect 416 530 418 532
rect 446 530 448 532
rect 476 530 478 532
rect 506 530 508 532
rect 536 530 538 532
rect 566 530 568 532
rect 38 461 40 463
rect 48 461 50 463
rect 58 461 60 463
rect 78 461 80 463
rect 88 461 90 463
rect 108 461 110 463
rect 118 461 120 463
rect 138 461 140 463
rect 148 461 150 463
rect 168 461 170 463
rect 178 461 180 463
rect 198 461 200 463
rect 208 461 210 463
rect 228 461 230 463
rect 238 461 240 463
rect 258 461 260 463
rect 268 461 270 463
rect 288 461 290 463
rect 298 461 300 463
rect 318 461 320 463
rect 328 461 330 463
rect 348 461 350 463
rect 358 461 360 463
rect 378 461 380 463
rect 388 461 390 463
rect 408 461 410 463
rect 418 461 420 463
rect 438 461 440 463
rect 448 461 450 463
rect 468 461 470 463
rect 478 461 480 463
rect 498 461 500 463
rect 508 461 510 463
rect 528 461 530 463
rect 538 461 540 463
rect 558 461 560 463
rect 40 459 42 461
rect 46 459 48 461
rect 60 459 62 461
rect 76 459 78 461
rect 90 459 92 461
rect 106 459 108 461
rect 120 459 122 461
rect 136 459 138 461
rect 150 459 152 461
rect 166 459 168 461
rect 180 459 182 461
rect 196 459 198 461
rect 210 459 212 461
rect 226 459 228 461
rect 240 459 242 461
rect 256 459 258 461
rect 270 459 272 461
rect 286 459 288 461
rect 300 459 302 461
rect 316 459 318 461
rect 330 459 332 461
rect 346 459 348 461
rect 360 459 362 461
rect 376 459 378 461
rect 390 459 392 461
rect 406 459 408 461
rect 420 459 422 461
rect 436 459 438 461
rect 450 459 452 461
rect 466 459 468 461
rect 480 459 482 461
rect 496 459 498 461
rect 510 459 512 461
rect 526 459 528 461
rect 540 459 542 461
rect 556 459 558 461
rect 68 451 70 453
rect 98 451 100 453
rect 128 451 130 453
rect 158 451 160 453
rect 188 451 190 453
rect 218 451 220 453
rect 248 451 250 453
rect 278 451 280 453
rect 308 451 310 453
rect 338 451 340 453
rect 368 451 370 453
rect 398 451 400 453
rect 428 451 430 453
rect 458 451 460 453
rect 488 451 490 453
rect 518 451 520 453
rect 548 451 550 453
rect 60 449 62 451
rect 66 449 68 451
rect 90 449 92 451
rect 96 449 98 451
rect 120 449 122 451
rect 126 449 128 451
rect 150 449 152 451
rect 156 449 158 451
rect 180 449 182 451
rect 186 449 188 451
rect 210 449 212 451
rect 216 449 218 451
rect 240 449 242 451
rect 246 449 248 451
rect 270 449 272 451
rect 276 449 278 451
rect 300 449 302 451
rect 306 449 308 451
rect 330 449 332 451
rect 336 449 338 451
rect 360 449 362 451
rect 366 449 368 451
rect 390 449 392 451
rect 396 449 398 451
rect 420 449 422 451
rect 426 449 428 451
rect 450 449 452 451
rect 456 449 458 451
rect 480 449 482 451
rect 486 449 488 451
rect 510 449 512 451
rect 516 449 518 451
rect 540 449 542 451
rect 546 449 548 451
rect 58 447 60 449
rect 88 447 90 449
rect 118 447 120 449
rect 148 447 150 449
rect 178 447 180 449
rect 208 447 210 449
rect 238 447 240 449
rect 268 447 270 449
rect 298 447 300 449
rect 328 447 330 449
rect 358 447 360 449
rect 388 447 390 449
rect 418 447 420 449
rect 448 447 450 449
rect 478 447 480 449
rect 508 447 510 449
rect 538 447 540 449
rect 58 441 60 443
rect 88 441 90 443
rect 118 441 120 443
rect 148 441 150 443
rect 178 441 180 443
rect 208 441 210 443
rect 238 441 240 443
rect 268 441 270 443
rect 298 441 300 443
rect 328 441 330 443
rect 358 441 360 443
rect 388 441 390 443
rect 418 441 420 443
rect 448 441 450 443
rect 478 441 480 443
rect 508 441 510 443
rect 538 441 540 443
rect 60 439 62 441
rect 66 439 68 441
rect 90 439 92 441
rect 96 439 98 441
rect 120 439 122 441
rect 126 439 128 441
rect 150 439 152 441
rect 156 439 158 441
rect 180 439 182 441
rect 186 439 188 441
rect 210 439 212 441
rect 216 439 218 441
rect 240 439 242 441
rect 246 439 248 441
rect 270 439 272 441
rect 276 439 278 441
rect 300 439 302 441
rect 306 439 308 441
rect 330 439 332 441
rect 336 439 338 441
rect 360 439 362 441
rect 366 439 368 441
rect 390 439 392 441
rect 396 439 398 441
rect 420 439 422 441
rect 426 439 428 441
rect 450 439 452 441
rect 456 439 458 441
rect 480 439 482 441
rect 486 439 488 441
rect 510 439 512 441
rect 516 439 518 441
rect 540 439 542 441
rect 546 439 548 441
rect 68 437 70 439
rect 98 437 100 439
rect 128 437 130 439
rect 158 437 160 439
rect 188 437 190 439
rect 218 437 220 439
rect 248 437 250 439
rect 278 437 280 439
rect 308 437 310 439
rect 338 437 340 439
rect 368 437 370 439
rect 398 437 400 439
rect 428 437 430 439
rect 458 437 460 439
rect 488 437 490 439
rect 518 437 520 439
rect 548 437 550 439
rect 68 431 70 433
rect 98 431 100 433
rect 128 431 130 433
rect 158 431 160 433
rect 188 431 190 433
rect 218 431 220 433
rect 248 431 250 433
rect 278 431 280 433
rect 308 431 310 433
rect 338 431 340 433
rect 368 431 370 433
rect 398 431 400 433
rect 428 431 430 433
rect 458 431 460 433
rect 488 431 490 433
rect 518 431 520 433
rect 548 431 550 433
rect 60 429 62 431
rect 66 429 68 431
rect 90 429 92 431
rect 96 429 98 431
rect 120 429 122 431
rect 126 429 128 431
rect 150 429 152 431
rect 156 429 158 431
rect 180 429 182 431
rect 186 429 188 431
rect 210 429 212 431
rect 216 429 218 431
rect 240 429 242 431
rect 246 429 248 431
rect 270 429 272 431
rect 276 429 278 431
rect 300 429 302 431
rect 306 429 308 431
rect 330 429 332 431
rect 336 429 338 431
rect 360 429 362 431
rect 366 429 368 431
rect 390 429 392 431
rect 396 429 398 431
rect 420 429 422 431
rect 426 429 428 431
rect 450 429 452 431
rect 456 429 458 431
rect 480 429 482 431
rect 486 429 488 431
rect 510 429 512 431
rect 516 429 518 431
rect 540 429 542 431
rect 546 429 548 431
rect 58 427 60 429
rect 88 427 90 429
rect 118 427 120 429
rect 148 427 150 429
rect 178 427 180 429
rect 208 427 210 429
rect 238 427 240 429
rect 268 427 270 429
rect 298 427 300 429
rect 328 427 330 429
rect 358 427 360 429
rect 388 427 390 429
rect 418 427 420 429
rect 448 427 450 429
rect 478 427 480 429
rect 508 427 510 429
rect 538 427 540 429
rect 58 421 60 423
rect 88 421 90 423
rect 118 421 120 423
rect 148 421 150 423
rect 178 421 180 423
rect 208 421 210 423
rect 238 421 240 423
rect 268 421 270 423
rect 298 421 300 423
rect 328 421 330 423
rect 358 421 360 423
rect 388 421 390 423
rect 418 421 420 423
rect 448 421 450 423
rect 478 421 480 423
rect 508 421 510 423
rect 538 421 540 423
rect 60 419 62 421
rect 66 419 68 421
rect 90 419 92 421
rect 96 419 98 421
rect 120 419 122 421
rect 126 419 128 421
rect 150 419 152 421
rect 156 419 158 421
rect 180 419 182 421
rect 186 419 188 421
rect 210 419 212 421
rect 216 419 218 421
rect 240 419 242 421
rect 246 419 248 421
rect 270 419 272 421
rect 276 419 278 421
rect 300 419 302 421
rect 306 419 308 421
rect 330 419 332 421
rect 336 419 338 421
rect 360 419 362 421
rect 366 419 368 421
rect 390 419 392 421
rect 396 419 398 421
rect 420 419 422 421
rect 426 419 428 421
rect 450 419 452 421
rect 456 419 458 421
rect 480 419 482 421
rect 486 419 488 421
rect 510 419 512 421
rect 516 419 518 421
rect 540 419 542 421
rect 546 419 548 421
rect 68 417 70 419
rect 98 417 100 419
rect 128 417 130 419
rect 158 417 160 419
rect 188 417 190 419
rect 218 417 220 419
rect 248 417 250 419
rect 278 417 280 419
rect 308 417 310 419
rect 338 417 340 419
rect 368 417 370 419
rect 398 417 400 419
rect 428 417 430 419
rect 458 417 460 419
rect 488 417 490 419
rect 518 417 520 419
rect 548 417 550 419
rect 68 411 70 413
rect 98 411 100 413
rect 128 411 130 413
rect 158 411 160 413
rect 188 411 190 413
rect 218 411 220 413
rect 248 411 250 413
rect 278 411 280 413
rect 308 411 310 413
rect 338 411 340 413
rect 368 411 370 413
rect 398 411 400 413
rect 428 411 430 413
rect 458 411 460 413
rect 488 411 490 413
rect 518 411 520 413
rect 548 411 550 413
rect 60 409 62 411
rect 66 409 68 411
rect 90 409 92 411
rect 96 409 98 411
rect 120 409 122 411
rect 126 409 128 411
rect 150 409 152 411
rect 156 409 158 411
rect 180 409 182 411
rect 186 409 188 411
rect 210 409 212 411
rect 216 409 218 411
rect 240 409 242 411
rect 246 409 248 411
rect 270 409 272 411
rect 276 409 278 411
rect 300 409 302 411
rect 306 409 308 411
rect 330 409 332 411
rect 336 409 338 411
rect 360 409 362 411
rect 366 409 368 411
rect 390 409 392 411
rect 396 409 398 411
rect 420 409 422 411
rect 426 409 428 411
rect 450 409 452 411
rect 456 409 458 411
rect 480 409 482 411
rect 486 409 488 411
rect 510 409 512 411
rect 516 409 518 411
rect 540 409 542 411
rect 546 409 548 411
rect 58 407 60 409
rect 88 407 90 409
rect 118 407 120 409
rect 148 407 150 409
rect 178 407 180 409
rect 208 407 210 409
rect 238 407 240 409
rect 268 407 270 409
rect 298 407 300 409
rect 328 407 330 409
rect 358 407 360 409
rect 388 407 390 409
rect 418 407 420 409
rect 448 407 450 409
rect 478 407 480 409
rect 508 407 510 409
rect 538 407 540 409
rect 58 401 60 403
rect 88 401 90 403
rect 118 401 120 403
rect 148 401 150 403
rect 178 401 180 403
rect 208 401 210 403
rect 238 401 240 403
rect 268 401 270 403
rect 298 401 300 403
rect 328 401 330 403
rect 358 401 360 403
rect 388 401 390 403
rect 418 401 420 403
rect 448 401 450 403
rect 478 401 480 403
rect 508 401 510 403
rect 538 401 540 403
rect 60 399 62 401
rect 66 399 68 401
rect 90 399 92 401
rect 96 399 98 401
rect 120 399 122 401
rect 126 399 128 401
rect 150 399 152 401
rect 156 399 158 401
rect 180 399 182 401
rect 186 399 188 401
rect 210 399 212 401
rect 216 399 218 401
rect 240 399 242 401
rect 246 399 248 401
rect 270 399 272 401
rect 276 399 278 401
rect 300 399 302 401
rect 306 399 308 401
rect 330 399 332 401
rect 336 399 338 401
rect 360 399 362 401
rect 366 399 368 401
rect 390 399 392 401
rect 396 399 398 401
rect 420 399 422 401
rect 426 399 428 401
rect 450 399 452 401
rect 456 399 458 401
rect 480 399 482 401
rect 486 399 488 401
rect 510 399 512 401
rect 516 399 518 401
rect 540 399 542 401
rect 546 399 548 401
rect 68 397 70 399
rect 98 397 100 399
rect 128 397 130 399
rect 158 397 160 399
rect 188 397 190 399
rect 218 397 220 399
rect 248 397 250 399
rect 278 397 280 399
rect 308 397 310 399
rect 338 397 340 399
rect 368 397 370 399
rect 398 397 400 399
rect 428 397 430 399
rect 458 397 460 399
rect 488 397 490 399
rect 518 397 520 399
rect 548 397 550 399
rect 98 391 100 393
rect 518 391 520 393
rect 548 391 550 393
rect 96 389 98 391
rect 516 389 518 391
rect 540 389 542 391
rect 546 389 548 391
rect 538 387 540 389
rect 538 381 540 383
rect 96 379 98 381
rect 516 379 518 381
rect 540 379 542 381
rect 546 379 548 381
rect 98 377 100 379
rect 518 377 520 379
rect 548 377 550 379
rect 68 371 70 373
rect 98 371 100 373
rect 128 371 130 373
rect 158 371 160 373
rect 188 371 190 373
rect 218 371 220 373
rect 248 371 250 373
rect 278 371 280 373
rect 308 371 310 373
rect 338 371 340 373
rect 368 371 370 373
rect 398 371 400 373
rect 428 371 430 373
rect 458 371 460 373
rect 488 371 490 373
rect 518 371 520 373
rect 548 371 550 373
rect 60 369 62 371
rect 66 369 68 371
rect 90 369 92 371
rect 96 369 98 371
rect 120 369 122 371
rect 126 369 128 371
rect 150 369 152 371
rect 156 369 158 371
rect 180 369 182 371
rect 186 369 188 371
rect 210 369 212 371
rect 216 369 218 371
rect 240 369 242 371
rect 246 369 248 371
rect 270 369 272 371
rect 276 369 278 371
rect 300 369 302 371
rect 306 369 308 371
rect 330 369 332 371
rect 336 369 338 371
rect 360 369 362 371
rect 366 369 368 371
rect 390 369 392 371
rect 396 369 398 371
rect 420 369 422 371
rect 426 369 428 371
rect 450 369 452 371
rect 456 369 458 371
rect 480 369 482 371
rect 486 369 488 371
rect 510 369 512 371
rect 516 369 518 371
rect 540 369 542 371
rect 546 369 548 371
rect 58 367 60 369
rect 88 367 90 369
rect 118 367 120 369
rect 148 367 150 369
rect 178 367 180 369
rect 208 367 210 369
rect 238 367 240 369
rect 268 367 270 369
rect 298 367 300 369
rect 328 367 330 369
rect 358 367 360 369
rect 388 367 390 369
rect 418 367 420 369
rect 448 367 450 369
rect 478 367 480 369
rect 508 367 510 369
rect 538 367 540 369
rect 58 361 60 363
rect 88 361 90 363
rect 118 361 120 363
rect 148 361 150 363
rect 178 361 180 363
rect 208 361 210 363
rect 238 361 240 363
rect 268 361 270 363
rect 298 361 300 363
rect 328 361 330 363
rect 358 361 360 363
rect 388 361 390 363
rect 418 361 420 363
rect 448 361 450 363
rect 478 361 480 363
rect 508 361 510 363
rect 538 361 540 363
rect 60 359 62 361
rect 66 359 68 361
rect 90 359 92 361
rect 96 359 98 361
rect 120 359 122 361
rect 126 359 128 361
rect 150 359 152 361
rect 156 359 158 361
rect 180 359 182 361
rect 186 359 188 361
rect 210 359 212 361
rect 216 359 218 361
rect 240 359 242 361
rect 246 359 248 361
rect 270 359 272 361
rect 276 359 278 361
rect 300 359 302 361
rect 306 359 308 361
rect 330 359 332 361
rect 336 359 338 361
rect 360 359 362 361
rect 366 359 368 361
rect 390 359 392 361
rect 396 359 398 361
rect 420 359 422 361
rect 426 359 428 361
rect 450 359 452 361
rect 456 359 458 361
rect 480 359 482 361
rect 486 359 488 361
rect 510 359 512 361
rect 516 359 518 361
rect 540 359 542 361
rect 546 359 548 361
rect 68 357 70 359
rect 98 357 100 359
rect 128 357 130 359
rect 158 357 160 359
rect 188 357 190 359
rect 218 357 220 359
rect 248 357 250 359
rect 278 357 280 359
rect 308 357 310 359
rect 338 357 340 359
rect 368 357 370 359
rect 398 357 400 359
rect 428 357 430 359
rect 458 357 460 359
rect 488 357 490 359
rect 518 357 520 359
rect 548 357 550 359
rect 68 351 70 353
rect 98 351 100 353
rect 128 351 130 353
rect 158 351 160 353
rect 188 351 190 353
rect 218 351 220 353
rect 248 351 250 353
rect 278 351 280 353
rect 308 351 310 353
rect 338 351 340 353
rect 368 351 370 353
rect 398 351 400 353
rect 428 351 430 353
rect 458 351 460 353
rect 488 351 490 353
rect 518 351 520 353
rect 548 351 550 353
rect 60 349 62 351
rect 66 349 68 351
rect 90 349 92 351
rect 96 349 98 351
rect 120 349 122 351
rect 126 349 128 351
rect 150 349 152 351
rect 156 349 158 351
rect 180 349 182 351
rect 186 349 188 351
rect 210 349 212 351
rect 216 349 218 351
rect 240 349 242 351
rect 246 349 248 351
rect 270 349 272 351
rect 276 349 278 351
rect 300 349 302 351
rect 306 349 308 351
rect 330 349 332 351
rect 336 349 338 351
rect 360 349 362 351
rect 366 349 368 351
rect 390 349 392 351
rect 396 349 398 351
rect 420 349 422 351
rect 426 349 428 351
rect 450 349 452 351
rect 456 349 458 351
rect 480 349 482 351
rect 486 349 488 351
rect 510 349 512 351
rect 516 349 518 351
rect 540 349 542 351
rect 546 349 548 351
rect 58 347 60 349
rect 88 347 90 349
rect 118 347 120 349
rect 148 347 150 349
rect 178 347 180 349
rect 208 347 210 349
rect 238 347 240 349
rect 268 347 270 349
rect 298 347 300 349
rect 328 347 330 349
rect 358 347 360 349
rect 388 347 390 349
rect 418 347 420 349
rect 448 347 450 349
rect 478 347 480 349
rect 508 347 510 349
rect 538 347 540 349
rect 58 341 60 343
rect 88 341 90 343
rect 118 341 120 343
rect 148 341 150 343
rect 178 341 180 343
rect 208 341 210 343
rect 238 341 240 343
rect 268 341 270 343
rect 298 341 300 343
rect 328 341 330 343
rect 358 341 360 343
rect 388 341 390 343
rect 418 341 420 343
rect 448 341 450 343
rect 478 341 480 343
rect 508 341 510 343
rect 538 341 540 343
rect 60 339 62 341
rect 66 339 68 341
rect 90 339 92 341
rect 96 339 98 341
rect 120 339 122 341
rect 126 339 128 341
rect 150 339 152 341
rect 156 339 158 341
rect 180 339 182 341
rect 186 339 188 341
rect 210 339 212 341
rect 216 339 218 341
rect 240 339 242 341
rect 246 339 248 341
rect 270 339 272 341
rect 276 339 278 341
rect 300 339 302 341
rect 306 339 308 341
rect 330 339 332 341
rect 336 339 338 341
rect 360 339 362 341
rect 366 339 368 341
rect 390 339 392 341
rect 396 339 398 341
rect 420 339 422 341
rect 426 339 428 341
rect 450 339 452 341
rect 456 339 458 341
rect 480 339 482 341
rect 486 339 488 341
rect 510 339 512 341
rect 516 339 518 341
rect 540 339 542 341
rect 546 339 548 341
rect 68 337 70 339
rect 98 337 100 339
rect 128 337 130 339
rect 158 337 160 339
rect 188 337 190 339
rect 218 337 220 339
rect 248 337 250 339
rect 278 337 280 339
rect 308 337 310 339
rect 338 337 340 339
rect 368 337 370 339
rect 398 337 400 339
rect 428 337 430 339
rect 458 337 460 339
rect 488 337 490 339
rect 518 337 520 339
rect 548 337 550 339
rect 68 331 70 333
rect 98 331 100 333
rect 128 331 130 333
rect 158 331 160 333
rect 188 331 190 333
rect 218 331 220 333
rect 248 331 250 333
rect 278 331 280 333
rect 308 331 310 333
rect 338 331 340 333
rect 368 331 370 333
rect 398 331 400 333
rect 428 331 430 333
rect 458 331 460 333
rect 488 331 490 333
rect 518 331 520 333
rect 548 331 550 333
rect 60 329 62 331
rect 66 329 68 331
rect 90 329 92 331
rect 96 329 98 331
rect 120 329 122 331
rect 126 329 128 331
rect 150 329 152 331
rect 156 329 158 331
rect 180 329 182 331
rect 186 329 188 331
rect 210 329 212 331
rect 216 329 218 331
rect 240 329 242 331
rect 246 329 248 331
rect 270 329 272 331
rect 276 329 278 331
rect 300 329 302 331
rect 306 329 308 331
rect 330 329 332 331
rect 336 329 338 331
rect 360 329 362 331
rect 366 329 368 331
rect 390 329 392 331
rect 396 329 398 331
rect 420 329 422 331
rect 426 329 428 331
rect 450 329 452 331
rect 456 329 458 331
rect 480 329 482 331
rect 486 329 488 331
rect 510 329 512 331
rect 516 329 518 331
rect 540 329 542 331
rect 546 329 548 331
rect 58 327 60 329
rect 88 327 90 329
rect 118 327 120 329
rect 148 327 150 329
rect 178 327 180 329
rect 208 327 210 329
rect 238 327 240 329
rect 268 327 270 329
rect 298 327 300 329
rect 328 327 330 329
rect 358 327 360 329
rect 388 327 390 329
rect 418 327 420 329
rect 448 327 450 329
rect 478 327 480 329
rect 508 327 510 329
rect 538 327 540 329
rect 58 321 60 323
rect 88 321 90 323
rect 118 321 120 323
rect 148 321 150 323
rect 178 321 180 323
rect 208 321 210 323
rect 238 321 240 323
rect 268 321 270 323
rect 298 321 300 323
rect 328 321 330 323
rect 358 321 360 323
rect 388 321 390 323
rect 418 321 420 323
rect 448 321 450 323
rect 478 321 480 323
rect 508 321 510 323
rect 538 321 540 323
rect 60 319 62 321
rect 66 319 68 321
rect 90 319 92 321
rect 96 319 98 321
rect 120 319 122 321
rect 126 319 128 321
rect 150 319 152 321
rect 156 319 158 321
rect 180 319 182 321
rect 186 319 188 321
rect 210 319 212 321
rect 216 319 218 321
rect 240 319 242 321
rect 246 319 248 321
rect 270 319 272 321
rect 276 319 278 321
rect 300 319 302 321
rect 306 319 308 321
rect 330 319 332 321
rect 336 319 338 321
rect 360 319 362 321
rect 366 319 368 321
rect 390 319 392 321
rect 396 319 398 321
rect 420 319 422 321
rect 426 319 428 321
rect 450 319 452 321
rect 456 319 458 321
rect 480 319 482 321
rect 486 319 488 321
rect 510 319 512 321
rect 516 319 518 321
rect 540 319 542 321
rect 546 319 548 321
rect 68 317 70 319
rect 98 317 100 319
rect 128 317 130 319
rect 158 317 160 319
rect 188 317 190 319
rect 218 317 220 319
rect 248 317 250 319
rect 278 317 280 319
rect 308 317 310 319
rect 338 317 340 319
rect 368 317 370 319
rect 398 317 400 319
rect 428 317 430 319
rect 458 317 460 319
rect 488 317 490 319
rect 518 317 520 319
rect 548 317 550 319
rect 68 311 70 313
rect 518 311 520 313
rect 548 311 550 313
rect 60 309 62 311
rect 66 309 68 311
rect 510 309 512 311
rect 516 309 518 311
rect 540 309 542 311
rect 546 309 548 311
rect 58 307 60 309
rect 508 307 510 309
rect 538 307 540 309
rect 58 301 60 303
rect 508 301 510 303
rect 538 301 540 303
rect 60 299 62 301
rect 66 299 68 301
rect 510 299 512 301
rect 516 299 518 301
rect 540 299 542 301
rect 546 299 548 301
rect 68 297 70 299
rect 518 297 520 299
rect 548 297 550 299
rect 68 291 70 293
rect 98 291 100 293
rect 128 291 130 293
rect 158 291 160 293
rect 188 291 190 293
rect 218 291 220 293
rect 248 291 250 293
rect 278 291 280 293
rect 308 291 310 293
rect 338 291 340 293
rect 368 291 370 293
rect 398 291 400 293
rect 428 291 430 293
rect 458 291 460 293
rect 488 291 490 293
rect 518 291 520 293
rect 548 291 550 293
rect 60 289 62 291
rect 66 289 68 291
rect 90 289 92 291
rect 96 289 98 291
rect 120 289 122 291
rect 126 289 128 291
rect 150 289 152 291
rect 156 289 158 291
rect 180 289 182 291
rect 186 289 188 291
rect 210 289 212 291
rect 216 289 218 291
rect 240 289 242 291
rect 246 289 248 291
rect 270 289 272 291
rect 276 289 278 291
rect 300 289 302 291
rect 306 289 308 291
rect 330 289 332 291
rect 336 289 338 291
rect 360 289 362 291
rect 366 289 368 291
rect 390 289 392 291
rect 396 289 398 291
rect 420 289 422 291
rect 426 289 428 291
rect 450 289 452 291
rect 456 289 458 291
rect 480 289 482 291
rect 486 289 488 291
rect 510 289 512 291
rect 516 289 518 291
rect 540 289 542 291
rect 546 289 548 291
rect 58 287 60 289
rect 88 287 90 289
rect 118 287 120 289
rect 148 287 150 289
rect 178 287 180 289
rect 208 287 210 289
rect 238 287 240 289
rect 268 287 270 289
rect 298 287 300 289
rect 328 287 330 289
rect 358 287 360 289
rect 388 287 390 289
rect 418 287 420 289
rect 448 287 450 289
rect 478 287 480 289
rect 508 287 510 289
rect 538 287 540 289
rect 58 281 60 283
rect 88 281 90 283
rect 118 281 120 283
rect 148 281 150 283
rect 178 281 180 283
rect 208 281 210 283
rect 238 281 240 283
rect 268 281 270 283
rect 298 281 300 283
rect 328 281 330 283
rect 358 281 360 283
rect 388 281 390 283
rect 418 281 420 283
rect 448 281 450 283
rect 478 281 480 283
rect 508 281 510 283
rect 538 281 540 283
rect 60 279 62 281
rect 66 279 68 281
rect 90 279 92 281
rect 96 279 98 281
rect 120 279 122 281
rect 126 279 128 281
rect 150 279 152 281
rect 156 279 158 281
rect 180 279 182 281
rect 186 279 188 281
rect 210 279 212 281
rect 216 279 218 281
rect 240 279 242 281
rect 246 279 248 281
rect 270 279 272 281
rect 276 279 278 281
rect 300 279 302 281
rect 306 279 308 281
rect 330 279 332 281
rect 336 279 338 281
rect 360 279 362 281
rect 366 279 368 281
rect 390 279 392 281
rect 396 279 398 281
rect 420 279 422 281
rect 426 279 428 281
rect 450 279 452 281
rect 456 279 458 281
rect 480 279 482 281
rect 486 279 488 281
rect 510 279 512 281
rect 516 279 518 281
rect 540 279 542 281
rect 546 279 548 281
rect 68 277 70 279
rect 98 277 100 279
rect 128 277 130 279
rect 158 277 160 279
rect 188 277 190 279
rect 218 277 220 279
rect 248 277 250 279
rect 278 277 280 279
rect 308 277 310 279
rect 338 277 340 279
rect 368 277 370 279
rect 398 277 400 279
rect 428 277 430 279
rect 458 277 460 279
rect 488 277 490 279
rect 518 277 520 279
rect 548 277 550 279
rect 68 271 70 273
rect 98 271 100 273
rect 128 271 130 273
rect 158 271 160 273
rect 188 271 190 273
rect 218 271 220 273
rect 248 271 250 273
rect 278 271 280 273
rect 308 271 310 273
rect 338 271 340 273
rect 368 271 370 273
rect 398 271 400 273
rect 428 271 430 273
rect 458 271 460 273
rect 488 271 490 273
rect 518 271 520 273
rect 548 271 550 273
rect 60 269 62 271
rect 66 269 68 271
rect 90 269 92 271
rect 96 269 98 271
rect 120 269 122 271
rect 126 269 128 271
rect 150 269 152 271
rect 156 269 158 271
rect 180 269 182 271
rect 186 269 188 271
rect 210 269 212 271
rect 216 269 218 271
rect 240 269 242 271
rect 246 269 248 271
rect 270 269 272 271
rect 276 269 278 271
rect 300 269 302 271
rect 306 269 308 271
rect 330 269 332 271
rect 336 269 338 271
rect 360 269 362 271
rect 366 269 368 271
rect 390 269 392 271
rect 396 269 398 271
rect 420 269 422 271
rect 426 269 428 271
rect 450 269 452 271
rect 456 269 458 271
rect 480 269 482 271
rect 486 269 488 271
rect 510 269 512 271
rect 516 269 518 271
rect 540 269 542 271
rect 546 269 548 271
rect 58 267 60 269
rect 88 267 90 269
rect 118 267 120 269
rect 148 267 150 269
rect 178 267 180 269
rect 208 267 210 269
rect 238 267 240 269
rect 268 267 270 269
rect 298 267 300 269
rect 328 267 330 269
rect 358 267 360 269
rect 388 267 390 269
rect 418 267 420 269
rect 448 267 450 269
rect 478 267 480 269
rect 508 267 510 269
rect 538 267 540 269
rect 58 261 60 263
rect 88 261 90 263
rect 118 261 120 263
rect 148 261 150 263
rect 178 261 180 263
rect 208 261 210 263
rect 238 261 240 263
rect 268 261 270 263
rect 298 261 300 263
rect 328 261 330 263
rect 358 261 360 263
rect 388 261 390 263
rect 418 261 420 263
rect 448 261 450 263
rect 478 261 480 263
rect 508 261 510 263
rect 538 261 540 263
rect 60 259 62 261
rect 66 259 68 261
rect 90 259 92 261
rect 96 259 98 261
rect 120 259 122 261
rect 126 259 128 261
rect 150 259 152 261
rect 156 259 158 261
rect 180 259 182 261
rect 186 259 188 261
rect 210 259 212 261
rect 216 259 218 261
rect 240 259 242 261
rect 246 259 248 261
rect 270 259 272 261
rect 276 259 278 261
rect 300 259 302 261
rect 306 259 308 261
rect 330 259 332 261
rect 336 259 338 261
rect 360 259 362 261
rect 366 259 368 261
rect 390 259 392 261
rect 396 259 398 261
rect 420 259 422 261
rect 426 259 428 261
rect 450 259 452 261
rect 456 259 458 261
rect 480 259 482 261
rect 486 259 488 261
rect 510 259 512 261
rect 516 259 518 261
rect 540 259 542 261
rect 546 259 548 261
rect 68 257 70 259
rect 98 257 100 259
rect 128 257 130 259
rect 158 257 160 259
rect 188 257 190 259
rect 218 257 220 259
rect 248 257 250 259
rect 278 257 280 259
rect 308 257 310 259
rect 338 257 340 259
rect 368 257 370 259
rect 398 257 400 259
rect 428 257 430 259
rect 458 257 460 259
rect 488 257 490 259
rect 518 257 520 259
rect 548 257 550 259
rect 68 251 70 253
rect 98 251 100 253
rect 128 251 130 253
rect 158 251 160 253
rect 188 251 190 253
rect 218 251 220 253
rect 248 251 250 253
rect 278 251 280 253
rect 308 251 310 253
rect 338 251 340 253
rect 368 251 370 253
rect 398 251 400 253
rect 428 251 430 253
rect 458 251 460 253
rect 488 251 490 253
rect 518 251 520 253
rect 548 251 550 253
rect 60 249 62 251
rect 66 249 68 251
rect 90 249 92 251
rect 96 249 98 251
rect 120 249 122 251
rect 126 249 128 251
rect 150 249 152 251
rect 156 249 158 251
rect 180 249 182 251
rect 186 249 188 251
rect 210 249 212 251
rect 216 249 218 251
rect 240 249 242 251
rect 246 249 248 251
rect 270 249 272 251
rect 276 249 278 251
rect 300 249 302 251
rect 306 249 308 251
rect 330 249 332 251
rect 336 249 338 251
rect 360 249 362 251
rect 366 249 368 251
rect 390 249 392 251
rect 396 249 398 251
rect 420 249 422 251
rect 426 249 428 251
rect 450 249 452 251
rect 456 249 458 251
rect 480 249 482 251
rect 486 249 488 251
rect 510 249 512 251
rect 516 249 518 251
rect 540 249 542 251
rect 546 249 548 251
rect 58 247 60 249
rect 88 247 90 249
rect 118 247 120 249
rect 148 247 150 249
rect 178 247 180 249
rect 208 247 210 249
rect 238 247 240 249
rect 268 247 270 249
rect 298 247 300 249
rect 328 247 330 249
rect 358 247 360 249
rect 388 247 390 249
rect 418 247 420 249
rect 448 247 450 249
rect 478 247 480 249
rect 508 247 510 249
rect 538 247 540 249
rect 58 241 60 243
rect 88 241 90 243
rect 508 241 510 243
rect 538 241 540 243
rect 60 239 62 241
rect 86 239 88 241
rect 506 239 508 241
rect 540 239 542 241
rect 546 239 548 241
rect 548 237 550 239
rect 548 231 550 233
rect 60 229 62 231
rect 86 229 88 231
rect 506 229 508 231
rect 540 229 542 231
rect 546 229 548 231
rect 58 227 60 229
rect 88 227 90 229
rect 508 227 510 229
rect 538 227 540 229
rect 58 221 60 223
rect 88 221 90 223
rect 118 221 120 223
rect 148 221 150 223
rect 178 221 180 223
rect 208 221 210 223
rect 238 221 240 223
rect 268 221 270 223
rect 298 221 300 223
rect 328 221 330 223
rect 358 221 360 223
rect 388 221 390 223
rect 418 221 420 223
rect 448 221 450 223
rect 478 221 480 223
rect 508 221 510 223
rect 538 221 540 223
rect 60 219 62 221
rect 66 219 68 221
rect 90 219 92 221
rect 96 219 98 221
rect 120 219 122 221
rect 126 219 128 221
rect 150 219 152 221
rect 156 219 158 221
rect 180 219 182 221
rect 186 219 188 221
rect 210 219 212 221
rect 216 219 218 221
rect 240 219 242 221
rect 246 219 248 221
rect 270 219 272 221
rect 276 219 278 221
rect 300 219 302 221
rect 306 219 308 221
rect 330 219 332 221
rect 336 219 338 221
rect 360 219 362 221
rect 366 219 368 221
rect 390 219 392 221
rect 396 219 398 221
rect 420 219 422 221
rect 426 219 428 221
rect 450 219 452 221
rect 456 219 458 221
rect 480 219 482 221
rect 486 219 488 221
rect 510 219 512 221
rect 516 219 518 221
rect 540 219 542 221
rect 546 219 548 221
rect 68 217 70 219
rect 98 217 100 219
rect 128 217 130 219
rect 158 217 160 219
rect 188 217 190 219
rect 218 217 220 219
rect 248 217 250 219
rect 278 217 280 219
rect 308 217 310 219
rect 338 217 340 219
rect 368 217 370 219
rect 398 217 400 219
rect 428 217 430 219
rect 458 217 460 219
rect 488 217 490 219
rect 518 217 520 219
rect 548 217 550 219
rect 68 211 70 213
rect 98 211 100 213
rect 128 211 130 213
rect 158 211 160 213
rect 188 211 190 213
rect 218 211 220 213
rect 248 211 250 213
rect 278 211 280 213
rect 308 211 310 213
rect 338 211 340 213
rect 368 211 370 213
rect 398 211 400 213
rect 428 211 430 213
rect 458 211 460 213
rect 488 211 490 213
rect 518 211 520 213
rect 548 211 550 213
rect 60 209 62 211
rect 66 209 68 211
rect 90 209 92 211
rect 96 209 98 211
rect 120 209 122 211
rect 126 209 128 211
rect 150 209 152 211
rect 156 209 158 211
rect 180 209 182 211
rect 186 209 188 211
rect 210 209 212 211
rect 216 209 218 211
rect 240 209 242 211
rect 246 209 248 211
rect 270 209 272 211
rect 276 209 278 211
rect 300 209 302 211
rect 306 209 308 211
rect 330 209 332 211
rect 336 209 338 211
rect 360 209 362 211
rect 366 209 368 211
rect 390 209 392 211
rect 396 209 398 211
rect 420 209 422 211
rect 426 209 428 211
rect 450 209 452 211
rect 456 209 458 211
rect 480 209 482 211
rect 486 209 488 211
rect 510 209 512 211
rect 516 209 518 211
rect 540 209 542 211
rect 546 209 548 211
rect 58 207 60 209
rect 88 207 90 209
rect 118 207 120 209
rect 148 207 150 209
rect 178 207 180 209
rect 208 207 210 209
rect 238 207 240 209
rect 268 207 270 209
rect 298 207 300 209
rect 328 207 330 209
rect 358 207 360 209
rect 388 207 390 209
rect 418 207 420 209
rect 448 207 450 209
rect 478 207 480 209
rect 508 207 510 209
rect 538 207 540 209
rect 58 201 60 203
rect 88 201 90 203
rect 118 201 120 203
rect 148 201 150 203
rect 178 201 180 203
rect 208 201 210 203
rect 238 201 240 203
rect 268 201 270 203
rect 298 201 300 203
rect 328 201 330 203
rect 358 201 360 203
rect 388 201 390 203
rect 418 201 420 203
rect 448 201 450 203
rect 478 201 480 203
rect 508 201 510 203
rect 538 201 540 203
rect 60 199 62 201
rect 66 199 68 201
rect 90 199 92 201
rect 96 199 98 201
rect 120 199 122 201
rect 126 199 128 201
rect 150 199 152 201
rect 156 199 158 201
rect 180 199 182 201
rect 186 199 188 201
rect 210 199 212 201
rect 216 199 218 201
rect 240 199 242 201
rect 246 199 248 201
rect 270 199 272 201
rect 276 199 278 201
rect 300 199 302 201
rect 306 199 308 201
rect 330 199 332 201
rect 336 199 338 201
rect 360 199 362 201
rect 366 199 368 201
rect 390 199 392 201
rect 396 199 398 201
rect 420 199 422 201
rect 426 199 428 201
rect 450 199 452 201
rect 456 199 458 201
rect 480 199 482 201
rect 486 199 488 201
rect 510 199 512 201
rect 516 199 518 201
rect 540 199 542 201
rect 546 199 548 201
rect 68 197 70 199
rect 98 197 100 199
rect 128 197 130 199
rect 158 197 160 199
rect 188 197 190 199
rect 218 197 220 199
rect 248 197 250 199
rect 278 197 280 199
rect 308 197 310 199
rect 338 197 340 199
rect 368 197 370 199
rect 398 197 400 199
rect 428 197 430 199
rect 458 197 460 199
rect 488 197 490 199
rect 518 197 520 199
rect 548 197 550 199
rect 68 191 70 193
rect 98 191 100 193
rect 128 191 130 193
rect 158 191 160 193
rect 188 191 190 193
rect 218 191 220 193
rect 248 191 250 193
rect 278 191 280 193
rect 308 191 310 193
rect 338 191 340 193
rect 368 191 370 193
rect 398 191 400 193
rect 428 191 430 193
rect 458 191 460 193
rect 488 191 490 193
rect 518 191 520 193
rect 548 191 550 193
rect 60 189 62 191
rect 66 189 68 191
rect 90 189 92 191
rect 96 189 98 191
rect 120 189 122 191
rect 126 189 128 191
rect 150 189 152 191
rect 156 189 158 191
rect 180 189 182 191
rect 186 189 188 191
rect 210 189 212 191
rect 216 189 218 191
rect 240 189 242 191
rect 246 189 248 191
rect 270 189 272 191
rect 276 189 278 191
rect 300 189 302 191
rect 306 189 308 191
rect 330 189 332 191
rect 336 189 338 191
rect 360 189 362 191
rect 366 189 368 191
rect 390 189 392 191
rect 396 189 398 191
rect 420 189 422 191
rect 426 189 428 191
rect 450 189 452 191
rect 456 189 458 191
rect 480 189 482 191
rect 486 189 488 191
rect 510 189 512 191
rect 516 189 518 191
rect 540 189 542 191
rect 546 189 548 191
rect 58 187 60 189
rect 88 187 90 189
rect 118 187 120 189
rect 148 187 150 189
rect 178 187 180 189
rect 208 187 210 189
rect 238 187 240 189
rect 268 187 270 189
rect 298 187 300 189
rect 328 187 330 189
rect 358 187 360 189
rect 388 187 390 189
rect 418 187 420 189
rect 448 187 450 189
rect 478 187 480 189
rect 508 187 510 189
rect 538 187 540 189
rect 58 181 60 183
rect 88 181 90 183
rect 118 181 120 183
rect 148 181 150 183
rect 178 181 180 183
rect 208 181 210 183
rect 238 181 240 183
rect 268 181 270 183
rect 298 181 300 183
rect 328 181 330 183
rect 358 181 360 183
rect 388 181 390 183
rect 418 181 420 183
rect 448 181 450 183
rect 478 181 480 183
rect 508 181 510 183
rect 538 181 540 183
rect 60 179 62 181
rect 66 179 68 181
rect 90 179 92 181
rect 96 179 98 181
rect 120 179 122 181
rect 126 179 128 181
rect 150 179 152 181
rect 156 179 158 181
rect 180 179 182 181
rect 186 179 188 181
rect 210 179 212 181
rect 216 179 218 181
rect 240 179 242 181
rect 246 179 248 181
rect 270 179 272 181
rect 276 179 278 181
rect 300 179 302 181
rect 306 179 308 181
rect 330 179 332 181
rect 336 179 338 181
rect 360 179 362 181
rect 366 179 368 181
rect 390 179 392 181
rect 396 179 398 181
rect 420 179 422 181
rect 426 179 428 181
rect 450 179 452 181
rect 456 179 458 181
rect 480 179 482 181
rect 486 179 488 181
rect 510 179 512 181
rect 516 179 518 181
rect 540 179 542 181
rect 546 179 548 181
rect 68 177 70 179
rect 98 177 100 179
rect 128 177 130 179
rect 158 177 160 179
rect 188 177 190 179
rect 218 177 220 179
rect 248 177 250 179
rect 278 177 280 179
rect 308 177 310 179
rect 338 177 340 179
rect 368 177 370 179
rect 398 177 400 179
rect 428 177 430 179
rect 458 177 460 179
rect 488 177 490 179
rect 518 177 520 179
rect 548 177 550 179
rect 68 171 70 173
rect 98 171 100 173
rect 128 171 130 173
rect 158 171 160 173
rect 188 171 190 173
rect 218 171 220 173
rect 248 171 250 173
rect 278 171 280 173
rect 308 171 310 173
rect 338 171 340 173
rect 368 171 370 173
rect 398 171 400 173
rect 428 171 430 173
rect 458 171 460 173
rect 488 171 490 173
rect 518 171 520 173
rect 548 171 550 173
rect 60 169 62 171
rect 66 169 68 171
rect 90 169 92 171
rect 96 169 98 171
rect 120 169 122 171
rect 126 169 128 171
rect 150 169 152 171
rect 156 169 158 171
rect 180 169 182 171
rect 186 169 188 171
rect 210 169 212 171
rect 216 169 218 171
rect 240 169 242 171
rect 246 169 248 171
rect 270 169 272 171
rect 276 169 278 171
rect 300 169 302 171
rect 306 169 308 171
rect 330 169 332 171
rect 336 169 338 171
rect 360 169 362 171
rect 366 169 368 171
rect 390 169 392 171
rect 396 169 398 171
rect 420 169 422 171
rect 426 169 428 171
rect 450 169 452 171
rect 456 169 458 171
rect 480 169 482 171
rect 486 169 488 171
rect 510 169 512 171
rect 516 169 518 171
rect 540 169 542 171
rect 546 169 548 171
rect 58 167 60 169
rect 88 167 90 169
rect 118 167 120 169
rect 148 167 150 169
rect 178 167 180 169
rect 208 167 210 169
rect 238 167 240 169
rect 268 167 270 169
rect 298 167 300 169
rect 328 167 330 169
rect 358 167 360 169
rect 388 167 390 169
rect 418 167 420 169
rect 448 167 450 169
rect 478 167 480 169
rect 508 167 510 169
rect 538 167 540 169
rect 58 161 60 163
rect 88 161 90 163
rect 508 161 510 163
rect 538 161 540 163
rect 60 159 62 161
rect 66 159 68 161
rect 90 159 92 161
rect 506 159 508 161
rect 540 159 542 161
rect 546 159 548 161
rect 68 157 70 159
rect 548 157 550 159
rect 68 151 70 153
rect 548 151 550 153
rect 60 149 62 151
rect 66 149 68 151
rect 90 149 92 151
rect 506 149 508 151
rect 540 149 542 151
rect 546 149 548 151
rect 58 147 60 149
rect 88 147 90 149
rect 508 147 510 149
rect 538 147 540 149
rect 58 141 60 143
rect 88 141 90 143
rect 118 141 120 143
rect 148 141 150 143
rect 178 141 180 143
rect 208 141 210 143
rect 238 141 240 143
rect 268 141 270 143
rect 298 141 300 143
rect 328 141 330 143
rect 358 141 360 143
rect 388 141 390 143
rect 418 141 420 143
rect 448 141 450 143
rect 478 141 480 143
rect 508 141 510 143
rect 538 141 540 143
rect 60 139 62 141
rect 66 139 68 141
rect 90 139 92 141
rect 96 139 98 141
rect 120 139 122 141
rect 126 139 128 141
rect 150 139 152 141
rect 156 139 158 141
rect 180 139 182 141
rect 186 139 188 141
rect 210 139 212 141
rect 216 139 218 141
rect 240 139 242 141
rect 246 139 248 141
rect 270 139 272 141
rect 276 139 278 141
rect 300 139 302 141
rect 306 139 308 141
rect 330 139 332 141
rect 336 139 338 141
rect 360 139 362 141
rect 366 139 368 141
rect 390 139 392 141
rect 396 139 398 141
rect 420 139 422 141
rect 426 139 428 141
rect 450 139 452 141
rect 456 139 458 141
rect 480 139 482 141
rect 486 139 488 141
rect 510 139 512 141
rect 516 139 518 141
rect 540 139 542 141
rect 546 139 548 141
rect 68 137 70 139
rect 98 137 100 139
rect 128 137 130 139
rect 158 137 160 139
rect 188 137 190 139
rect 218 137 220 139
rect 248 137 250 139
rect 278 137 280 139
rect 308 137 310 139
rect 338 137 340 139
rect 368 137 370 139
rect 398 137 400 139
rect 428 137 430 139
rect 458 137 460 139
rect 488 137 490 139
rect 518 137 520 139
rect 548 137 550 139
rect 68 131 70 133
rect 98 131 100 133
rect 128 131 130 133
rect 158 131 160 133
rect 188 131 190 133
rect 218 131 220 133
rect 248 131 250 133
rect 278 131 280 133
rect 308 131 310 133
rect 338 131 340 133
rect 368 131 370 133
rect 398 131 400 133
rect 428 131 430 133
rect 458 131 460 133
rect 488 131 490 133
rect 518 131 520 133
rect 548 131 550 133
rect 60 129 62 131
rect 66 129 68 131
rect 90 129 92 131
rect 96 129 98 131
rect 120 129 122 131
rect 126 129 128 131
rect 150 129 152 131
rect 156 129 158 131
rect 180 129 182 131
rect 186 129 188 131
rect 210 129 212 131
rect 216 129 218 131
rect 240 129 242 131
rect 246 129 248 131
rect 270 129 272 131
rect 276 129 278 131
rect 300 129 302 131
rect 306 129 308 131
rect 330 129 332 131
rect 336 129 338 131
rect 360 129 362 131
rect 366 129 368 131
rect 390 129 392 131
rect 396 129 398 131
rect 420 129 422 131
rect 426 129 428 131
rect 450 129 452 131
rect 456 129 458 131
rect 480 129 482 131
rect 486 129 488 131
rect 510 129 512 131
rect 516 129 518 131
rect 540 129 542 131
rect 546 129 548 131
rect 58 127 60 129
rect 88 127 90 129
rect 118 127 120 129
rect 148 127 150 129
rect 178 127 180 129
rect 208 127 210 129
rect 238 127 240 129
rect 268 127 270 129
rect 298 127 300 129
rect 328 127 330 129
rect 358 127 360 129
rect 388 127 390 129
rect 418 127 420 129
rect 448 127 450 129
rect 478 127 480 129
rect 508 127 510 129
rect 538 127 540 129
rect 58 121 60 123
rect 88 121 90 123
rect 118 121 120 123
rect 148 121 150 123
rect 178 121 180 123
rect 208 121 210 123
rect 238 121 240 123
rect 268 121 270 123
rect 298 121 300 123
rect 328 121 330 123
rect 358 121 360 123
rect 388 121 390 123
rect 418 121 420 123
rect 448 121 450 123
rect 478 121 480 123
rect 508 121 510 123
rect 538 121 540 123
rect 60 119 62 121
rect 66 119 68 121
rect 90 119 92 121
rect 96 119 98 121
rect 120 119 122 121
rect 126 119 128 121
rect 150 119 152 121
rect 156 119 158 121
rect 180 119 182 121
rect 186 119 188 121
rect 210 119 212 121
rect 216 119 218 121
rect 240 119 242 121
rect 246 119 248 121
rect 270 119 272 121
rect 276 119 278 121
rect 300 119 302 121
rect 306 119 308 121
rect 330 119 332 121
rect 336 119 338 121
rect 360 119 362 121
rect 366 119 368 121
rect 390 119 392 121
rect 396 119 398 121
rect 420 119 422 121
rect 426 119 428 121
rect 450 119 452 121
rect 456 119 458 121
rect 480 119 482 121
rect 486 119 488 121
rect 510 119 512 121
rect 516 119 518 121
rect 540 119 542 121
rect 546 119 548 121
rect 68 117 70 119
rect 98 117 100 119
rect 128 117 130 119
rect 158 117 160 119
rect 188 117 190 119
rect 218 117 220 119
rect 248 117 250 119
rect 278 117 280 119
rect 308 117 310 119
rect 338 117 340 119
rect 368 117 370 119
rect 398 117 400 119
rect 428 117 430 119
rect 458 117 460 119
rect 488 117 490 119
rect 518 117 520 119
rect 548 117 550 119
rect 68 111 70 113
rect 98 111 100 113
rect 128 111 130 113
rect 158 111 160 113
rect 188 111 190 113
rect 218 111 220 113
rect 248 111 250 113
rect 278 111 280 113
rect 308 111 310 113
rect 338 111 340 113
rect 368 111 370 113
rect 398 111 400 113
rect 428 111 430 113
rect 458 111 460 113
rect 488 111 490 113
rect 518 111 520 113
rect 548 111 550 113
rect 60 109 62 111
rect 66 109 68 111
rect 90 109 92 111
rect 96 109 98 111
rect 120 109 122 111
rect 126 109 128 111
rect 150 109 152 111
rect 156 109 158 111
rect 180 109 182 111
rect 186 109 188 111
rect 210 109 212 111
rect 216 109 218 111
rect 240 109 242 111
rect 246 109 248 111
rect 270 109 272 111
rect 276 109 278 111
rect 300 109 302 111
rect 306 109 308 111
rect 330 109 332 111
rect 336 109 338 111
rect 360 109 362 111
rect 366 109 368 111
rect 390 109 392 111
rect 396 109 398 111
rect 420 109 422 111
rect 426 109 428 111
rect 450 109 452 111
rect 456 109 458 111
rect 480 109 482 111
rect 486 109 488 111
rect 510 109 512 111
rect 516 109 518 111
rect 540 109 542 111
rect 546 109 548 111
rect 58 107 60 109
rect 88 107 90 109
rect 118 107 120 109
rect 148 107 150 109
rect 178 107 180 109
rect 208 107 210 109
rect 238 107 240 109
rect 268 107 270 109
rect 298 107 300 109
rect 328 107 330 109
rect 358 107 360 109
rect 388 107 390 109
rect 418 107 420 109
rect 448 107 450 109
rect 478 107 480 109
rect 508 107 510 109
rect 538 107 540 109
rect 58 101 60 103
rect 88 101 90 103
rect 118 101 120 103
rect 148 101 150 103
rect 178 101 180 103
rect 208 101 210 103
rect 238 101 240 103
rect 268 101 270 103
rect 298 101 300 103
rect 328 101 330 103
rect 358 101 360 103
rect 388 101 390 103
rect 418 101 420 103
rect 448 101 450 103
rect 478 101 480 103
rect 508 101 510 103
rect 538 101 540 103
rect 60 99 62 101
rect 66 99 68 101
rect 90 99 92 101
rect 96 99 98 101
rect 120 99 122 101
rect 126 99 128 101
rect 150 99 152 101
rect 156 99 158 101
rect 180 99 182 101
rect 186 99 188 101
rect 210 99 212 101
rect 216 99 218 101
rect 240 99 242 101
rect 246 99 248 101
rect 270 99 272 101
rect 276 99 278 101
rect 300 99 302 101
rect 306 99 308 101
rect 330 99 332 101
rect 336 99 338 101
rect 360 99 362 101
rect 366 99 368 101
rect 390 99 392 101
rect 396 99 398 101
rect 420 99 422 101
rect 426 99 428 101
rect 450 99 452 101
rect 456 99 458 101
rect 480 99 482 101
rect 486 99 488 101
rect 510 99 512 101
rect 516 99 518 101
rect 540 99 542 101
rect 546 99 548 101
rect 68 97 70 99
rect 98 97 100 99
rect 128 97 130 99
rect 158 97 160 99
rect 188 97 190 99
rect 218 97 220 99
rect 248 97 250 99
rect 278 97 280 99
rect 308 97 310 99
rect 338 97 340 99
rect 368 97 370 99
rect 398 97 400 99
rect 428 97 430 99
rect 458 97 460 99
rect 488 97 490 99
rect 518 97 520 99
rect 548 97 550 99
rect 68 91 70 93
rect 98 91 100 93
rect 128 91 130 93
rect 158 91 160 93
rect 188 91 190 93
rect 218 91 220 93
rect 248 91 250 93
rect 278 91 280 93
rect 308 91 310 93
rect 338 91 340 93
rect 368 91 370 93
rect 398 91 400 93
rect 428 91 430 93
rect 458 91 460 93
rect 488 91 490 93
rect 518 91 520 93
rect 548 91 550 93
rect 60 89 62 91
rect 66 89 68 91
rect 90 89 92 91
rect 96 89 98 91
rect 120 89 122 91
rect 126 89 128 91
rect 150 89 152 91
rect 156 89 158 91
rect 180 89 182 91
rect 186 89 188 91
rect 210 89 212 91
rect 216 89 218 91
rect 240 89 242 91
rect 246 89 248 91
rect 270 89 272 91
rect 276 89 278 91
rect 300 89 302 91
rect 306 89 308 91
rect 330 89 332 91
rect 336 89 338 91
rect 360 89 362 91
rect 366 89 368 91
rect 390 89 392 91
rect 396 89 398 91
rect 420 89 422 91
rect 426 89 428 91
rect 450 89 452 91
rect 456 89 458 91
rect 480 89 482 91
rect 486 89 488 91
rect 510 89 512 91
rect 516 89 518 91
rect 540 89 542 91
rect 546 89 548 91
rect 58 87 60 89
rect 88 87 90 89
rect 118 87 120 89
rect 148 87 150 89
rect 178 87 180 89
rect 208 87 210 89
rect 238 87 240 89
rect 268 87 270 89
rect 298 87 300 89
rect 328 87 330 89
rect 358 87 360 89
rect 388 87 390 89
rect 418 87 420 89
rect 448 87 450 89
rect 478 87 480 89
rect 508 87 510 89
rect 538 87 540 89
rect 58 81 60 83
rect 88 81 90 83
rect 118 81 120 83
rect 148 81 150 83
rect 178 81 180 83
rect 208 81 210 83
rect 238 81 240 83
rect 268 81 270 83
rect 298 81 300 83
rect 328 81 330 83
rect 358 81 360 83
rect 388 81 390 83
rect 418 81 420 83
rect 448 81 450 83
rect 478 81 480 83
rect 508 81 510 83
rect 538 81 540 83
rect 60 79 62 81
rect 66 79 68 81
rect 90 79 92 81
rect 96 79 98 81
rect 120 79 122 81
rect 126 79 128 81
rect 150 79 152 81
rect 156 79 158 81
rect 180 79 182 81
rect 186 79 188 81
rect 210 79 212 81
rect 216 79 218 81
rect 240 79 242 81
rect 246 79 248 81
rect 270 79 272 81
rect 276 79 278 81
rect 300 79 302 81
rect 306 79 308 81
rect 330 79 332 81
rect 336 79 338 81
rect 360 79 362 81
rect 366 79 368 81
rect 390 79 392 81
rect 396 79 398 81
rect 420 79 422 81
rect 426 79 428 81
rect 450 79 452 81
rect 456 79 458 81
rect 480 79 482 81
rect 486 79 488 81
rect 510 79 512 81
rect 516 79 518 81
rect 540 79 542 81
rect 546 79 548 81
rect 68 77 70 79
rect 98 77 100 79
rect 128 77 130 79
rect 158 77 160 79
rect 188 77 190 79
rect 218 77 220 79
rect 248 77 250 79
rect 278 77 280 79
rect 308 77 310 79
rect 338 77 340 79
rect 368 77 370 79
rect 398 77 400 79
rect 428 77 430 79
rect 458 77 460 79
rect 488 77 490 79
rect 518 77 520 79
rect 548 77 550 79
rect 68 71 70 73
rect 98 71 100 73
rect 128 71 130 73
rect 158 71 160 73
rect 188 71 190 73
rect 218 71 220 73
rect 248 71 250 73
rect 278 71 280 73
rect 308 71 310 73
rect 338 71 340 73
rect 368 71 370 73
rect 398 71 400 73
rect 428 71 430 73
rect 458 71 460 73
rect 488 71 490 73
rect 518 71 520 73
rect 548 71 550 73
rect 60 69 62 71
rect 66 69 68 71
rect 90 69 92 71
rect 96 69 98 71
rect 120 69 122 71
rect 126 69 128 71
rect 150 69 152 71
rect 156 69 158 71
rect 180 69 182 71
rect 186 69 188 71
rect 210 69 212 71
rect 216 69 218 71
rect 240 69 242 71
rect 246 69 248 71
rect 270 69 272 71
rect 276 69 278 71
rect 300 69 302 71
rect 306 69 308 71
rect 330 69 332 71
rect 336 69 338 71
rect 360 69 362 71
rect 366 69 368 71
rect 390 69 392 71
rect 396 69 398 71
rect 420 69 422 71
rect 426 69 428 71
rect 450 69 452 71
rect 456 69 458 71
rect 480 69 482 71
rect 486 69 488 71
rect 510 69 512 71
rect 516 69 518 71
rect 540 69 542 71
rect 546 69 548 71
rect 58 67 60 69
rect 88 67 90 69
rect 118 67 120 69
rect 148 67 150 69
rect 178 67 180 69
rect 208 67 210 69
rect 238 67 240 69
rect 268 67 270 69
rect 298 67 300 69
rect 328 67 330 69
rect 358 67 360 69
rect 388 67 390 69
rect 418 67 420 69
rect 448 67 450 69
rect 478 67 480 69
rect 508 67 510 69
rect 538 67 540 69
rect 58 61 60 63
rect 88 61 90 63
rect 118 61 120 63
rect 148 61 150 63
rect 178 61 180 63
rect 208 61 210 63
rect 238 61 240 63
rect 268 61 270 63
rect 298 61 300 63
rect 328 61 330 63
rect 358 61 360 63
rect 388 61 390 63
rect 418 61 420 63
rect 448 61 450 63
rect 478 61 480 63
rect 508 61 510 63
rect 538 61 540 63
rect 60 59 62 61
rect 66 59 68 61
rect 90 59 92 61
rect 96 59 98 61
rect 120 59 122 61
rect 126 59 128 61
rect 150 59 152 61
rect 156 59 158 61
rect 180 59 182 61
rect 186 59 188 61
rect 210 59 212 61
rect 216 59 218 61
rect 240 59 242 61
rect 246 59 248 61
rect 270 59 272 61
rect 276 59 278 61
rect 300 59 302 61
rect 306 59 308 61
rect 330 59 332 61
rect 336 59 338 61
rect 360 59 362 61
rect 366 59 368 61
rect 390 59 392 61
rect 396 59 398 61
rect 420 59 422 61
rect 426 59 428 61
rect 450 59 452 61
rect 456 59 458 61
rect 480 59 482 61
rect 486 59 488 61
rect 510 59 512 61
rect 516 59 518 61
rect 540 59 542 61
rect 546 59 548 61
rect 68 57 70 59
rect 98 57 100 59
rect 128 57 130 59
rect 158 57 160 59
rect 188 57 190 59
rect 218 57 220 59
rect 248 57 250 59
rect 278 57 280 59
rect 308 57 310 59
rect 338 57 340 59
rect 368 57 370 59
rect 398 57 400 59
rect 428 57 430 59
rect 458 57 460 59
rect 488 57 490 59
rect 518 57 520 59
rect 548 57 550 59
rect 68 51 70 53
rect 98 51 100 53
rect 128 51 130 53
rect 158 51 160 53
rect 188 51 190 53
rect 218 51 220 53
rect 248 51 250 53
rect 278 51 280 53
rect 308 51 310 53
rect 338 51 340 53
rect 368 51 370 53
rect 398 51 400 53
rect 428 51 430 53
rect 458 51 460 53
rect 488 51 490 53
rect 518 51 520 53
rect 548 51 550 53
rect 60 49 62 51
rect 66 49 68 51
rect 90 49 92 51
rect 96 49 98 51
rect 120 49 122 51
rect 126 49 128 51
rect 150 49 152 51
rect 156 49 158 51
rect 180 49 182 51
rect 186 49 188 51
rect 210 49 212 51
rect 216 49 218 51
rect 240 49 242 51
rect 246 49 248 51
rect 270 49 272 51
rect 276 49 278 51
rect 300 49 302 51
rect 306 49 308 51
rect 330 49 332 51
rect 336 49 338 51
rect 360 49 362 51
rect 366 49 368 51
rect 390 49 392 51
rect 396 49 398 51
rect 420 49 422 51
rect 426 49 428 51
rect 450 49 452 51
rect 456 49 458 51
rect 480 49 482 51
rect 486 49 488 51
rect 510 49 512 51
rect 516 49 518 51
rect 540 49 542 51
rect 546 49 548 51
rect 58 47 60 49
rect 88 47 90 49
rect 118 47 120 49
rect 148 47 150 49
rect 178 47 180 49
rect 208 47 210 49
rect 238 47 240 49
rect 268 47 270 49
rect 298 47 300 49
rect 328 47 330 49
rect 358 47 360 49
rect 388 47 390 49
rect 418 47 420 49
rect 448 47 450 49
rect 478 47 480 49
rect 508 47 510 49
rect 538 47 540 49
rect 58 41 60 43
rect 88 41 90 43
rect 118 41 120 43
rect 148 41 150 43
rect 178 41 180 43
rect 208 41 210 43
rect 238 41 240 43
rect 268 41 270 43
rect 298 41 300 43
rect 328 41 330 43
rect 358 41 360 43
rect 388 41 390 43
rect 418 41 420 43
rect 448 41 450 43
rect 478 41 480 43
rect 508 41 510 43
rect 538 41 540 43
rect 60 39 62 41
rect 66 39 68 41
rect 90 39 92 41
rect 96 39 98 41
rect 120 39 122 41
rect 126 39 128 41
rect 150 39 152 41
rect 156 39 158 41
rect 180 39 182 41
rect 186 39 188 41
rect 210 39 212 41
rect 216 39 218 41
rect 240 39 242 41
rect 246 39 248 41
rect 270 39 272 41
rect 276 39 278 41
rect 300 39 302 41
rect 306 39 308 41
rect 330 39 332 41
rect 336 39 338 41
rect 360 39 362 41
rect 366 39 368 41
rect 390 39 392 41
rect 396 39 398 41
rect 420 39 422 41
rect 426 39 428 41
rect 450 39 452 41
rect 456 39 458 41
rect 480 39 482 41
rect 486 39 488 41
rect 510 39 512 41
rect 516 39 518 41
rect 540 39 542 41
rect 546 39 548 41
rect 68 37 70 39
rect 98 37 100 39
rect 128 37 130 39
rect 158 37 160 39
rect 188 37 190 39
rect 218 37 220 39
rect 248 37 250 39
rect 278 37 280 39
rect 308 37 310 39
rect 338 37 340 39
rect 368 37 370 39
rect 398 37 400 39
rect 428 37 430 39
rect 458 37 460 39
rect 488 37 490 39
rect 518 37 520 39
rect 548 37 550 39
rect 10 12 12 14
rect 588 12 590 14
rect 12 10 14 12
rect 586 10 588 12
<< error_s >>
rect 110 1598 118 1600
rect 134 1598 142 1600
rect 158 1598 166 1600
rect 182 1598 190 1600
rect 206 1598 214 1600
rect 230 1598 238 1600
rect 254 1598 262 1600
rect 278 1598 286 1600
rect 302 1598 310 1600
rect 326 1598 334 1600
rect 350 1598 358 1600
rect 374 1598 382 1600
rect 398 1598 406 1600
rect 422 1598 430 1600
rect 446 1598 454 1600
rect 470 1598 478 1600
rect 494 1598 502 1600
rect 98 1592 106 1594
rect 98 1588 100 1592
rect 104 1588 106 1592
rect 98 1586 106 1588
rect 122 1592 130 1594
rect 122 1588 124 1592
rect 128 1588 130 1592
rect 122 1586 130 1588
rect 146 1592 154 1594
rect 146 1588 148 1592
rect 152 1588 154 1592
rect 146 1586 154 1588
rect 170 1592 178 1594
rect 170 1588 172 1592
rect 176 1588 178 1592
rect 170 1586 178 1588
rect 194 1592 202 1594
rect 194 1588 196 1592
rect 200 1588 202 1592
rect 194 1586 202 1588
rect 218 1592 226 1594
rect 218 1588 220 1592
rect 224 1588 226 1592
rect 218 1586 226 1588
rect 242 1592 250 1594
rect 242 1588 244 1592
rect 248 1588 250 1592
rect 242 1586 250 1588
rect 266 1592 274 1594
rect 266 1588 268 1592
rect 272 1588 274 1592
rect 266 1586 274 1588
rect 290 1592 298 1594
rect 290 1588 292 1592
rect 296 1588 298 1592
rect 290 1586 298 1588
rect 314 1592 322 1594
rect 314 1588 316 1592
rect 320 1588 322 1592
rect 314 1586 322 1588
rect 338 1592 346 1594
rect 338 1588 340 1592
rect 344 1588 346 1592
rect 338 1586 346 1588
rect 362 1592 370 1594
rect 362 1588 364 1592
rect 368 1588 370 1592
rect 362 1586 370 1588
rect 386 1592 394 1594
rect 386 1588 388 1592
rect 392 1588 394 1592
rect 386 1586 394 1588
rect 410 1592 418 1594
rect 410 1588 412 1592
rect 416 1588 418 1592
rect 410 1586 418 1588
rect 434 1592 442 1594
rect 434 1588 436 1592
rect 440 1588 442 1592
rect 434 1586 442 1588
rect 458 1592 466 1594
rect 458 1588 460 1592
rect 464 1588 466 1592
rect 458 1586 466 1588
rect 482 1592 490 1594
rect 482 1588 484 1592
rect 488 1588 490 1592
rect 482 1586 490 1588
rect 110 1580 118 1582
rect 110 1576 112 1580
rect 116 1576 118 1580
rect 110 1574 118 1576
rect 134 1580 142 1582
rect 134 1576 136 1580
rect 140 1576 142 1580
rect 134 1574 142 1576
rect 158 1580 166 1582
rect 158 1576 160 1580
rect 164 1576 166 1580
rect 158 1574 166 1576
rect 182 1580 190 1582
rect 182 1576 184 1580
rect 188 1576 190 1580
rect 182 1574 190 1576
rect 206 1580 214 1582
rect 206 1576 208 1580
rect 212 1576 214 1580
rect 206 1574 214 1576
rect 230 1580 238 1582
rect 230 1576 232 1580
rect 236 1576 238 1580
rect 230 1574 238 1576
rect 254 1580 262 1582
rect 254 1576 256 1580
rect 260 1576 262 1580
rect 254 1574 262 1576
rect 278 1580 286 1582
rect 278 1576 280 1580
rect 284 1576 286 1580
rect 278 1574 286 1576
rect 302 1580 310 1582
rect 302 1576 304 1580
rect 308 1576 310 1580
rect 302 1574 310 1576
rect 326 1580 334 1582
rect 326 1576 328 1580
rect 332 1576 334 1580
rect 326 1574 334 1576
rect 350 1580 358 1582
rect 350 1576 352 1580
rect 356 1576 358 1580
rect 350 1574 358 1576
rect 374 1580 382 1582
rect 374 1576 376 1580
rect 380 1576 382 1580
rect 374 1574 382 1576
rect 398 1580 406 1582
rect 398 1576 400 1580
rect 404 1576 406 1580
rect 398 1574 406 1576
rect 422 1580 430 1582
rect 422 1576 424 1580
rect 428 1576 430 1580
rect 422 1574 430 1576
rect 446 1580 454 1582
rect 446 1576 448 1580
rect 452 1576 454 1580
rect 446 1574 454 1576
rect 470 1580 478 1582
rect 470 1576 472 1580
rect 476 1576 478 1580
rect 470 1574 478 1576
rect 494 1580 502 1582
rect 494 1576 496 1580
rect 500 1576 502 1580
rect 494 1574 502 1576
rect 98 1568 106 1570
rect 98 1564 100 1568
rect 104 1564 106 1568
rect 98 1562 106 1564
rect 122 1568 130 1570
rect 122 1564 124 1568
rect 128 1564 130 1568
rect 122 1562 130 1564
rect 146 1568 154 1570
rect 146 1564 148 1568
rect 152 1564 154 1568
rect 146 1562 154 1564
rect 170 1568 178 1570
rect 170 1564 172 1568
rect 176 1564 178 1568
rect 170 1562 178 1564
rect 194 1568 202 1570
rect 194 1564 196 1568
rect 200 1564 202 1568
rect 194 1562 202 1564
rect 218 1568 226 1570
rect 218 1564 220 1568
rect 224 1564 226 1568
rect 218 1562 226 1564
rect 242 1568 250 1570
rect 242 1564 244 1568
rect 248 1564 250 1568
rect 242 1562 250 1564
rect 266 1568 274 1570
rect 266 1564 268 1568
rect 272 1564 274 1568
rect 266 1562 274 1564
rect 290 1568 298 1570
rect 290 1564 292 1568
rect 296 1564 298 1568
rect 290 1562 298 1564
rect 314 1568 322 1570
rect 314 1564 316 1568
rect 320 1564 322 1568
rect 314 1562 322 1564
rect 338 1568 346 1570
rect 338 1564 340 1568
rect 344 1564 346 1568
rect 338 1562 346 1564
rect 362 1568 370 1570
rect 362 1564 364 1568
rect 368 1564 370 1568
rect 362 1562 370 1564
rect 386 1568 394 1570
rect 386 1564 388 1568
rect 392 1564 394 1568
rect 386 1562 394 1564
rect 410 1568 418 1570
rect 410 1564 412 1568
rect 416 1564 418 1568
rect 410 1562 418 1564
rect 434 1568 442 1570
rect 434 1564 436 1568
rect 440 1564 442 1568
rect 434 1562 442 1564
rect 458 1568 466 1570
rect 458 1564 460 1568
rect 464 1564 466 1568
rect 458 1562 466 1564
rect 482 1568 490 1570
rect 482 1564 484 1568
rect 488 1564 490 1568
rect 482 1562 490 1564
rect 110 1556 118 1558
rect 110 1552 112 1556
rect 116 1552 118 1556
rect 110 1550 118 1552
rect 134 1556 142 1558
rect 134 1552 136 1556
rect 140 1552 142 1556
rect 134 1550 142 1552
rect 158 1556 166 1558
rect 158 1552 160 1556
rect 164 1552 166 1556
rect 158 1550 166 1552
rect 182 1556 190 1558
rect 182 1552 184 1556
rect 188 1552 190 1556
rect 182 1550 190 1552
rect 206 1556 214 1558
rect 206 1552 208 1556
rect 212 1552 214 1556
rect 206 1550 214 1552
rect 230 1556 238 1558
rect 230 1552 232 1556
rect 236 1552 238 1556
rect 230 1550 238 1552
rect 254 1556 262 1558
rect 254 1552 256 1556
rect 260 1552 262 1556
rect 254 1550 262 1552
rect 278 1556 286 1558
rect 278 1552 280 1556
rect 284 1552 286 1556
rect 278 1550 286 1552
rect 302 1556 310 1558
rect 302 1552 304 1556
rect 308 1552 310 1556
rect 302 1550 310 1552
rect 326 1556 334 1558
rect 326 1552 328 1556
rect 332 1552 334 1556
rect 326 1550 334 1552
rect 350 1556 358 1558
rect 350 1552 352 1556
rect 356 1552 358 1556
rect 350 1550 358 1552
rect 374 1556 382 1558
rect 374 1552 376 1556
rect 380 1552 382 1556
rect 374 1550 382 1552
rect 398 1556 406 1558
rect 398 1552 400 1556
rect 404 1552 406 1556
rect 398 1550 406 1552
rect 422 1556 430 1558
rect 422 1552 424 1556
rect 428 1552 430 1556
rect 422 1550 430 1552
rect 446 1556 454 1558
rect 446 1552 448 1556
rect 452 1552 454 1556
rect 446 1550 454 1552
rect 470 1556 478 1558
rect 470 1552 472 1556
rect 476 1552 478 1556
rect 470 1550 478 1552
rect 494 1556 502 1558
rect 494 1552 496 1556
rect 500 1552 502 1556
rect 494 1550 502 1552
rect 98 1544 106 1546
rect 98 1540 100 1544
rect 104 1540 106 1544
rect 98 1538 106 1540
rect 122 1544 130 1546
rect 122 1540 124 1544
rect 128 1540 130 1544
rect 122 1538 130 1540
rect 146 1544 154 1546
rect 146 1540 148 1544
rect 152 1540 154 1544
rect 146 1538 154 1540
rect 170 1544 178 1546
rect 170 1540 172 1544
rect 176 1540 178 1544
rect 170 1538 178 1540
rect 194 1544 202 1546
rect 194 1540 196 1544
rect 200 1540 202 1544
rect 194 1538 202 1540
rect 218 1544 226 1546
rect 218 1540 220 1544
rect 224 1540 226 1544
rect 218 1538 226 1540
rect 242 1544 250 1546
rect 242 1540 244 1544
rect 248 1540 250 1544
rect 242 1538 250 1540
rect 266 1544 274 1546
rect 266 1540 268 1544
rect 272 1540 274 1544
rect 266 1538 274 1540
rect 290 1544 298 1546
rect 290 1540 292 1544
rect 296 1540 298 1544
rect 290 1538 298 1540
rect 314 1544 322 1546
rect 314 1540 316 1544
rect 320 1540 322 1544
rect 314 1538 322 1540
rect 338 1544 346 1546
rect 338 1540 340 1544
rect 344 1540 346 1544
rect 338 1538 346 1540
rect 362 1544 370 1546
rect 362 1540 364 1544
rect 368 1540 370 1544
rect 362 1538 370 1540
rect 386 1544 394 1546
rect 386 1540 388 1544
rect 392 1540 394 1544
rect 386 1538 394 1540
rect 410 1544 418 1546
rect 410 1540 412 1544
rect 416 1540 418 1544
rect 410 1538 418 1540
rect 434 1544 442 1546
rect 434 1540 436 1544
rect 440 1540 442 1544
rect 434 1538 442 1540
rect 458 1544 466 1546
rect 458 1540 460 1544
rect 464 1540 466 1544
rect 458 1538 466 1540
rect 482 1544 490 1546
rect 482 1540 484 1544
rect 488 1540 490 1544
rect 482 1538 490 1540
<< nwell >>
rect 34 858 566 1306
rect -6 498 606 660
rect -6 22 22 498
rect 578 22 606 498
rect -6 -6 606 22
<< ptransistor >>
rect 76 1252 276 1258
rect 324 1252 524 1258
rect 76 1164 276 1170
rect 76 1124 276 1130
rect 324 1164 524 1170
rect 324 1124 524 1130
rect 76 1036 276 1042
rect 76 994 276 1000
rect 324 1036 524 1042
rect 324 994 524 1000
rect 76 906 276 912
rect 324 906 524 912
<< pdiffusion >>
rect 76 1274 276 1276
rect 76 1266 82 1274
rect 240 1266 276 1274
rect 76 1258 276 1266
rect 76 1220 276 1252
rect 76 1202 112 1220
rect 240 1202 276 1220
rect 76 1170 276 1202
rect 324 1274 524 1276
rect 324 1266 360 1274
rect 518 1266 524 1274
rect 324 1258 524 1266
rect 76 1156 276 1164
rect 76 1138 82 1156
rect 240 1138 276 1156
rect 76 1130 276 1138
rect 76 1092 276 1124
rect 76 1074 112 1092
rect 240 1074 276 1092
rect 76 1042 276 1074
rect 324 1220 524 1252
rect 324 1202 360 1220
rect 488 1202 524 1220
rect 324 1170 524 1202
rect 324 1156 524 1164
rect 324 1138 360 1156
rect 518 1138 524 1156
rect 324 1130 524 1138
rect 76 1028 276 1036
rect 76 1020 82 1028
rect 240 1020 276 1028
rect 76 1016 276 1020
rect 76 1008 82 1016
rect 240 1008 276 1016
rect 76 1000 276 1008
rect 76 962 276 994
rect 76 944 112 962
rect 240 944 276 962
rect 76 912 276 944
rect 324 1092 524 1124
rect 324 1074 360 1092
rect 488 1074 524 1092
rect 324 1042 524 1074
rect 324 1028 524 1036
rect 324 1020 360 1028
rect 518 1020 524 1028
rect 324 1016 524 1020
rect 324 1008 360 1016
rect 518 1008 524 1016
rect 324 1000 524 1008
rect 76 898 276 906
rect 76 890 82 898
rect 240 890 276 898
rect 76 888 276 890
rect 324 962 524 994
rect 324 944 360 962
rect 488 944 524 962
rect 324 912 524 944
rect 324 898 524 906
rect 324 890 360 898
rect 518 890 524 898
rect 324 888 524 890
<< pdcontact >>
rect 82 1266 240 1274
rect 112 1202 240 1220
rect 360 1266 518 1274
rect 82 1138 240 1156
rect 112 1074 240 1092
rect 360 1202 488 1220
rect 360 1138 518 1156
rect 82 1020 240 1028
rect 82 1008 240 1016
rect 112 944 240 962
rect 360 1074 488 1092
rect 360 1020 518 1028
rect 360 1008 518 1016
rect 82 890 240 898
rect 360 944 488 962
rect 360 890 518 898
<< psubstratepdiff >>
rect 0 1338 600 1340
rect 0 840 2 1338
rect 260 1320 340 1338
rect 20 1318 580 1320
rect 20 846 22 1318
rect 578 846 580 1318
rect 20 844 580 846
rect 20 840 44 844
rect 0 836 44 840
rect 52 836 74 844
rect 82 836 104 844
rect 112 836 134 844
rect 142 836 164 844
rect 172 836 194 844
rect 202 836 224 844
rect 232 836 244 844
rect 262 836 274 844
rect 282 836 296 844
rect 304 836 318 844
rect 326 836 338 844
rect 356 836 368 844
rect 376 836 398 844
rect 406 836 428 844
rect 436 836 458 844
rect 466 836 488 844
rect 496 836 518 844
rect 526 836 548 844
rect 556 840 580 844
rect 598 840 600 1338
rect 556 836 600 840
rect 0 828 4 836
rect 12 828 24 836
rect 42 828 54 836
rect 72 828 84 836
rect 102 828 114 836
rect 132 828 144 836
rect 162 828 174 836
rect 192 828 204 836
rect 222 828 234 836
rect 242 828 264 836
rect 272 828 286 836
rect 294 828 306 836
rect 314 828 328 836
rect 336 828 358 836
rect 366 828 378 836
rect 396 828 408 836
rect 426 828 438 836
rect 456 828 468 836
rect 486 828 498 836
rect 516 828 528 836
rect 546 828 558 836
rect 576 828 588 836
rect 596 828 600 836
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 184 828
rect 192 826 214 828
rect 222 826 378 828
rect 386 826 408 828
rect 416 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 0 818 14 826
rect 22 818 34 826
rect 52 818 64 826
rect 82 818 94 826
rect 112 818 124 826
rect 142 818 154 826
rect 172 818 184 826
rect 202 818 214 826
rect 232 818 244 826
rect 262 818 274 826
rect 282 818 296 826
rect 304 818 318 826
rect 326 818 338 826
rect 356 818 368 826
rect 386 818 398 826
rect 416 818 428 826
rect 446 818 458 826
rect 476 818 488 826
rect 506 818 518 826
rect 536 818 548 826
rect 566 818 578 826
rect 586 818 600 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 184 818
rect 192 816 214 818
rect 222 816 378 818
rect 386 816 408 818
rect 416 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 0 808 4 816
rect 12 808 24 816
rect 42 808 54 816
rect 72 808 84 816
rect 102 808 114 816
rect 132 808 144 816
rect 162 808 174 816
rect 192 808 204 816
rect 222 808 234 816
rect 242 808 264 816
rect 272 808 286 816
rect 294 808 306 816
rect 314 808 328 816
rect 336 808 358 816
rect 366 808 378 816
rect 396 808 408 816
rect 426 808 438 816
rect 456 808 468 816
rect 486 808 498 816
rect 516 808 528 816
rect 546 808 558 816
rect 576 808 588 816
rect 596 808 600 816
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 184 808
rect 192 806 214 808
rect 222 806 378 808
rect 386 806 408 808
rect 416 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 0 798 14 806
rect 22 798 34 806
rect 52 798 64 806
rect 82 798 94 806
rect 112 798 124 806
rect 142 798 154 806
rect 172 798 184 806
rect 202 798 214 806
rect 232 798 244 806
rect 262 798 274 806
rect 282 798 296 806
rect 304 798 318 806
rect 326 798 338 806
rect 356 798 368 806
rect 386 798 398 806
rect 416 798 428 806
rect 446 798 458 806
rect 476 798 488 806
rect 506 798 518 806
rect 536 798 548 806
rect 566 798 578 806
rect 586 798 600 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 184 798
rect 192 796 214 798
rect 222 796 378 798
rect 386 796 408 798
rect 416 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 0 788 4 796
rect 12 788 24 796
rect 42 788 54 796
rect 72 788 84 796
rect 102 788 114 796
rect 132 788 144 796
rect 162 788 174 796
rect 192 788 204 796
rect 222 788 234 796
rect 242 788 264 796
rect 272 788 286 796
rect 294 788 306 796
rect 314 788 328 796
rect 336 788 358 796
rect 366 788 378 796
rect 396 788 408 796
rect 426 788 438 796
rect 456 788 468 796
rect 486 788 498 796
rect 516 788 528 796
rect 546 788 558 796
rect 576 788 588 796
rect 596 788 600 796
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 184 788
rect 192 786 214 788
rect 222 786 378 788
rect 386 786 408 788
rect 416 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 0 778 14 786
rect 22 778 34 786
rect 52 778 64 786
rect 82 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 776 124 786
rect 142 776 154 786
rect 172 776 184 786
rect 202 776 214 786
rect 232 776 244 786
rect 262 776 274 786
rect 282 776 296 786
rect 0 768 4 776
rect 12 768 24 776
rect 42 768 54 776
rect 72 768 84 776
rect 292 768 296 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 14 766
rect 22 758 34 766
rect 52 758 64 766
rect 82 758 94 766
rect 112 758 124 768
rect 142 758 154 768
rect 172 758 184 768
rect 202 758 214 768
rect 232 758 244 768
rect 262 758 274 768
rect 282 758 296 768
rect 304 776 318 786
rect 326 776 338 786
rect 356 776 368 786
rect 386 776 398 786
rect 416 776 428 786
rect 446 776 458 786
rect 476 776 488 786
rect 506 778 518 786
rect 536 778 548 786
rect 566 778 578 786
rect 586 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 304 768 308 776
rect 516 768 528 776
rect 546 768 558 776
rect 576 768 588 776
rect 596 768 600 776
rect 304 758 318 768
rect 326 758 338 768
rect 356 758 368 768
rect 386 758 398 768
rect 416 758 428 768
rect 446 758 458 768
rect 476 758 488 768
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 518 766
rect 536 758 548 766
rect 566 758 578 766
rect 586 758 600 766
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 184 758
rect 192 756 214 758
rect 222 756 378 758
rect 386 756 408 758
rect 416 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 0 748 4 756
rect 12 748 24 756
rect 42 748 54 756
rect 72 748 84 756
rect 102 748 114 756
rect 132 748 144 756
rect 162 748 174 756
rect 192 748 204 756
rect 222 748 234 756
rect 242 748 264 756
rect 272 748 286 756
rect 294 748 306 756
rect 314 748 328 756
rect 336 748 358 756
rect 366 748 378 756
rect 396 748 408 756
rect 426 748 438 756
rect 456 748 468 756
rect 486 748 498 756
rect 516 748 528 756
rect 546 748 558 756
rect 576 748 588 756
rect 596 748 600 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 184 748
rect 192 746 214 748
rect 222 746 378 748
rect 386 746 408 748
rect 416 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 0 738 14 746
rect 22 738 34 746
rect 52 738 64 746
rect 82 738 94 746
rect 112 738 124 746
rect 142 738 154 746
rect 172 738 184 746
rect 202 738 214 746
rect 232 738 244 746
rect 262 738 274 746
rect 282 738 296 746
rect 304 738 318 746
rect 326 738 338 746
rect 356 738 368 746
rect 386 738 398 746
rect 416 738 428 746
rect 446 738 458 746
rect 476 738 488 746
rect 506 738 518 746
rect 536 738 548 746
rect 566 738 578 746
rect 586 738 600 746
rect 0 736 214 738
rect 0 728 4 736
rect 12 728 24 736
rect 32 728 214 736
rect 0 726 214 728
rect 222 736 378 738
rect 222 728 234 736
rect 242 728 286 736
rect 294 728 306 736
rect 314 728 358 736
rect 366 728 378 736
rect 222 726 378 728
rect 386 736 600 738
rect 386 728 568 736
rect 576 728 588 736
rect 596 728 600 736
rect 386 726 600 728
rect 0 718 14 726
rect 22 718 34 726
rect 52 718 64 726
rect 82 718 94 726
rect 112 718 124 726
rect 142 718 154 726
rect 172 718 184 726
rect 202 718 214 726
rect 232 718 244 726
rect 262 718 296 726
rect 304 718 338 726
rect 356 718 368 726
rect 386 718 398 726
rect 416 718 428 726
rect 446 718 458 726
rect 476 718 488 726
rect 506 718 518 726
rect 536 718 548 726
rect 566 718 578 726
rect 586 718 600 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 184 718
rect 192 716 214 718
rect 222 716 378 718
rect 386 716 408 718
rect 416 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 0 708 4 716
rect 12 708 24 716
rect 42 708 54 716
rect 72 708 84 716
rect 102 708 114 716
rect 132 708 144 716
rect 162 708 174 716
rect 192 708 204 716
rect 222 708 234 716
rect 242 708 264 716
rect 272 708 286 716
rect 294 708 306 716
rect 314 708 328 716
rect 336 708 358 716
rect 366 708 378 716
rect 396 708 408 716
rect 426 708 438 716
rect 456 708 468 716
rect 486 708 498 716
rect 516 708 528 716
rect 546 708 558 716
rect 576 708 588 716
rect 596 708 600 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 184 708
rect 192 706 214 708
rect 222 706 378 708
rect 386 706 408 708
rect 416 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 0 698 14 706
rect 22 698 34 706
rect 52 698 64 706
rect 82 698 94 706
rect 112 698 124 706
rect 142 698 154 706
rect 172 698 184 706
rect 202 698 214 706
rect 232 698 244 706
rect 262 698 274 706
rect 282 698 296 706
rect 304 698 318 706
rect 326 698 338 706
rect 356 698 368 706
rect 386 698 398 706
rect 416 698 428 706
rect 446 698 458 706
rect 476 698 488 706
rect 506 698 518 706
rect 536 698 548 706
rect 566 698 578 706
rect 586 698 600 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 184 698
rect 192 696 214 698
rect 222 697 378 698
rect 222 696 286 697
rect 0 688 4 696
rect 12 688 24 696
rect 42 688 54 696
rect 72 688 84 696
rect 102 688 114 696
rect 132 688 144 696
rect 162 688 174 696
rect 192 688 204 696
rect 222 688 234 696
rect 242 689 286 696
rect 294 689 306 697
rect 314 696 378 697
rect 386 696 408 698
rect 416 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 314 689 358 696
rect 242 688 358 689
rect 366 688 378 696
rect 396 688 408 696
rect 426 688 438 696
rect 456 688 468 696
rect 486 688 498 696
rect 516 688 528 696
rect 546 688 558 696
rect 576 688 588 696
rect 596 688 600 696
rect 0 686 600 688
rect 28 489 572 492
rect 28 461 30 489
rect 568 461 572 489
rect 28 451 40 461
rect 48 451 60 461
rect 78 451 90 461
rect 108 451 120 461
rect 138 451 150 461
rect 168 451 180 461
rect 198 451 210 461
rect 228 451 240 461
rect 258 451 270 461
rect 288 451 300 461
rect 318 451 330 461
rect 348 451 360 461
rect 378 451 390 461
rect 408 451 420 461
rect 438 451 450 461
rect 468 451 480 461
rect 498 451 510 461
rect 528 451 540 461
rect 558 451 572 461
rect 28 449 60 451
rect 68 449 90 451
rect 98 449 120 451
rect 128 449 150 451
rect 158 449 180 451
rect 188 449 210 451
rect 218 449 240 451
rect 248 449 270 451
rect 278 449 300 451
rect 308 449 330 451
rect 338 449 360 451
rect 368 449 390 451
rect 398 449 420 451
rect 428 449 450 451
rect 458 449 480 451
rect 488 449 510 451
rect 518 449 540 451
rect 548 449 572 451
rect 28 441 30 449
rect 38 441 50 449
rect 68 441 80 449
rect 98 441 110 449
rect 128 441 140 449
rect 158 441 170 449
rect 188 441 200 449
rect 218 441 230 449
rect 248 441 260 449
rect 278 441 290 449
rect 308 441 320 449
rect 338 441 350 449
rect 368 441 380 449
rect 398 441 410 449
rect 428 441 440 449
rect 458 441 470 449
rect 488 441 500 449
rect 518 441 530 449
rect 548 441 560 449
rect 568 441 572 449
rect 28 439 60 441
rect 68 439 90 441
rect 98 439 120 441
rect 128 439 150 441
rect 158 439 180 441
rect 188 439 210 441
rect 218 439 240 441
rect 248 439 270 441
rect 278 439 300 441
rect 308 439 330 441
rect 338 439 360 441
rect 368 439 390 441
rect 398 439 420 441
rect 428 439 450 441
rect 458 439 480 441
rect 488 439 510 441
rect 518 439 540 441
rect 548 439 572 441
rect 28 431 40 439
rect 48 431 60 439
rect 78 431 90 439
rect 108 431 120 439
rect 138 431 150 439
rect 168 431 180 439
rect 198 431 210 439
rect 228 431 240 439
rect 258 431 270 439
rect 288 431 300 439
rect 318 431 330 439
rect 348 431 360 439
rect 378 431 390 439
rect 408 431 420 439
rect 438 431 450 439
rect 468 431 480 439
rect 498 431 510 439
rect 528 431 540 439
rect 558 431 572 439
rect 28 429 60 431
rect 68 429 90 431
rect 98 429 120 431
rect 128 429 150 431
rect 158 429 180 431
rect 188 429 210 431
rect 218 429 240 431
rect 248 429 270 431
rect 278 429 300 431
rect 308 429 330 431
rect 338 429 360 431
rect 368 429 390 431
rect 398 429 420 431
rect 428 429 450 431
rect 458 429 480 431
rect 488 429 510 431
rect 518 429 540 431
rect 548 429 572 431
rect 28 421 30 429
rect 38 421 50 429
rect 68 421 80 429
rect 98 421 110 429
rect 128 421 140 429
rect 158 421 170 429
rect 188 421 200 429
rect 218 421 230 429
rect 248 421 260 429
rect 278 421 290 429
rect 308 421 320 429
rect 338 421 350 429
rect 368 421 380 429
rect 398 421 410 429
rect 428 421 440 429
rect 458 421 470 429
rect 488 421 500 429
rect 518 421 530 429
rect 548 421 560 429
rect 568 421 572 429
rect 28 419 60 421
rect 68 419 90 421
rect 98 419 120 421
rect 128 419 150 421
rect 158 419 180 421
rect 188 419 210 421
rect 218 419 240 421
rect 248 419 270 421
rect 278 419 300 421
rect 308 419 330 421
rect 338 419 360 421
rect 368 419 390 421
rect 398 419 420 421
rect 428 419 450 421
rect 458 419 480 421
rect 488 419 510 421
rect 518 419 540 421
rect 548 419 572 421
rect 28 411 40 419
rect 48 411 60 419
rect 78 411 90 419
rect 108 411 120 419
rect 138 411 150 419
rect 168 411 180 419
rect 198 411 210 419
rect 228 411 240 419
rect 258 411 270 419
rect 288 411 300 419
rect 318 411 330 419
rect 348 411 360 419
rect 378 411 390 419
rect 408 411 420 419
rect 438 411 450 419
rect 468 411 480 419
rect 498 411 510 419
rect 528 411 540 419
rect 558 411 572 419
rect 28 409 60 411
rect 68 409 90 411
rect 98 409 120 411
rect 128 409 150 411
rect 158 409 180 411
rect 188 409 210 411
rect 218 409 240 411
rect 248 409 270 411
rect 278 409 300 411
rect 308 409 330 411
rect 338 409 360 411
rect 368 409 390 411
rect 398 409 420 411
rect 428 409 450 411
rect 458 409 480 411
rect 488 409 510 411
rect 518 409 540 411
rect 548 409 572 411
rect 28 401 30 409
rect 38 401 50 409
rect 68 401 80 409
rect 98 401 110 409
rect 128 401 140 409
rect 158 401 170 409
rect 188 401 200 409
rect 218 401 230 409
rect 248 401 260 409
rect 278 401 290 409
rect 308 401 320 409
rect 338 401 350 409
rect 368 401 380 409
rect 398 401 410 409
rect 428 401 440 409
rect 458 401 470 409
rect 488 401 500 409
rect 518 401 530 409
rect 548 401 560 409
rect 568 401 572 409
rect 28 399 60 401
rect 68 399 90 401
rect 98 399 120 401
rect 128 399 150 401
rect 158 399 180 401
rect 188 399 210 401
rect 218 399 240 401
rect 248 399 270 401
rect 278 399 300 401
rect 308 399 330 401
rect 338 399 360 401
rect 368 399 390 401
rect 398 399 420 401
rect 428 399 450 401
rect 458 399 480 401
rect 488 399 510 401
rect 518 399 540 401
rect 548 399 572 401
rect 28 371 40 399
rect 48 371 60 399
rect 78 371 90 399
rect 108 391 120 399
rect 138 391 150 399
rect 168 391 180 399
rect 198 391 210 399
rect 228 391 240 399
rect 258 391 270 399
rect 288 391 300 399
rect 318 391 330 399
rect 348 391 360 399
rect 378 391 390 399
rect 408 391 420 399
rect 438 391 450 399
rect 468 391 480 399
rect 498 391 510 399
rect 528 391 540 399
rect 558 391 572 399
rect 98 379 510 391
rect 518 389 540 391
rect 548 389 572 391
rect 518 381 530 389
rect 548 381 560 389
rect 568 381 572 389
rect 518 379 540 381
rect 548 379 572 381
rect 108 371 120 379
rect 138 371 150 379
rect 168 371 180 379
rect 198 371 210 379
rect 228 371 240 379
rect 258 371 270 379
rect 288 371 300 379
rect 318 371 330 379
rect 348 371 360 379
rect 378 371 390 379
rect 408 371 420 379
rect 438 371 450 379
rect 468 371 480 379
rect 498 371 510 379
rect 528 371 540 379
rect 558 371 572 379
rect 28 369 60 371
rect 68 369 90 371
rect 98 369 120 371
rect 128 369 150 371
rect 158 369 180 371
rect 188 369 210 371
rect 218 369 240 371
rect 248 369 270 371
rect 278 369 300 371
rect 308 369 330 371
rect 338 369 360 371
rect 368 369 390 371
rect 398 369 420 371
rect 428 369 450 371
rect 458 369 480 371
rect 488 369 510 371
rect 518 369 540 371
rect 548 369 572 371
rect 28 361 30 369
rect 38 361 50 369
rect 68 361 80 369
rect 98 361 110 369
rect 128 361 140 369
rect 158 361 170 369
rect 188 361 200 369
rect 218 361 230 369
rect 248 361 260 369
rect 278 361 290 369
rect 308 361 320 369
rect 338 361 350 369
rect 368 361 380 369
rect 398 361 410 369
rect 428 361 440 369
rect 458 361 470 369
rect 488 361 500 369
rect 518 361 530 369
rect 548 361 560 369
rect 568 361 572 369
rect 28 359 60 361
rect 68 359 90 361
rect 98 359 120 361
rect 128 359 150 361
rect 158 359 180 361
rect 188 359 210 361
rect 218 359 240 361
rect 248 359 270 361
rect 278 359 300 361
rect 308 359 330 361
rect 338 359 360 361
rect 368 359 390 361
rect 398 359 420 361
rect 428 359 450 361
rect 458 359 480 361
rect 488 359 510 361
rect 518 359 540 361
rect 548 359 572 361
rect 28 351 40 359
rect 48 351 60 359
rect 78 351 90 359
rect 108 351 120 359
rect 138 351 150 359
rect 168 351 180 359
rect 198 351 210 359
rect 228 351 240 359
rect 258 351 270 359
rect 288 351 300 359
rect 318 351 330 359
rect 348 351 360 359
rect 378 351 390 359
rect 408 351 420 359
rect 438 351 450 359
rect 468 351 480 359
rect 498 351 510 359
rect 528 351 540 359
rect 558 351 572 359
rect 28 349 60 351
rect 68 349 90 351
rect 98 349 120 351
rect 128 349 150 351
rect 158 349 180 351
rect 188 349 210 351
rect 218 349 240 351
rect 248 349 270 351
rect 278 349 300 351
rect 308 349 330 351
rect 338 349 360 351
rect 368 349 390 351
rect 398 349 420 351
rect 428 349 450 351
rect 458 349 480 351
rect 488 349 510 351
rect 518 349 540 351
rect 548 349 572 351
rect 28 341 30 349
rect 38 341 50 349
rect 68 341 80 349
rect 98 341 110 349
rect 128 341 140 349
rect 158 341 170 349
rect 188 341 200 349
rect 218 341 230 349
rect 248 341 260 349
rect 278 341 290 349
rect 308 341 320 349
rect 338 341 350 349
rect 368 341 380 349
rect 398 341 410 349
rect 428 341 440 349
rect 458 341 470 349
rect 488 341 500 349
rect 518 341 530 349
rect 548 341 560 349
rect 568 341 572 349
rect 28 339 60 341
rect 68 339 90 341
rect 98 339 120 341
rect 128 339 150 341
rect 158 339 180 341
rect 188 339 210 341
rect 218 339 240 341
rect 248 339 270 341
rect 278 339 300 341
rect 308 339 330 341
rect 338 339 360 341
rect 368 339 390 341
rect 398 339 420 341
rect 428 339 450 341
rect 458 339 480 341
rect 488 339 510 341
rect 518 339 540 341
rect 548 339 572 341
rect 28 331 40 339
rect 48 331 60 339
rect 78 331 90 339
rect 108 331 120 339
rect 138 331 150 339
rect 168 331 180 339
rect 198 331 210 339
rect 228 331 240 339
rect 258 331 270 339
rect 288 331 300 339
rect 318 331 330 339
rect 348 331 360 339
rect 378 331 390 339
rect 408 331 420 339
rect 438 331 450 339
rect 468 331 480 339
rect 498 331 510 339
rect 528 331 540 339
rect 558 331 572 339
rect 28 329 60 331
rect 68 329 90 331
rect 98 329 120 331
rect 128 329 150 331
rect 158 329 180 331
rect 188 329 210 331
rect 218 329 240 331
rect 248 329 270 331
rect 278 329 300 331
rect 308 329 330 331
rect 338 329 360 331
rect 368 329 390 331
rect 398 329 420 331
rect 428 329 450 331
rect 458 329 480 331
rect 488 329 510 331
rect 518 329 540 331
rect 548 329 572 331
rect 28 321 30 329
rect 38 321 50 329
rect 68 321 80 329
rect 98 321 110 329
rect 128 321 140 329
rect 158 321 170 329
rect 188 321 200 329
rect 218 321 230 329
rect 248 321 260 329
rect 278 321 290 329
rect 308 321 320 329
rect 338 321 350 329
rect 368 321 380 329
rect 398 321 410 329
rect 428 321 440 329
rect 458 321 470 329
rect 488 321 500 329
rect 518 321 530 329
rect 548 321 560 329
rect 568 321 572 329
rect 28 319 60 321
rect 68 319 90 321
rect 98 319 120 321
rect 128 319 150 321
rect 158 319 180 321
rect 188 319 210 321
rect 218 319 240 321
rect 248 319 270 321
rect 278 319 300 321
rect 308 319 330 321
rect 338 319 360 321
rect 368 319 390 321
rect 398 319 420 321
rect 428 319 450 321
rect 458 319 480 321
rect 488 319 510 321
rect 518 319 540 321
rect 548 319 572 321
rect 28 311 40 319
rect 48 311 60 319
rect 78 311 90 319
rect 108 311 120 319
rect 138 311 150 319
rect 168 311 180 319
rect 198 311 210 319
rect 228 311 240 319
rect 258 311 270 319
rect 288 311 300 319
rect 318 311 330 319
rect 348 311 360 319
rect 378 311 390 319
rect 408 311 420 319
rect 438 311 450 319
rect 468 311 480 319
rect 498 311 510 319
rect 528 311 540 319
rect 558 311 572 319
rect 28 309 60 311
rect 68 309 510 311
rect 518 309 540 311
rect 548 309 572 311
rect 28 301 30 309
rect 38 301 50 309
rect 68 301 80 309
rect 88 301 500 309
rect 518 301 530 309
rect 548 301 560 309
rect 568 301 572 309
rect 28 299 60 301
rect 68 299 510 301
rect 518 299 540 301
rect 548 299 572 301
rect 28 291 40 299
rect 48 291 60 299
rect 78 291 90 299
rect 108 291 120 299
rect 138 291 150 299
rect 168 291 180 299
rect 198 291 210 299
rect 228 291 240 299
rect 258 291 270 299
rect 288 291 300 299
rect 318 291 330 299
rect 348 291 360 299
rect 378 291 390 299
rect 408 291 420 299
rect 438 291 450 299
rect 468 291 480 299
rect 498 291 510 299
rect 528 291 540 299
rect 558 291 572 299
rect 28 289 60 291
rect 68 289 90 291
rect 98 289 120 291
rect 128 289 150 291
rect 158 289 180 291
rect 188 289 210 291
rect 218 289 240 291
rect 248 289 270 291
rect 278 289 300 291
rect 308 289 330 291
rect 338 289 360 291
rect 368 289 390 291
rect 398 289 420 291
rect 428 289 450 291
rect 458 289 480 291
rect 488 289 510 291
rect 518 289 540 291
rect 548 289 572 291
rect 28 281 30 289
rect 38 281 50 289
rect 68 281 80 289
rect 98 281 110 289
rect 128 281 140 289
rect 158 281 170 289
rect 188 281 200 289
rect 218 281 230 289
rect 248 281 260 289
rect 278 281 290 289
rect 308 281 320 289
rect 338 281 350 289
rect 368 281 380 289
rect 398 281 410 289
rect 428 281 440 289
rect 458 281 470 289
rect 488 281 500 289
rect 518 281 530 289
rect 548 281 560 289
rect 568 281 572 289
rect 28 279 60 281
rect 68 279 90 281
rect 98 279 120 281
rect 128 279 150 281
rect 158 279 180 281
rect 188 279 210 281
rect 218 279 240 281
rect 248 279 270 281
rect 278 279 300 281
rect 308 279 330 281
rect 338 279 360 281
rect 368 279 390 281
rect 398 279 420 281
rect 428 279 450 281
rect 458 279 480 281
rect 488 279 510 281
rect 518 279 540 281
rect 548 279 572 281
rect 28 271 40 279
rect 48 271 60 279
rect 78 271 90 279
rect 108 271 120 279
rect 138 271 150 279
rect 168 271 180 279
rect 198 271 210 279
rect 228 271 240 279
rect 258 271 270 279
rect 288 271 300 279
rect 318 271 330 279
rect 348 271 360 279
rect 378 271 390 279
rect 408 271 420 279
rect 438 271 450 279
rect 468 271 480 279
rect 498 271 510 279
rect 528 271 540 279
rect 558 271 572 279
rect 28 269 60 271
rect 68 269 90 271
rect 98 269 120 271
rect 128 269 150 271
rect 158 269 180 271
rect 188 269 210 271
rect 218 269 240 271
rect 248 269 270 271
rect 278 269 300 271
rect 308 269 330 271
rect 338 269 360 271
rect 368 269 390 271
rect 398 269 420 271
rect 428 269 450 271
rect 458 269 480 271
rect 488 269 510 271
rect 518 269 540 271
rect 548 269 572 271
rect 28 261 30 269
rect 38 261 50 269
rect 68 261 80 269
rect 98 261 110 269
rect 128 261 140 269
rect 158 261 170 269
rect 188 261 200 269
rect 218 261 230 269
rect 248 261 260 269
rect 278 261 290 269
rect 308 261 320 269
rect 338 261 350 269
rect 368 261 380 269
rect 398 261 410 269
rect 428 261 440 269
rect 458 261 470 269
rect 488 261 500 269
rect 518 261 530 269
rect 548 261 560 269
rect 568 261 572 269
rect 28 259 60 261
rect 68 259 90 261
rect 98 259 120 261
rect 128 259 150 261
rect 158 259 180 261
rect 188 259 210 261
rect 218 259 240 261
rect 248 259 270 261
rect 278 259 300 261
rect 308 259 330 261
rect 338 259 360 261
rect 368 259 390 261
rect 398 259 420 261
rect 428 259 450 261
rect 458 259 480 261
rect 488 259 510 261
rect 518 259 540 261
rect 548 259 572 261
rect 28 251 40 259
rect 48 251 60 259
rect 78 251 90 259
rect 108 251 120 259
rect 138 251 150 259
rect 168 251 180 259
rect 198 251 210 259
rect 228 251 240 259
rect 258 251 270 259
rect 288 251 300 259
rect 318 251 330 259
rect 348 251 360 259
rect 378 251 390 259
rect 408 251 420 259
rect 438 251 450 259
rect 468 251 480 259
rect 498 251 510 259
rect 528 251 540 259
rect 558 251 572 259
rect 28 249 60 251
rect 68 249 90 251
rect 98 249 120 251
rect 128 249 150 251
rect 158 249 180 251
rect 188 249 210 251
rect 218 249 240 251
rect 248 249 270 251
rect 278 249 300 251
rect 308 249 330 251
rect 338 249 360 251
rect 368 249 390 251
rect 398 249 420 251
rect 428 249 450 251
rect 458 249 480 251
rect 488 249 510 251
rect 518 249 540 251
rect 548 249 572 251
rect 28 241 30 249
rect 38 241 50 249
rect 28 239 60 241
rect 28 231 40 239
rect 48 231 60 239
rect 28 229 60 231
rect 28 221 30 229
rect 38 221 50 229
rect 68 221 80 249
rect 98 241 110 249
rect 128 241 140 249
rect 158 241 170 249
rect 188 241 200 249
rect 218 241 230 249
rect 248 241 260 249
rect 278 241 290 249
rect 308 241 320 249
rect 338 241 350 249
rect 368 241 380 249
rect 398 241 410 249
rect 428 241 440 249
rect 458 241 470 249
rect 488 241 500 249
rect 518 241 530 249
rect 548 241 560 249
rect 568 241 572 249
rect 88 229 500 241
rect 508 239 540 241
rect 548 239 572 241
rect 508 231 520 239
rect 528 231 540 239
rect 558 231 572 239
rect 508 229 540 231
rect 548 229 572 231
rect 98 221 110 229
rect 128 221 140 229
rect 158 221 170 229
rect 188 221 200 229
rect 218 221 230 229
rect 248 221 260 229
rect 278 221 290 229
rect 308 221 320 229
rect 338 221 350 229
rect 368 221 380 229
rect 398 221 410 229
rect 428 221 440 229
rect 458 221 470 229
rect 488 221 500 229
rect 518 221 530 229
rect 548 221 560 229
rect 568 221 572 229
rect 28 219 60 221
rect 68 219 90 221
rect 98 219 120 221
rect 128 219 150 221
rect 158 219 180 221
rect 188 219 210 221
rect 218 219 240 221
rect 248 219 270 221
rect 278 219 300 221
rect 308 219 330 221
rect 338 219 360 221
rect 368 219 390 221
rect 398 219 420 221
rect 428 219 450 221
rect 458 219 480 221
rect 488 219 510 221
rect 518 219 540 221
rect 548 219 572 221
rect 28 211 40 219
rect 48 211 60 219
rect 78 211 90 219
rect 108 211 120 219
rect 138 211 150 219
rect 168 211 180 219
rect 198 211 210 219
rect 228 211 240 219
rect 258 211 270 219
rect 288 211 300 219
rect 318 211 330 219
rect 348 211 360 219
rect 378 211 390 219
rect 408 211 420 219
rect 438 211 450 219
rect 468 211 480 219
rect 498 211 510 219
rect 528 211 540 219
rect 558 211 572 219
rect 28 209 60 211
rect 68 209 90 211
rect 98 209 120 211
rect 128 209 150 211
rect 158 209 180 211
rect 188 209 210 211
rect 218 209 240 211
rect 248 209 270 211
rect 278 209 300 211
rect 308 209 330 211
rect 338 209 360 211
rect 368 209 390 211
rect 398 209 420 211
rect 428 209 450 211
rect 458 209 480 211
rect 488 209 510 211
rect 518 209 540 211
rect 548 209 572 211
rect 28 201 30 209
rect 38 201 50 209
rect 68 201 80 209
rect 98 201 110 209
rect 128 201 140 209
rect 158 201 170 209
rect 188 201 200 209
rect 218 201 230 209
rect 248 201 260 209
rect 278 201 290 209
rect 308 201 320 209
rect 338 201 350 209
rect 368 201 380 209
rect 398 201 410 209
rect 428 201 440 209
rect 458 201 470 209
rect 488 201 500 209
rect 518 201 530 209
rect 548 201 560 209
rect 568 201 572 209
rect 28 199 60 201
rect 68 199 90 201
rect 98 199 120 201
rect 128 199 150 201
rect 158 199 180 201
rect 188 199 210 201
rect 218 199 240 201
rect 248 199 270 201
rect 278 199 300 201
rect 308 199 330 201
rect 338 199 360 201
rect 368 199 390 201
rect 398 199 420 201
rect 428 199 450 201
rect 458 199 480 201
rect 488 199 510 201
rect 518 199 540 201
rect 548 199 572 201
rect 28 191 40 199
rect 48 191 60 199
rect 78 191 90 199
rect 108 191 120 199
rect 138 191 150 199
rect 168 191 180 199
rect 198 191 210 199
rect 228 191 240 199
rect 258 191 270 199
rect 288 191 300 199
rect 318 191 330 199
rect 348 191 360 199
rect 378 191 390 199
rect 408 191 420 199
rect 438 191 450 199
rect 468 191 480 199
rect 498 191 510 199
rect 528 191 540 199
rect 558 191 572 199
rect 28 189 60 191
rect 68 189 90 191
rect 98 189 120 191
rect 128 189 150 191
rect 158 189 180 191
rect 188 189 210 191
rect 218 189 240 191
rect 248 189 270 191
rect 278 189 300 191
rect 308 189 330 191
rect 338 189 360 191
rect 368 189 390 191
rect 398 189 420 191
rect 428 189 450 191
rect 458 189 480 191
rect 488 189 510 191
rect 518 189 540 191
rect 548 189 572 191
rect 28 181 30 189
rect 38 181 50 189
rect 68 181 80 189
rect 98 181 110 189
rect 128 181 140 189
rect 158 181 170 189
rect 188 181 200 189
rect 218 181 230 189
rect 248 181 260 189
rect 278 181 290 189
rect 308 181 320 189
rect 338 181 350 189
rect 368 181 380 189
rect 398 181 410 189
rect 428 181 440 189
rect 458 181 470 189
rect 488 181 500 189
rect 518 181 530 189
rect 548 181 560 189
rect 568 181 572 189
rect 28 179 60 181
rect 68 179 90 181
rect 98 179 120 181
rect 128 179 150 181
rect 158 179 180 181
rect 188 179 210 181
rect 218 179 240 181
rect 248 179 270 181
rect 278 179 300 181
rect 308 179 330 181
rect 338 179 360 181
rect 368 179 390 181
rect 398 179 420 181
rect 428 179 450 181
rect 458 179 480 181
rect 488 179 510 181
rect 518 179 540 181
rect 548 179 572 181
rect 28 171 40 179
rect 48 171 60 179
rect 78 171 90 179
rect 108 171 120 179
rect 138 171 150 179
rect 168 171 180 179
rect 198 171 210 179
rect 228 171 240 179
rect 258 171 270 179
rect 288 171 300 179
rect 318 171 330 179
rect 348 171 360 179
rect 378 171 390 179
rect 408 171 420 179
rect 438 171 450 179
rect 468 171 480 179
rect 498 171 510 179
rect 528 171 540 179
rect 558 171 572 179
rect 28 169 60 171
rect 68 169 90 171
rect 98 169 120 171
rect 128 169 150 171
rect 158 169 180 171
rect 188 169 210 171
rect 218 169 240 171
rect 248 169 270 171
rect 278 169 300 171
rect 308 169 330 171
rect 338 169 360 171
rect 368 169 390 171
rect 398 169 420 171
rect 428 169 450 171
rect 458 169 480 171
rect 488 169 510 171
rect 518 169 540 171
rect 548 169 572 171
rect 28 161 30 169
rect 38 161 50 169
rect 68 161 80 169
rect 98 161 110 169
rect 128 161 140 169
rect 158 161 170 169
rect 188 161 200 169
rect 218 161 230 169
rect 248 161 260 169
rect 278 161 290 169
rect 308 161 320 169
rect 338 161 350 169
rect 368 161 380 169
rect 398 161 410 169
rect 428 161 440 169
rect 458 161 470 169
rect 488 161 500 169
rect 518 161 530 169
rect 548 161 560 169
rect 568 161 572 169
rect 28 159 60 161
rect 68 159 90 161
rect 28 151 40 159
rect 48 151 60 159
rect 78 151 90 159
rect 28 149 60 151
rect 68 149 90 151
rect 98 149 500 161
rect 508 159 540 161
rect 548 159 572 161
rect 508 151 520 159
rect 528 151 540 159
rect 558 151 572 159
rect 508 149 540 151
rect 548 149 572 151
rect 28 141 30 149
rect 38 141 50 149
rect 68 141 80 149
rect 98 141 110 149
rect 128 141 140 149
rect 158 141 170 149
rect 188 141 200 149
rect 218 141 230 149
rect 248 141 260 149
rect 278 141 290 149
rect 308 141 320 149
rect 338 141 350 149
rect 368 141 380 149
rect 398 141 410 149
rect 428 141 440 149
rect 458 141 470 149
rect 488 141 500 149
rect 518 141 530 149
rect 548 141 560 149
rect 568 141 572 149
rect 28 139 60 141
rect 68 139 90 141
rect 98 139 120 141
rect 128 139 150 141
rect 158 139 180 141
rect 188 139 210 141
rect 218 139 240 141
rect 248 139 270 141
rect 278 139 300 141
rect 308 139 330 141
rect 338 139 360 141
rect 368 139 390 141
rect 398 139 420 141
rect 428 139 450 141
rect 458 139 480 141
rect 488 139 510 141
rect 518 139 540 141
rect 548 139 572 141
rect 28 131 40 139
rect 48 131 60 139
rect 78 131 90 139
rect 108 131 120 139
rect 138 131 150 139
rect 168 131 180 139
rect 198 131 210 139
rect 228 131 240 139
rect 258 131 270 139
rect 288 131 300 139
rect 318 131 330 139
rect 348 131 360 139
rect 378 131 390 139
rect 408 131 420 139
rect 438 131 450 139
rect 468 131 480 139
rect 498 131 510 139
rect 528 131 540 139
rect 558 131 572 139
rect 28 129 60 131
rect 68 129 90 131
rect 98 129 120 131
rect 128 129 150 131
rect 158 129 180 131
rect 188 129 210 131
rect 218 129 240 131
rect 248 129 270 131
rect 278 129 300 131
rect 308 129 330 131
rect 338 129 360 131
rect 368 129 390 131
rect 398 129 420 131
rect 428 129 450 131
rect 458 129 480 131
rect 488 129 510 131
rect 518 129 540 131
rect 548 129 572 131
rect 28 121 30 129
rect 38 121 50 129
rect 68 121 80 129
rect 98 121 110 129
rect 128 121 140 129
rect 158 121 170 129
rect 188 121 200 129
rect 218 121 230 129
rect 248 121 260 129
rect 278 121 290 129
rect 308 121 320 129
rect 338 121 350 129
rect 368 121 380 129
rect 398 121 410 129
rect 428 121 440 129
rect 458 121 470 129
rect 488 121 500 129
rect 518 121 530 129
rect 548 121 560 129
rect 568 121 572 129
rect 28 119 60 121
rect 68 119 90 121
rect 98 119 120 121
rect 128 119 150 121
rect 158 119 180 121
rect 188 119 210 121
rect 218 119 240 121
rect 248 119 270 121
rect 278 119 300 121
rect 308 119 330 121
rect 338 119 360 121
rect 368 119 390 121
rect 398 119 420 121
rect 428 119 450 121
rect 458 119 480 121
rect 488 119 510 121
rect 518 119 540 121
rect 548 119 572 121
rect 28 111 40 119
rect 48 111 60 119
rect 78 111 90 119
rect 108 111 120 119
rect 138 111 150 119
rect 168 111 180 119
rect 198 111 210 119
rect 228 111 240 119
rect 258 111 270 119
rect 288 111 300 119
rect 318 111 330 119
rect 348 111 360 119
rect 378 111 390 119
rect 408 111 420 119
rect 438 111 450 119
rect 468 111 480 119
rect 498 111 510 119
rect 528 111 540 119
rect 558 111 572 119
rect 28 109 60 111
rect 68 109 90 111
rect 98 109 120 111
rect 128 109 150 111
rect 158 109 180 111
rect 188 109 210 111
rect 218 109 240 111
rect 248 109 270 111
rect 278 109 300 111
rect 308 109 330 111
rect 338 109 360 111
rect 368 109 390 111
rect 398 109 420 111
rect 428 109 450 111
rect 458 109 480 111
rect 488 109 510 111
rect 518 109 540 111
rect 548 109 572 111
rect 28 101 30 109
rect 38 101 50 109
rect 68 101 80 109
rect 98 101 110 109
rect 128 101 140 109
rect 158 101 170 109
rect 188 101 200 109
rect 218 101 230 109
rect 248 101 260 109
rect 278 101 290 109
rect 308 101 320 109
rect 338 101 350 109
rect 368 101 380 109
rect 398 101 410 109
rect 428 101 440 109
rect 458 101 470 109
rect 488 101 500 109
rect 518 101 530 109
rect 548 101 560 109
rect 568 101 572 109
rect 28 99 60 101
rect 68 99 90 101
rect 98 99 120 101
rect 128 99 150 101
rect 158 99 180 101
rect 188 99 210 101
rect 218 99 240 101
rect 248 99 270 101
rect 278 99 300 101
rect 308 99 330 101
rect 338 99 360 101
rect 368 99 390 101
rect 398 99 420 101
rect 428 99 450 101
rect 458 99 480 101
rect 488 99 510 101
rect 518 99 540 101
rect 548 99 572 101
rect 28 91 40 99
rect 48 91 60 99
rect 78 91 90 99
rect 108 91 120 99
rect 138 91 150 99
rect 168 91 180 99
rect 198 91 210 99
rect 228 91 240 99
rect 258 91 270 99
rect 288 91 300 99
rect 318 91 330 99
rect 348 91 360 99
rect 378 91 390 99
rect 408 91 420 99
rect 438 91 450 99
rect 468 91 480 99
rect 498 91 510 99
rect 528 91 540 99
rect 558 91 572 99
rect 28 89 60 91
rect 68 89 90 91
rect 98 89 120 91
rect 128 89 150 91
rect 158 89 180 91
rect 188 89 210 91
rect 218 89 240 91
rect 248 89 270 91
rect 278 89 300 91
rect 308 89 330 91
rect 338 89 360 91
rect 368 89 390 91
rect 398 89 420 91
rect 428 89 450 91
rect 458 89 480 91
rect 488 89 510 91
rect 518 89 540 91
rect 548 89 572 91
rect 28 81 30 89
rect 38 81 50 89
rect 68 81 80 89
rect 98 81 110 89
rect 128 81 140 89
rect 158 81 170 89
rect 188 81 200 89
rect 218 81 230 89
rect 248 81 260 89
rect 278 81 290 89
rect 308 81 320 89
rect 338 81 350 89
rect 368 81 380 89
rect 398 81 410 89
rect 428 81 440 89
rect 458 81 470 89
rect 488 81 500 89
rect 518 81 530 89
rect 548 81 560 89
rect 568 81 572 89
rect 28 79 60 81
rect 68 79 90 81
rect 98 79 120 81
rect 128 79 150 81
rect 158 79 180 81
rect 188 79 210 81
rect 218 79 240 81
rect 248 79 270 81
rect 278 79 300 81
rect 308 79 330 81
rect 338 79 360 81
rect 368 79 390 81
rect 398 79 420 81
rect 428 79 450 81
rect 458 79 480 81
rect 488 79 510 81
rect 518 79 540 81
rect 548 79 572 81
rect 28 71 40 79
rect 48 71 60 79
rect 78 71 90 79
rect 108 71 120 79
rect 138 71 150 79
rect 168 71 180 79
rect 198 71 210 79
rect 228 71 240 79
rect 258 71 270 79
rect 288 71 300 79
rect 318 71 330 79
rect 348 71 360 79
rect 378 71 390 79
rect 408 71 420 79
rect 438 71 450 79
rect 468 71 480 79
rect 498 71 510 79
rect 528 71 540 79
rect 558 71 572 79
rect 28 69 60 71
rect 68 69 90 71
rect 98 69 120 71
rect 128 69 150 71
rect 158 69 180 71
rect 188 69 210 71
rect 218 69 240 71
rect 248 69 270 71
rect 278 69 300 71
rect 308 69 330 71
rect 338 69 360 71
rect 368 69 390 71
rect 398 69 420 71
rect 428 69 450 71
rect 458 69 480 71
rect 488 69 510 71
rect 518 69 540 71
rect 548 69 572 71
rect 28 61 30 69
rect 38 61 50 69
rect 68 61 80 69
rect 98 61 110 69
rect 128 61 140 69
rect 158 61 170 69
rect 188 61 200 69
rect 218 61 230 69
rect 248 61 260 69
rect 278 61 290 69
rect 308 61 320 69
rect 338 61 350 69
rect 368 61 380 69
rect 398 61 410 69
rect 428 61 440 69
rect 458 61 470 69
rect 488 61 500 69
rect 518 61 530 69
rect 548 61 560 69
rect 568 61 572 69
rect 28 59 60 61
rect 68 59 90 61
rect 98 59 120 61
rect 128 59 150 61
rect 158 59 180 61
rect 188 59 210 61
rect 218 59 240 61
rect 248 59 270 61
rect 278 59 300 61
rect 308 59 330 61
rect 338 59 360 61
rect 368 59 390 61
rect 398 59 420 61
rect 428 59 450 61
rect 458 59 480 61
rect 488 59 510 61
rect 518 59 540 61
rect 548 59 572 61
rect 28 51 40 59
rect 48 51 60 59
rect 78 51 90 59
rect 108 51 120 59
rect 138 51 150 59
rect 168 51 180 59
rect 198 51 210 59
rect 228 51 240 59
rect 258 51 270 59
rect 288 51 300 59
rect 318 51 330 59
rect 348 51 360 59
rect 378 51 390 59
rect 408 51 420 59
rect 438 51 450 59
rect 468 51 480 59
rect 498 51 510 59
rect 528 51 540 59
rect 558 51 572 59
rect 28 49 60 51
rect 68 49 90 51
rect 98 49 120 51
rect 128 49 150 51
rect 158 49 180 51
rect 188 49 210 51
rect 218 49 240 51
rect 248 49 270 51
rect 278 49 300 51
rect 308 49 330 51
rect 338 49 360 51
rect 368 49 390 51
rect 398 49 420 51
rect 428 49 450 51
rect 458 49 480 51
rect 488 49 510 51
rect 518 49 540 51
rect 548 49 572 51
rect 28 41 30 49
rect 38 41 50 49
rect 68 41 80 49
rect 98 41 110 49
rect 128 41 140 49
rect 158 41 170 49
rect 188 41 200 49
rect 218 41 230 49
rect 248 41 260 49
rect 278 41 290 49
rect 308 41 320 49
rect 338 41 350 49
rect 368 41 380 49
rect 398 41 410 49
rect 428 41 440 49
rect 458 41 470 49
rect 488 41 500 49
rect 518 41 530 49
rect 548 41 560 49
rect 568 41 572 49
rect 28 39 60 41
rect 68 39 90 41
rect 98 39 120 41
rect 128 39 150 41
rect 158 39 180 41
rect 188 39 210 41
rect 218 39 240 41
rect 248 39 270 41
rect 278 39 300 41
rect 308 39 330 41
rect 338 39 360 41
rect 368 39 390 41
rect 398 39 420 41
rect 428 39 450 41
rect 458 39 480 41
rect 488 39 510 41
rect 518 39 540 41
rect 548 39 572 41
rect 28 31 40 39
rect 48 31 60 39
rect 78 31 90 39
rect 108 31 120 39
rect 138 31 150 39
rect 168 31 180 39
rect 198 31 210 39
rect 228 31 240 39
rect 258 31 270 39
rect 288 31 300 39
rect 318 31 330 39
rect 348 31 360 39
rect 378 31 390 39
rect 408 31 420 39
rect 438 31 450 39
rect 468 31 480 39
rect 498 31 510 39
rect 528 31 540 39
rect 558 31 572 39
rect 28 28 572 31
<< nsubstratendiff >>
rect 40 1298 560 1300
rect 40 1290 51 1298
rect 59 1290 72 1298
rect 80 1294 520 1298
rect 40 1289 82 1290
rect 40 1288 62 1289
rect 40 1280 41 1288
rect 49 1281 62 1288
rect 70 1286 82 1289
rect 90 1286 102 1294
rect 110 1286 122 1294
rect 130 1286 142 1294
rect 150 1286 162 1294
rect 170 1286 182 1294
rect 190 1286 202 1294
rect 210 1286 222 1294
rect 230 1286 370 1294
rect 378 1286 390 1294
rect 398 1286 410 1294
rect 418 1286 430 1294
rect 438 1286 450 1294
rect 458 1286 470 1294
rect 478 1286 490 1294
rect 498 1286 510 1294
rect 528 1290 541 1298
rect 549 1290 560 1298
rect 518 1289 560 1290
rect 518 1286 530 1289
rect 70 1284 530 1286
rect 70 1281 92 1284
rect 49 1280 92 1281
rect 40 1278 60 1280
rect 40 1270 51 1278
rect 59 1270 60 1278
rect 40 1268 60 1270
rect 40 1260 41 1268
rect 49 1260 60 1268
rect 40 1258 60 1260
rect 76 1276 92 1280
rect 100 1276 112 1284
rect 120 1276 132 1284
rect 140 1276 152 1284
rect 160 1276 172 1284
rect 180 1276 192 1284
rect 200 1276 212 1284
rect 220 1276 232 1284
rect 240 1280 360 1284
rect 240 1276 276 1280
rect 40 1250 51 1258
rect 59 1250 60 1258
rect 40 1248 60 1250
rect 40 1240 41 1248
rect 49 1240 60 1248
rect 40 1238 60 1240
rect 40 1230 51 1238
rect 59 1230 60 1238
rect 40 1228 60 1230
rect 40 1220 41 1228
rect 49 1220 60 1228
rect 40 1218 60 1220
rect 40 1210 51 1218
rect 59 1210 60 1218
rect 40 1208 60 1210
rect 40 1200 41 1208
rect 49 1200 60 1208
rect 40 1198 60 1200
rect 40 1190 51 1198
rect 59 1190 60 1198
rect 40 1188 60 1190
rect 40 1180 41 1188
rect 49 1180 60 1188
rect 40 1178 60 1180
rect 40 1170 51 1178
rect 59 1170 60 1178
rect 40 1168 60 1170
rect 40 1160 41 1168
rect 49 1160 60 1168
rect 40 1158 60 1160
rect 40 1150 51 1158
rect 59 1150 60 1158
rect 40 1148 60 1150
rect 40 1140 41 1148
rect 49 1140 60 1148
rect 40 1138 60 1140
rect 40 1130 51 1138
rect 59 1130 60 1138
rect 40 1128 60 1130
rect 40 1120 41 1128
rect 49 1120 60 1128
rect 40 1118 60 1120
rect 40 1110 51 1118
rect 59 1110 60 1118
rect 40 1108 60 1110
rect 40 1100 41 1108
rect 49 1100 60 1108
rect 40 1098 60 1100
rect 40 1090 51 1098
rect 59 1090 60 1098
rect 40 1088 60 1090
rect 40 1080 41 1088
rect 49 1080 60 1088
rect 40 1078 60 1080
rect 40 1070 51 1078
rect 59 1070 60 1078
rect 40 1068 60 1070
rect 40 1060 41 1068
rect 49 1060 60 1068
rect 40 1058 60 1060
rect 40 1050 51 1058
rect 59 1050 60 1058
rect 40 1048 60 1050
rect 40 1040 41 1048
rect 49 1040 60 1048
rect 40 1038 60 1040
rect 40 1030 51 1038
rect 59 1030 60 1038
rect 40 1028 60 1030
rect 40 1020 41 1028
rect 49 1020 60 1028
rect 40 1018 60 1020
rect 40 1010 51 1018
rect 59 1010 60 1018
rect 40 1008 60 1010
rect 40 1000 41 1008
rect 49 1000 60 1008
rect 40 998 60 1000
rect 40 990 51 998
rect 59 990 60 998
rect 40 988 60 990
rect 40 980 41 988
rect 49 980 60 988
rect 40 978 60 980
rect 40 970 51 978
rect 59 970 60 978
rect 40 968 60 970
rect 40 960 41 968
rect 49 960 60 968
rect 40 958 60 960
rect 40 950 51 958
rect 59 950 60 958
rect 40 948 60 950
rect 40 940 41 948
rect 49 940 60 948
rect 40 938 60 940
rect 40 930 51 938
rect 59 930 60 938
rect 40 928 60 930
rect 40 920 41 928
rect 49 920 60 928
rect 40 918 60 920
rect 40 910 51 918
rect 59 910 60 918
rect 40 908 60 910
rect 40 900 41 908
rect 49 900 60 908
rect 284 1230 316 1280
rect 324 1276 360 1280
rect 368 1276 380 1284
rect 388 1276 400 1284
rect 408 1276 420 1284
rect 428 1276 440 1284
rect 448 1276 460 1284
rect 468 1276 480 1284
rect 488 1276 500 1284
rect 508 1281 530 1284
rect 538 1288 560 1289
rect 538 1281 551 1288
rect 508 1280 551 1281
rect 559 1280 560 1288
rect 508 1276 524 1280
rect 540 1278 560 1280
rect 540 1270 541 1278
rect 549 1270 560 1278
rect 540 1268 560 1270
rect 540 1260 551 1268
rect 559 1260 560 1268
rect 540 1258 560 1260
rect 284 1222 286 1230
rect 314 1222 316 1230
rect 284 1210 316 1222
rect 284 1202 286 1210
rect 314 1202 316 1210
rect 284 1190 316 1202
rect 284 1182 286 1190
rect 314 1182 316 1190
rect 284 1102 316 1182
rect 284 1094 286 1102
rect 314 1094 316 1102
rect 284 1082 316 1094
rect 284 1074 286 1082
rect 314 1074 316 1082
rect 284 1062 316 1074
rect 284 1054 286 1062
rect 314 1054 316 1062
rect 284 972 316 1054
rect 284 964 286 972
rect 314 964 316 972
rect 284 952 316 964
rect 284 944 286 952
rect 314 944 316 952
rect 284 932 316 944
rect 284 924 286 932
rect 314 924 316 932
rect 40 898 60 900
rect 40 890 51 898
rect 59 890 60 898
rect 40 888 60 890
rect 40 880 41 888
rect 49 884 60 888
rect 76 884 276 888
rect 284 884 316 924
rect 540 1250 541 1258
rect 549 1250 560 1258
rect 540 1248 560 1250
rect 540 1240 551 1248
rect 559 1240 560 1248
rect 540 1238 560 1240
rect 540 1230 541 1238
rect 549 1230 560 1238
rect 540 1228 560 1230
rect 540 1220 551 1228
rect 559 1220 560 1228
rect 540 1218 560 1220
rect 540 1210 541 1218
rect 549 1210 560 1218
rect 540 1208 560 1210
rect 540 1200 551 1208
rect 559 1200 560 1208
rect 540 1198 560 1200
rect 540 1190 541 1198
rect 549 1190 560 1198
rect 540 1188 560 1190
rect 540 1180 551 1188
rect 559 1180 560 1188
rect 540 1178 560 1180
rect 540 1170 541 1178
rect 549 1170 560 1178
rect 540 1168 560 1170
rect 540 1160 551 1168
rect 559 1160 560 1168
rect 540 1158 560 1160
rect 540 1150 541 1158
rect 549 1150 560 1158
rect 540 1148 560 1150
rect 540 1140 551 1148
rect 559 1140 560 1148
rect 540 1138 560 1140
rect 540 1130 541 1138
rect 549 1130 560 1138
rect 540 1128 560 1130
rect 540 1120 551 1128
rect 559 1120 560 1128
rect 540 1118 560 1120
rect 540 1110 541 1118
rect 549 1110 560 1118
rect 540 1108 560 1110
rect 540 1100 551 1108
rect 559 1100 560 1108
rect 540 1098 560 1100
rect 540 1090 541 1098
rect 549 1090 560 1098
rect 540 1088 560 1090
rect 540 1080 551 1088
rect 559 1080 560 1088
rect 540 1078 560 1080
rect 540 1070 541 1078
rect 549 1070 560 1078
rect 540 1068 560 1070
rect 540 1060 551 1068
rect 559 1060 560 1068
rect 540 1058 560 1060
rect 540 1050 541 1058
rect 549 1050 560 1058
rect 540 1048 560 1050
rect 540 1040 551 1048
rect 559 1040 560 1048
rect 540 1038 560 1040
rect 540 1030 541 1038
rect 549 1030 560 1038
rect 540 1028 560 1030
rect 540 1020 551 1028
rect 559 1020 560 1028
rect 540 1018 560 1020
rect 540 1010 541 1018
rect 549 1010 560 1018
rect 540 1008 560 1010
rect 540 1000 551 1008
rect 559 1000 560 1008
rect 540 998 560 1000
rect 540 990 541 998
rect 549 990 560 998
rect 540 988 560 990
rect 540 980 551 988
rect 559 980 560 988
rect 540 978 560 980
rect 540 970 541 978
rect 549 970 560 978
rect 540 968 560 970
rect 540 960 551 968
rect 559 960 560 968
rect 540 958 560 960
rect 540 950 541 958
rect 549 950 560 958
rect 540 948 560 950
rect 540 940 551 948
rect 559 940 560 948
rect 540 938 560 940
rect 540 930 541 938
rect 549 930 560 938
rect 540 928 560 930
rect 540 920 551 928
rect 559 920 560 928
rect 540 918 560 920
rect 540 910 541 918
rect 549 910 560 918
rect 540 908 560 910
rect 324 884 524 888
rect 540 900 551 908
rect 559 900 560 908
rect 540 898 560 900
rect 540 890 541 898
rect 549 890 560 898
rect 540 888 560 890
rect 540 884 551 888
rect 49 883 551 884
rect 49 880 62 883
rect 40 873 62 880
rect 40 865 42 873
rect 240 865 360 883
rect 538 880 551 883
rect 559 880 560 888
rect 538 873 560 880
rect 558 865 560 873
rect 40 864 560 865
rect 0 652 600 654
rect 0 644 4 652
rect 12 644 24 652
rect 42 644 54 652
rect 72 644 84 652
rect 102 644 114 652
rect 132 644 144 652
rect 162 644 174 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 0 634 14 642
rect 22 634 34 642
rect 52 634 64 642
rect 82 634 94 642
rect 112 634 124 642
rect 142 634 154 642
rect 172 634 184 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 192 642 408 652
rect 426 644 438 652
rect 456 644 468 652
rect 486 644 498 652
rect 516 644 528 652
rect 546 644 558 652
rect 576 644 588 652
rect 596 644 600 652
rect 192 634 286 642
rect 314 634 408 642
rect 0 624 4 632
rect 12 624 24 632
rect 42 624 54 632
rect 72 624 84 632
rect 102 624 114 632
rect 132 624 144 632
rect 162 624 174 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 0 614 14 622
rect 22 614 34 622
rect 52 614 64 622
rect 82 614 94 622
rect 112 614 124 622
rect 142 614 154 622
rect 172 614 184 622
rect 192 622 408 634
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 416 634 428 642
rect 446 634 458 642
rect 476 634 488 642
rect 506 634 518 642
rect 536 634 548 642
rect 566 634 578 642
rect 586 634 600 642
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 426 624 438 632
rect 456 624 468 632
rect 486 624 498 632
rect 516 624 528 632
rect 546 624 558 632
rect 576 624 588 632
rect 596 624 600 632
rect 192 614 286 622
rect 314 614 408 622
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 416 614 428 622
rect 446 614 458 622
rect 476 614 488 622
rect 506 614 518 622
rect 536 614 548 622
rect 566 614 578 622
rect 586 614 600 622
rect 0 612 600 614
rect 0 604 4 612
rect 12 604 24 612
rect 32 604 568 612
rect 576 604 588 612
rect 596 604 600 612
rect 0 602 600 604
rect 0 594 14 602
rect 22 594 34 602
rect 52 594 64 602
rect 82 594 94 602
rect 112 594 124 602
rect 142 594 154 602
rect 172 594 184 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 192 594 286 602
rect 314 594 408 602
rect 0 584 4 592
rect 12 584 24 592
rect 42 584 54 592
rect 72 584 84 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 592
rect 132 582 144 592
rect 162 582 174 592
rect 192 584 408 594
rect 416 594 428 602
rect 446 594 458 602
rect 476 594 488 602
rect 506 594 518 602
rect 536 594 548 602
rect 566 594 578 602
rect 586 594 600 602
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 0 574 14 582
rect 22 574 34 582
rect 52 574 64 582
rect 82 574 94 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 0 564 4 572
rect 12 564 24 572
rect 42 564 54 572
rect 72 564 84 572
rect 102 564 114 574
rect 132 564 144 574
rect 162 564 174 574
rect 192 566 286 584
rect 314 566 408 584
rect 426 582 438 592
rect 456 582 468 592
rect 486 582 498 592
rect 516 584 528 592
rect 546 584 558 592
rect 576 584 588 592
rect 596 584 600 592
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 506 574 518 582
rect 536 574 548 582
rect 566 574 578 582
rect 586 574 600 582
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 0 554 14 562
rect 22 554 34 562
rect 52 554 64 562
rect 82 554 94 562
rect 112 554 124 562
rect 142 554 154 562
rect 172 554 184 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 192 554 408 566
rect 426 564 438 574
rect 456 564 468 574
rect 486 564 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 516 564 528 572
rect 546 564 558 572
rect 576 564 588 572
rect 596 564 600 572
rect 0 544 4 552
rect 12 544 24 552
rect 42 544 54 552
rect 72 544 84 552
rect 102 544 114 552
rect 132 544 144 552
rect 162 544 174 552
rect 192 546 286 554
rect 314 546 408 554
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 416 554 428 562
rect 446 554 458 562
rect 476 554 488 562
rect 506 554 518 562
rect 536 554 548 562
rect 566 554 578 562
rect 586 554 600 562
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 0 534 14 542
rect 22 534 34 542
rect 52 534 64 542
rect 82 534 94 542
rect 112 534 124 542
rect 142 534 154 542
rect 172 534 184 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 192 534 408 546
rect 426 544 438 552
rect 456 544 468 552
rect 486 544 498 552
rect 516 544 528 552
rect 546 544 558 552
rect 576 544 588 552
rect 596 544 600 552
rect 0 524 4 532
rect 12 524 24 532
rect 42 524 54 532
rect 72 524 84 532
rect 102 524 114 532
rect 132 524 144 532
rect 162 524 174 532
rect 192 526 286 534
rect 314 526 408 534
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 416 534 428 542
rect 446 534 458 542
rect 476 534 488 542
rect 506 534 518 542
rect 536 534 548 542
rect 566 534 578 542
rect 586 534 600 542
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 192 524 408 526
rect 426 524 438 532
rect 456 524 468 532
rect 486 524 498 532
rect 516 524 528 532
rect 546 524 558 532
rect 576 524 588 532
rect 596 524 600 532
rect 0 516 600 524
rect 0 512 24 516
rect 0 4 4 512
rect 12 508 24 512
rect 32 508 44 516
rect 52 508 64 516
rect 72 508 84 516
rect 92 508 104 516
rect 112 508 124 516
rect 132 508 144 516
rect 152 508 164 516
rect 172 508 184 516
rect 192 514 408 516
rect 192 508 286 514
rect 12 506 286 508
rect 314 508 408 514
rect 416 508 428 516
rect 436 508 448 516
rect 456 508 468 516
rect 476 508 488 516
rect 496 508 508 516
rect 516 508 528 516
rect 536 508 548 516
rect 556 508 568 516
rect 576 512 600 516
rect 576 508 588 512
rect 314 506 588 508
rect 12 504 588 506
rect 12 16 16 504
rect 584 16 588 504
rect 12 12 588 16
rect 192 4 408 12
rect 596 4 600 512
rect 0 0 600 4
<< psubstratepcontact >>
rect 2 1320 260 1338
rect 340 1320 598 1338
rect 2 840 20 1320
rect 44 836 52 844
rect 74 836 82 844
rect 104 836 112 844
rect 134 836 142 844
rect 164 836 172 844
rect 194 836 202 844
rect 224 836 232 844
rect 244 836 262 844
rect 274 836 282 844
rect 296 836 304 844
rect 318 836 326 844
rect 338 836 356 844
rect 368 836 376 844
rect 398 836 406 844
rect 428 836 436 844
rect 458 836 466 844
rect 488 836 496 844
rect 518 836 526 844
rect 548 836 556 844
rect 580 840 598 1320
rect 4 828 12 836
rect 24 828 42 836
rect 54 828 72 836
rect 84 828 102 836
rect 114 828 132 836
rect 144 828 162 836
rect 174 828 192 836
rect 204 828 222 836
rect 234 828 242 836
rect 264 828 272 836
rect 286 828 294 836
rect 306 828 314 836
rect 328 828 336 836
rect 358 828 366 836
rect 378 828 396 836
rect 408 828 426 836
rect 438 828 456 836
rect 468 828 486 836
rect 498 828 516 836
rect 528 828 546 836
rect 558 828 576 836
rect 588 828 596 836
rect 34 826 42 828
rect 64 826 72 828
rect 94 826 102 828
rect 124 826 132 828
rect 154 826 162 828
rect 184 826 192 828
rect 214 826 222 828
rect 378 826 386 828
rect 408 826 416 828
rect 438 826 446 828
rect 468 826 476 828
rect 498 826 506 828
rect 528 826 536 828
rect 558 826 566 828
rect 14 818 22 826
rect 34 818 52 826
rect 64 818 82 826
rect 94 818 112 826
rect 124 818 142 826
rect 154 818 172 826
rect 184 818 202 826
rect 214 818 232 826
rect 244 818 262 826
rect 274 818 282 826
rect 296 818 304 826
rect 318 818 326 826
rect 338 818 356 826
rect 368 818 386 826
rect 398 818 416 826
rect 428 818 446 826
rect 458 818 476 826
rect 488 818 506 826
rect 518 818 536 826
rect 548 818 566 826
rect 578 818 586 826
rect 34 816 42 818
rect 64 816 72 818
rect 94 816 102 818
rect 124 816 132 818
rect 154 816 162 818
rect 184 816 192 818
rect 214 816 222 818
rect 378 816 386 818
rect 408 816 416 818
rect 438 816 446 818
rect 468 816 476 818
rect 498 816 506 818
rect 528 816 536 818
rect 558 816 566 818
rect 4 808 12 816
rect 24 808 42 816
rect 54 808 72 816
rect 84 808 102 816
rect 114 808 132 816
rect 144 808 162 816
rect 174 808 192 816
rect 204 808 222 816
rect 234 808 242 816
rect 264 808 272 816
rect 286 808 294 816
rect 306 808 314 816
rect 328 808 336 816
rect 358 808 366 816
rect 378 808 396 816
rect 408 808 426 816
rect 438 808 456 816
rect 468 808 486 816
rect 498 808 516 816
rect 528 808 546 816
rect 558 808 576 816
rect 588 808 596 816
rect 34 806 42 808
rect 64 806 72 808
rect 94 806 102 808
rect 124 806 132 808
rect 154 806 162 808
rect 184 806 192 808
rect 214 806 222 808
rect 378 806 386 808
rect 408 806 416 808
rect 438 806 446 808
rect 468 806 476 808
rect 498 806 506 808
rect 528 806 536 808
rect 558 806 566 808
rect 14 798 22 806
rect 34 798 52 806
rect 64 798 82 806
rect 94 798 112 806
rect 124 798 142 806
rect 154 798 172 806
rect 184 798 202 806
rect 214 798 232 806
rect 244 798 262 806
rect 274 798 282 806
rect 296 798 304 806
rect 318 798 326 806
rect 338 798 356 806
rect 368 798 386 806
rect 398 798 416 806
rect 428 798 446 806
rect 458 798 476 806
rect 488 798 506 806
rect 518 798 536 806
rect 548 798 566 806
rect 578 798 586 806
rect 34 796 42 798
rect 64 796 72 798
rect 94 796 102 798
rect 124 796 132 798
rect 154 796 162 798
rect 184 796 192 798
rect 214 796 222 798
rect 378 796 386 798
rect 408 796 416 798
rect 438 796 446 798
rect 468 796 476 798
rect 498 796 506 798
rect 528 796 536 798
rect 558 796 566 798
rect 4 788 12 796
rect 24 788 42 796
rect 54 788 72 796
rect 84 788 102 796
rect 114 788 132 796
rect 144 788 162 796
rect 174 788 192 796
rect 204 788 222 796
rect 234 788 242 796
rect 264 788 272 796
rect 286 788 294 796
rect 306 788 314 796
rect 328 788 336 796
rect 358 788 366 796
rect 378 788 396 796
rect 408 788 426 796
rect 438 788 456 796
rect 468 788 486 796
rect 498 788 516 796
rect 528 788 546 796
rect 558 788 576 796
rect 588 788 596 796
rect 34 786 42 788
rect 64 786 72 788
rect 94 786 102 788
rect 124 786 132 788
rect 154 786 162 788
rect 184 786 192 788
rect 214 786 222 788
rect 378 786 386 788
rect 408 786 416 788
rect 438 786 446 788
rect 468 786 476 788
rect 498 786 506 788
rect 528 786 536 788
rect 558 786 566 788
rect 14 778 22 786
rect 34 778 52 786
rect 64 778 82 786
rect 34 776 42 778
rect 64 776 72 778
rect 94 776 112 786
rect 124 776 142 786
rect 154 776 172 786
rect 184 776 202 786
rect 214 776 232 786
rect 244 776 262 786
rect 274 776 282 786
rect 4 768 12 776
rect 24 768 42 776
rect 54 768 72 776
rect 84 768 292 776
rect 34 766 42 768
rect 64 766 72 768
rect 14 758 22 766
rect 34 758 52 766
rect 64 758 82 766
rect 94 758 112 768
rect 124 758 142 768
rect 154 758 172 768
rect 184 758 202 768
rect 214 758 232 768
rect 244 758 262 768
rect 274 758 282 768
rect 296 758 304 786
rect 318 776 326 786
rect 338 776 356 786
rect 368 776 386 786
rect 398 776 416 786
rect 428 776 446 786
rect 458 776 476 786
rect 488 776 506 786
rect 518 778 536 786
rect 548 778 566 786
rect 578 778 586 786
rect 528 776 536 778
rect 558 776 566 778
rect 308 768 516 776
rect 528 768 546 776
rect 558 768 576 776
rect 588 768 596 776
rect 318 758 326 768
rect 338 758 356 768
rect 368 758 386 768
rect 398 758 416 768
rect 428 758 446 768
rect 458 758 476 768
rect 488 758 506 768
rect 528 766 536 768
rect 558 766 566 768
rect 518 758 536 766
rect 548 758 566 766
rect 578 758 586 766
rect 34 756 42 758
rect 64 756 72 758
rect 94 756 102 758
rect 124 756 132 758
rect 154 756 162 758
rect 184 756 192 758
rect 214 756 222 758
rect 378 756 386 758
rect 408 756 416 758
rect 438 756 446 758
rect 468 756 476 758
rect 498 756 506 758
rect 528 756 536 758
rect 558 756 566 758
rect 4 748 12 756
rect 24 748 42 756
rect 54 748 72 756
rect 84 748 102 756
rect 114 748 132 756
rect 144 748 162 756
rect 174 748 192 756
rect 204 748 222 756
rect 234 748 242 756
rect 264 748 272 756
rect 286 748 294 756
rect 306 748 314 756
rect 328 748 336 756
rect 358 748 366 756
rect 378 748 396 756
rect 408 748 426 756
rect 438 748 456 756
rect 468 748 486 756
rect 498 748 516 756
rect 528 748 546 756
rect 558 748 576 756
rect 588 748 596 756
rect 34 746 42 748
rect 64 746 72 748
rect 94 746 102 748
rect 124 746 132 748
rect 154 746 162 748
rect 184 746 192 748
rect 214 746 222 748
rect 378 746 386 748
rect 408 746 416 748
rect 438 746 446 748
rect 468 746 476 748
rect 498 746 506 748
rect 528 746 536 748
rect 558 746 566 748
rect 14 738 22 746
rect 34 738 52 746
rect 64 738 82 746
rect 94 738 112 746
rect 124 738 142 746
rect 154 738 172 746
rect 184 738 202 746
rect 214 738 232 746
rect 244 738 262 746
rect 274 738 282 746
rect 296 738 304 746
rect 318 738 326 746
rect 338 738 356 746
rect 368 738 386 746
rect 398 738 416 746
rect 428 738 446 746
rect 458 738 476 746
rect 488 738 506 746
rect 518 738 536 746
rect 548 738 566 746
rect 578 738 586 746
rect 4 728 12 736
rect 24 728 32 736
rect 214 726 222 738
rect 234 728 242 736
rect 286 728 294 736
rect 306 728 314 736
rect 358 728 366 736
rect 378 726 386 738
rect 568 728 576 736
rect 588 728 596 736
rect 14 718 22 726
rect 34 718 52 726
rect 64 718 82 726
rect 94 718 112 726
rect 124 718 142 726
rect 154 718 172 726
rect 184 718 202 726
rect 214 718 232 726
rect 244 718 262 726
rect 296 718 304 726
rect 338 718 356 726
rect 368 718 386 726
rect 398 718 416 726
rect 428 718 446 726
rect 458 718 476 726
rect 488 718 506 726
rect 518 718 536 726
rect 548 718 566 726
rect 578 718 586 726
rect 34 716 42 718
rect 64 716 72 718
rect 94 716 102 718
rect 124 716 132 718
rect 154 716 162 718
rect 184 716 192 718
rect 214 716 222 718
rect 378 716 386 718
rect 408 716 416 718
rect 438 716 446 718
rect 468 716 476 718
rect 498 716 506 718
rect 528 716 536 718
rect 558 716 566 718
rect 4 708 12 716
rect 24 708 42 716
rect 54 708 72 716
rect 84 708 102 716
rect 114 708 132 716
rect 144 708 162 716
rect 174 708 192 716
rect 204 708 222 716
rect 234 708 242 716
rect 264 708 272 716
rect 286 708 294 716
rect 306 708 314 716
rect 328 708 336 716
rect 358 708 366 716
rect 378 708 396 716
rect 408 708 426 716
rect 438 708 456 716
rect 468 708 486 716
rect 498 708 516 716
rect 528 708 546 716
rect 558 708 576 716
rect 588 708 596 716
rect 34 706 42 708
rect 64 706 72 708
rect 94 706 102 708
rect 124 706 132 708
rect 154 706 162 708
rect 184 706 192 708
rect 214 706 222 708
rect 378 706 386 708
rect 408 706 416 708
rect 438 706 446 708
rect 468 706 476 708
rect 498 706 506 708
rect 528 706 536 708
rect 558 706 566 708
rect 14 698 22 706
rect 34 698 52 706
rect 64 698 82 706
rect 94 698 112 706
rect 124 698 142 706
rect 154 698 172 706
rect 184 698 202 706
rect 214 698 232 706
rect 244 698 262 706
rect 274 698 282 706
rect 296 698 304 706
rect 318 698 326 706
rect 338 698 356 706
rect 368 698 386 706
rect 398 698 416 706
rect 428 698 446 706
rect 458 698 476 706
rect 488 698 506 706
rect 518 698 536 706
rect 548 698 566 706
rect 578 698 586 706
rect 34 696 42 698
rect 64 696 72 698
rect 94 696 102 698
rect 124 696 132 698
rect 154 696 162 698
rect 184 696 192 698
rect 214 696 222 698
rect 4 688 12 696
rect 24 688 42 696
rect 54 688 72 696
rect 84 688 102 696
rect 114 688 132 696
rect 144 688 162 696
rect 174 688 192 696
rect 204 688 222 696
rect 234 688 242 696
rect 286 689 294 697
rect 306 689 314 697
rect 378 696 386 698
rect 408 696 416 698
rect 438 696 446 698
rect 468 696 476 698
rect 498 696 506 698
rect 528 696 536 698
rect 558 696 566 698
rect 358 688 366 696
rect 378 688 396 696
rect 408 688 426 696
rect 438 688 456 696
rect 468 688 486 696
rect 498 688 516 696
rect 528 688 546 696
rect 558 688 576 696
rect 588 688 596 696
rect 30 461 568 489
rect 40 451 48 461
rect 60 451 78 461
rect 90 451 108 461
rect 120 451 138 461
rect 150 451 168 461
rect 180 451 198 461
rect 210 451 228 461
rect 240 451 258 461
rect 270 451 288 461
rect 300 451 318 461
rect 330 451 348 461
rect 360 451 378 461
rect 390 451 408 461
rect 420 451 438 461
rect 450 451 468 461
rect 480 451 498 461
rect 510 451 528 461
rect 540 451 558 461
rect 60 449 68 451
rect 90 449 98 451
rect 120 449 128 451
rect 150 449 158 451
rect 180 449 188 451
rect 210 449 218 451
rect 240 449 248 451
rect 270 449 278 451
rect 300 449 308 451
rect 330 449 338 451
rect 360 449 368 451
rect 390 449 398 451
rect 420 449 428 451
rect 450 449 458 451
rect 480 449 488 451
rect 510 449 518 451
rect 540 449 548 451
rect 30 441 38 449
rect 50 441 68 449
rect 80 441 98 449
rect 110 441 128 449
rect 140 441 158 449
rect 170 441 188 449
rect 200 441 218 449
rect 230 441 248 449
rect 260 441 278 449
rect 290 441 308 449
rect 320 441 338 449
rect 350 441 368 449
rect 380 441 398 449
rect 410 441 428 449
rect 440 441 458 449
rect 470 441 488 449
rect 500 441 518 449
rect 530 441 548 449
rect 560 441 568 449
rect 60 439 68 441
rect 90 439 98 441
rect 120 439 128 441
rect 150 439 158 441
rect 180 439 188 441
rect 210 439 218 441
rect 240 439 248 441
rect 270 439 278 441
rect 300 439 308 441
rect 330 439 338 441
rect 360 439 368 441
rect 390 439 398 441
rect 420 439 428 441
rect 450 439 458 441
rect 480 439 488 441
rect 510 439 518 441
rect 540 439 548 441
rect 40 431 48 439
rect 60 431 78 439
rect 90 431 108 439
rect 120 431 138 439
rect 150 431 168 439
rect 180 431 198 439
rect 210 431 228 439
rect 240 431 258 439
rect 270 431 288 439
rect 300 431 318 439
rect 330 431 348 439
rect 360 431 378 439
rect 390 431 408 439
rect 420 431 438 439
rect 450 431 468 439
rect 480 431 498 439
rect 510 431 528 439
rect 540 431 558 439
rect 60 429 68 431
rect 90 429 98 431
rect 120 429 128 431
rect 150 429 158 431
rect 180 429 188 431
rect 210 429 218 431
rect 240 429 248 431
rect 270 429 278 431
rect 300 429 308 431
rect 330 429 338 431
rect 360 429 368 431
rect 390 429 398 431
rect 420 429 428 431
rect 450 429 458 431
rect 480 429 488 431
rect 510 429 518 431
rect 540 429 548 431
rect 30 421 38 429
rect 50 421 68 429
rect 80 421 98 429
rect 110 421 128 429
rect 140 421 158 429
rect 170 421 188 429
rect 200 421 218 429
rect 230 421 248 429
rect 260 421 278 429
rect 290 421 308 429
rect 320 421 338 429
rect 350 421 368 429
rect 380 421 398 429
rect 410 421 428 429
rect 440 421 458 429
rect 470 421 488 429
rect 500 421 518 429
rect 530 421 548 429
rect 560 421 568 429
rect 60 419 68 421
rect 90 419 98 421
rect 120 419 128 421
rect 150 419 158 421
rect 180 419 188 421
rect 210 419 218 421
rect 240 419 248 421
rect 270 419 278 421
rect 300 419 308 421
rect 330 419 338 421
rect 360 419 368 421
rect 390 419 398 421
rect 420 419 428 421
rect 450 419 458 421
rect 480 419 488 421
rect 510 419 518 421
rect 540 419 548 421
rect 40 411 48 419
rect 60 411 78 419
rect 90 411 108 419
rect 120 411 138 419
rect 150 411 168 419
rect 180 411 198 419
rect 210 411 228 419
rect 240 411 258 419
rect 270 411 288 419
rect 300 411 318 419
rect 330 411 348 419
rect 360 411 378 419
rect 390 411 408 419
rect 420 411 438 419
rect 450 411 468 419
rect 480 411 498 419
rect 510 411 528 419
rect 540 411 558 419
rect 60 409 68 411
rect 90 409 98 411
rect 120 409 128 411
rect 150 409 158 411
rect 180 409 188 411
rect 210 409 218 411
rect 240 409 248 411
rect 270 409 278 411
rect 300 409 308 411
rect 330 409 338 411
rect 360 409 368 411
rect 390 409 398 411
rect 420 409 428 411
rect 450 409 458 411
rect 480 409 488 411
rect 510 409 518 411
rect 540 409 548 411
rect 30 401 38 409
rect 50 401 68 409
rect 80 401 98 409
rect 110 401 128 409
rect 140 401 158 409
rect 170 401 188 409
rect 200 401 218 409
rect 230 401 248 409
rect 260 401 278 409
rect 290 401 308 409
rect 320 401 338 409
rect 350 401 368 409
rect 380 401 398 409
rect 410 401 428 409
rect 440 401 458 409
rect 470 401 488 409
rect 500 401 518 409
rect 530 401 548 409
rect 560 401 568 409
rect 60 399 68 401
rect 90 399 98 401
rect 120 399 128 401
rect 150 399 158 401
rect 180 399 188 401
rect 210 399 218 401
rect 240 399 248 401
rect 270 399 278 401
rect 300 399 308 401
rect 330 399 338 401
rect 360 399 368 401
rect 390 399 398 401
rect 420 399 428 401
rect 450 399 458 401
rect 480 399 488 401
rect 510 399 518 401
rect 540 399 548 401
rect 40 371 48 399
rect 60 371 78 399
rect 90 391 108 399
rect 120 391 138 399
rect 150 391 168 399
rect 180 391 198 399
rect 210 391 228 399
rect 240 391 258 399
rect 270 391 288 399
rect 300 391 318 399
rect 330 391 348 399
rect 360 391 378 399
rect 390 391 408 399
rect 420 391 438 399
rect 450 391 468 399
rect 480 391 498 399
rect 510 391 528 399
rect 540 391 558 399
rect 90 379 98 391
rect 510 379 518 391
rect 540 389 548 391
rect 530 381 548 389
rect 560 381 568 389
rect 540 379 548 381
rect 90 371 108 379
rect 120 371 138 379
rect 150 371 168 379
rect 180 371 198 379
rect 210 371 228 379
rect 240 371 258 379
rect 270 371 288 379
rect 300 371 318 379
rect 330 371 348 379
rect 360 371 378 379
rect 390 371 408 379
rect 420 371 438 379
rect 450 371 468 379
rect 480 371 498 379
rect 510 371 528 379
rect 540 371 558 379
rect 60 369 68 371
rect 90 369 98 371
rect 120 369 128 371
rect 150 369 158 371
rect 180 369 188 371
rect 210 369 218 371
rect 240 369 248 371
rect 270 369 278 371
rect 300 369 308 371
rect 330 369 338 371
rect 360 369 368 371
rect 390 369 398 371
rect 420 369 428 371
rect 450 369 458 371
rect 480 369 488 371
rect 510 369 518 371
rect 540 369 548 371
rect 30 361 38 369
rect 50 361 68 369
rect 80 361 98 369
rect 110 361 128 369
rect 140 361 158 369
rect 170 361 188 369
rect 200 361 218 369
rect 230 361 248 369
rect 260 361 278 369
rect 290 361 308 369
rect 320 361 338 369
rect 350 361 368 369
rect 380 361 398 369
rect 410 361 428 369
rect 440 361 458 369
rect 470 361 488 369
rect 500 361 518 369
rect 530 361 548 369
rect 560 361 568 369
rect 60 359 68 361
rect 90 359 98 361
rect 120 359 128 361
rect 150 359 158 361
rect 180 359 188 361
rect 210 359 218 361
rect 240 359 248 361
rect 270 359 278 361
rect 300 359 308 361
rect 330 359 338 361
rect 360 359 368 361
rect 390 359 398 361
rect 420 359 428 361
rect 450 359 458 361
rect 480 359 488 361
rect 510 359 518 361
rect 540 359 548 361
rect 40 351 48 359
rect 60 351 78 359
rect 90 351 108 359
rect 120 351 138 359
rect 150 351 168 359
rect 180 351 198 359
rect 210 351 228 359
rect 240 351 258 359
rect 270 351 288 359
rect 300 351 318 359
rect 330 351 348 359
rect 360 351 378 359
rect 390 351 408 359
rect 420 351 438 359
rect 450 351 468 359
rect 480 351 498 359
rect 510 351 528 359
rect 540 351 558 359
rect 60 349 68 351
rect 90 349 98 351
rect 120 349 128 351
rect 150 349 158 351
rect 180 349 188 351
rect 210 349 218 351
rect 240 349 248 351
rect 270 349 278 351
rect 300 349 308 351
rect 330 349 338 351
rect 360 349 368 351
rect 390 349 398 351
rect 420 349 428 351
rect 450 349 458 351
rect 480 349 488 351
rect 510 349 518 351
rect 540 349 548 351
rect 30 341 38 349
rect 50 341 68 349
rect 80 341 98 349
rect 110 341 128 349
rect 140 341 158 349
rect 170 341 188 349
rect 200 341 218 349
rect 230 341 248 349
rect 260 341 278 349
rect 290 341 308 349
rect 320 341 338 349
rect 350 341 368 349
rect 380 341 398 349
rect 410 341 428 349
rect 440 341 458 349
rect 470 341 488 349
rect 500 341 518 349
rect 530 341 548 349
rect 560 341 568 349
rect 60 339 68 341
rect 90 339 98 341
rect 120 339 128 341
rect 150 339 158 341
rect 180 339 188 341
rect 210 339 218 341
rect 240 339 248 341
rect 270 339 278 341
rect 300 339 308 341
rect 330 339 338 341
rect 360 339 368 341
rect 390 339 398 341
rect 420 339 428 341
rect 450 339 458 341
rect 480 339 488 341
rect 510 339 518 341
rect 540 339 548 341
rect 40 331 48 339
rect 60 331 78 339
rect 90 331 108 339
rect 120 331 138 339
rect 150 331 168 339
rect 180 331 198 339
rect 210 331 228 339
rect 240 331 258 339
rect 270 331 288 339
rect 300 331 318 339
rect 330 331 348 339
rect 360 331 378 339
rect 390 331 408 339
rect 420 331 438 339
rect 450 331 468 339
rect 480 331 498 339
rect 510 331 528 339
rect 540 331 558 339
rect 60 329 68 331
rect 90 329 98 331
rect 120 329 128 331
rect 150 329 158 331
rect 180 329 188 331
rect 210 329 218 331
rect 240 329 248 331
rect 270 329 278 331
rect 300 329 308 331
rect 330 329 338 331
rect 360 329 368 331
rect 390 329 398 331
rect 420 329 428 331
rect 450 329 458 331
rect 480 329 488 331
rect 510 329 518 331
rect 540 329 548 331
rect 30 321 38 329
rect 50 321 68 329
rect 80 321 98 329
rect 110 321 128 329
rect 140 321 158 329
rect 170 321 188 329
rect 200 321 218 329
rect 230 321 248 329
rect 260 321 278 329
rect 290 321 308 329
rect 320 321 338 329
rect 350 321 368 329
rect 380 321 398 329
rect 410 321 428 329
rect 440 321 458 329
rect 470 321 488 329
rect 500 321 518 329
rect 530 321 548 329
rect 560 321 568 329
rect 60 319 68 321
rect 90 319 98 321
rect 120 319 128 321
rect 150 319 158 321
rect 180 319 188 321
rect 210 319 218 321
rect 240 319 248 321
rect 270 319 278 321
rect 300 319 308 321
rect 330 319 338 321
rect 360 319 368 321
rect 390 319 398 321
rect 420 319 428 321
rect 450 319 458 321
rect 480 319 488 321
rect 510 319 518 321
rect 540 319 548 321
rect 40 311 48 319
rect 60 311 78 319
rect 90 311 108 319
rect 120 311 138 319
rect 150 311 168 319
rect 180 311 198 319
rect 210 311 228 319
rect 240 311 258 319
rect 270 311 288 319
rect 300 311 318 319
rect 330 311 348 319
rect 360 311 378 319
rect 390 311 408 319
rect 420 311 438 319
rect 450 311 468 319
rect 480 311 498 319
rect 510 311 528 319
rect 540 311 558 319
rect 60 309 68 311
rect 510 309 518 311
rect 540 309 548 311
rect 30 301 38 309
rect 50 301 68 309
rect 80 301 88 309
rect 500 301 518 309
rect 530 301 548 309
rect 560 301 568 309
rect 60 299 68 301
rect 510 299 518 301
rect 540 299 548 301
rect 40 291 48 299
rect 60 291 78 299
rect 90 291 108 299
rect 120 291 138 299
rect 150 291 168 299
rect 180 291 198 299
rect 210 291 228 299
rect 240 291 258 299
rect 270 291 288 299
rect 300 291 318 299
rect 330 291 348 299
rect 360 291 378 299
rect 390 291 408 299
rect 420 291 438 299
rect 450 291 468 299
rect 480 291 498 299
rect 510 291 528 299
rect 540 291 558 299
rect 60 289 68 291
rect 90 289 98 291
rect 120 289 128 291
rect 150 289 158 291
rect 180 289 188 291
rect 210 289 218 291
rect 240 289 248 291
rect 270 289 278 291
rect 300 289 308 291
rect 330 289 338 291
rect 360 289 368 291
rect 390 289 398 291
rect 420 289 428 291
rect 450 289 458 291
rect 480 289 488 291
rect 510 289 518 291
rect 540 289 548 291
rect 30 281 38 289
rect 50 281 68 289
rect 80 281 98 289
rect 110 281 128 289
rect 140 281 158 289
rect 170 281 188 289
rect 200 281 218 289
rect 230 281 248 289
rect 260 281 278 289
rect 290 281 308 289
rect 320 281 338 289
rect 350 281 368 289
rect 380 281 398 289
rect 410 281 428 289
rect 440 281 458 289
rect 470 281 488 289
rect 500 281 518 289
rect 530 281 548 289
rect 560 281 568 289
rect 60 279 68 281
rect 90 279 98 281
rect 120 279 128 281
rect 150 279 158 281
rect 180 279 188 281
rect 210 279 218 281
rect 240 279 248 281
rect 270 279 278 281
rect 300 279 308 281
rect 330 279 338 281
rect 360 279 368 281
rect 390 279 398 281
rect 420 279 428 281
rect 450 279 458 281
rect 480 279 488 281
rect 510 279 518 281
rect 540 279 548 281
rect 40 271 48 279
rect 60 271 78 279
rect 90 271 108 279
rect 120 271 138 279
rect 150 271 168 279
rect 180 271 198 279
rect 210 271 228 279
rect 240 271 258 279
rect 270 271 288 279
rect 300 271 318 279
rect 330 271 348 279
rect 360 271 378 279
rect 390 271 408 279
rect 420 271 438 279
rect 450 271 468 279
rect 480 271 498 279
rect 510 271 528 279
rect 540 271 558 279
rect 60 269 68 271
rect 90 269 98 271
rect 120 269 128 271
rect 150 269 158 271
rect 180 269 188 271
rect 210 269 218 271
rect 240 269 248 271
rect 270 269 278 271
rect 300 269 308 271
rect 330 269 338 271
rect 360 269 368 271
rect 390 269 398 271
rect 420 269 428 271
rect 450 269 458 271
rect 480 269 488 271
rect 510 269 518 271
rect 540 269 548 271
rect 30 261 38 269
rect 50 261 68 269
rect 80 261 98 269
rect 110 261 128 269
rect 140 261 158 269
rect 170 261 188 269
rect 200 261 218 269
rect 230 261 248 269
rect 260 261 278 269
rect 290 261 308 269
rect 320 261 338 269
rect 350 261 368 269
rect 380 261 398 269
rect 410 261 428 269
rect 440 261 458 269
rect 470 261 488 269
rect 500 261 518 269
rect 530 261 548 269
rect 560 261 568 269
rect 60 259 68 261
rect 90 259 98 261
rect 120 259 128 261
rect 150 259 158 261
rect 180 259 188 261
rect 210 259 218 261
rect 240 259 248 261
rect 270 259 278 261
rect 300 259 308 261
rect 330 259 338 261
rect 360 259 368 261
rect 390 259 398 261
rect 420 259 428 261
rect 450 259 458 261
rect 480 259 488 261
rect 510 259 518 261
rect 540 259 548 261
rect 40 251 48 259
rect 60 251 78 259
rect 90 251 108 259
rect 120 251 138 259
rect 150 251 168 259
rect 180 251 198 259
rect 210 251 228 259
rect 240 251 258 259
rect 270 251 288 259
rect 300 251 318 259
rect 330 251 348 259
rect 360 251 378 259
rect 390 251 408 259
rect 420 251 438 259
rect 450 251 468 259
rect 480 251 498 259
rect 510 251 528 259
rect 540 251 558 259
rect 60 249 68 251
rect 90 249 98 251
rect 120 249 128 251
rect 150 249 158 251
rect 180 249 188 251
rect 210 249 218 251
rect 240 249 248 251
rect 270 249 278 251
rect 300 249 308 251
rect 330 249 338 251
rect 360 249 368 251
rect 390 249 398 251
rect 420 249 428 251
rect 450 249 458 251
rect 480 249 488 251
rect 510 249 518 251
rect 540 249 548 251
rect 30 241 38 249
rect 50 241 68 249
rect 40 231 48 239
rect 60 229 68 241
rect 30 221 38 229
rect 50 221 68 229
rect 80 241 98 249
rect 110 241 128 249
rect 140 241 158 249
rect 170 241 188 249
rect 200 241 218 249
rect 230 241 248 249
rect 260 241 278 249
rect 290 241 308 249
rect 320 241 338 249
rect 350 241 368 249
rect 380 241 398 249
rect 410 241 428 249
rect 440 241 458 249
rect 470 241 488 249
rect 500 241 518 249
rect 530 241 548 249
rect 560 241 568 249
rect 80 229 88 241
rect 500 229 508 241
rect 540 239 548 241
rect 520 231 528 239
rect 540 231 558 239
rect 540 229 548 231
rect 80 221 98 229
rect 110 221 128 229
rect 140 221 158 229
rect 170 221 188 229
rect 200 221 218 229
rect 230 221 248 229
rect 260 221 278 229
rect 290 221 308 229
rect 320 221 338 229
rect 350 221 368 229
rect 380 221 398 229
rect 410 221 428 229
rect 440 221 458 229
rect 470 221 488 229
rect 500 221 518 229
rect 530 221 548 229
rect 560 221 568 229
rect 60 219 68 221
rect 90 219 98 221
rect 120 219 128 221
rect 150 219 158 221
rect 180 219 188 221
rect 210 219 218 221
rect 240 219 248 221
rect 270 219 278 221
rect 300 219 308 221
rect 330 219 338 221
rect 360 219 368 221
rect 390 219 398 221
rect 420 219 428 221
rect 450 219 458 221
rect 480 219 488 221
rect 510 219 518 221
rect 540 219 548 221
rect 40 211 48 219
rect 60 211 78 219
rect 90 211 108 219
rect 120 211 138 219
rect 150 211 168 219
rect 180 211 198 219
rect 210 211 228 219
rect 240 211 258 219
rect 270 211 288 219
rect 300 211 318 219
rect 330 211 348 219
rect 360 211 378 219
rect 390 211 408 219
rect 420 211 438 219
rect 450 211 468 219
rect 480 211 498 219
rect 510 211 528 219
rect 540 211 558 219
rect 60 209 68 211
rect 90 209 98 211
rect 120 209 128 211
rect 150 209 158 211
rect 180 209 188 211
rect 210 209 218 211
rect 240 209 248 211
rect 270 209 278 211
rect 300 209 308 211
rect 330 209 338 211
rect 360 209 368 211
rect 390 209 398 211
rect 420 209 428 211
rect 450 209 458 211
rect 480 209 488 211
rect 510 209 518 211
rect 540 209 548 211
rect 30 201 38 209
rect 50 201 68 209
rect 80 201 98 209
rect 110 201 128 209
rect 140 201 158 209
rect 170 201 188 209
rect 200 201 218 209
rect 230 201 248 209
rect 260 201 278 209
rect 290 201 308 209
rect 320 201 338 209
rect 350 201 368 209
rect 380 201 398 209
rect 410 201 428 209
rect 440 201 458 209
rect 470 201 488 209
rect 500 201 518 209
rect 530 201 548 209
rect 560 201 568 209
rect 60 199 68 201
rect 90 199 98 201
rect 120 199 128 201
rect 150 199 158 201
rect 180 199 188 201
rect 210 199 218 201
rect 240 199 248 201
rect 270 199 278 201
rect 300 199 308 201
rect 330 199 338 201
rect 360 199 368 201
rect 390 199 398 201
rect 420 199 428 201
rect 450 199 458 201
rect 480 199 488 201
rect 510 199 518 201
rect 540 199 548 201
rect 40 191 48 199
rect 60 191 78 199
rect 90 191 108 199
rect 120 191 138 199
rect 150 191 168 199
rect 180 191 198 199
rect 210 191 228 199
rect 240 191 258 199
rect 270 191 288 199
rect 300 191 318 199
rect 330 191 348 199
rect 360 191 378 199
rect 390 191 408 199
rect 420 191 438 199
rect 450 191 468 199
rect 480 191 498 199
rect 510 191 528 199
rect 540 191 558 199
rect 60 189 68 191
rect 90 189 98 191
rect 120 189 128 191
rect 150 189 158 191
rect 180 189 188 191
rect 210 189 218 191
rect 240 189 248 191
rect 270 189 278 191
rect 300 189 308 191
rect 330 189 338 191
rect 360 189 368 191
rect 390 189 398 191
rect 420 189 428 191
rect 450 189 458 191
rect 480 189 488 191
rect 510 189 518 191
rect 540 189 548 191
rect 30 181 38 189
rect 50 181 68 189
rect 80 181 98 189
rect 110 181 128 189
rect 140 181 158 189
rect 170 181 188 189
rect 200 181 218 189
rect 230 181 248 189
rect 260 181 278 189
rect 290 181 308 189
rect 320 181 338 189
rect 350 181 368 189
rect 380 181 398 189
rect 410 181 428 189
rect 440 181 458 189
rect 470 181 488 189
rect 500 181 518 189
rect 530 181 548 189
rect 560 181 568 189
rect 60 179 68 181
rect 90 179 98 181
rect 120 179 128 181
rect 150 179 158 181
rect 180 179 188 181
rect 210 179 218 181
rect 240 179 248 181
rect 270 179 278 181
rect 300 179 308 181
rect 330 179 338 181
rect 360 179 368 181
rect 390 179 398 181
rect 420 179 428 181
rect 450 179 458 181
rect 480 179 488 181
rect 510 179 518 181
rect 540 179 548 181
rect 40 171 48 179
rect 60 171 78 179
rect 90 171 108 179
rect 120 171 138 179
rect 150 171 168 179
rect 180 171 198 179
rect 210 171 228 179
rect 240 171 258 179
rect 270 171 288 179
rect 300 171 318 179
rect 330 171 348 179
rect 360 171 378 179
rect 390 171 408 179
rect 420 171 438 179
rect 450 171 468 179
rect 480 171 498 179
rect 510 171 528 179
rect 540 171 558 179
rect 60 169 68 171
rect 90 169 98 171
rect 120 169 128 171
rect 150 169 158 171
rect 180 169 188 171
rect 210 169 218 171
rect 240 169 248 171
rect 270 169 278 171
rect 300 169 308 171
rect 330 169 338 171
rect 360 169 368 171
rect 390 169 398 171
rect 420 169 428 171
rect 450 169 458 171
rect 480 169 488 171
rect 510 169 518 171
rect 540 169 548 171
rect 30 161 38 169
rect 50 161 68 169
rect 80 161 98 169
rect 110 161 128 169
rect 140 161 158 169
rect 170 161 188 169
rect 200 161 218 169
rect 230 161 248 169
rect 260 161 278 169
rect 290 161 308 169
rect 320 161 338 169
rect 350 161 368 169
rect 380 161 398 169
rect 410 161 428 169
rect 440 161 458 169
rect 470 161 488 169
rect 500 161 518 169
rect 530 161 548 169
rect 560 161 568 169
rect 60 159 68 161
rect 40 151 48 159
rect 60 151 78 159
rect 60 149 68 151
rect 90 149 98 161
rect 500 149 508 161
rect 540 159 548 161
rect 520 151 528 159
rect 540 151 558 159
rect 540 149 548 151
rect 30 141 38 149
rect 50 141 68 149
rect 80 141 98 149
rect 110 141 128 149
rect 140 141 158 149
rect 170 141 188 149
rect 200 141 218 149
rect 230 141 248 149
rect 260 141 278 149
rect 290 141 308 149
rect 320 141 338 149
rect 350 141 368 149
rect 380 141 398 149
rect 410 141 428 149
rect 440 141 458 149
rect 470 141 488 149
rect 500 141 518 149
rect 530 141 548 149
rect 560 141 568 149
rect 60 139 68 141
rect 90 139 98 141
rect 120 139 128 141
rect 150 139 158 141
rect 180 139 188 141
rect 210 139 218 141
rect 240 139 248 141
rect 270 139 278 141
rect 300 139 308 141
rect 330 139 338 141
rect 360 139 368 141
rect 390 139 398 141
rect 420 139 428 141
rect 450 139 458 141
rect 480 139 488 141
rect 510 139 518 141
rect 540 139 548 141
rect 40 131 48 139
rect 60 131 78 139
rect 90 131 108 139
rect 120 131 138 139
rect 150 131 168 139
rect 180 131 198 139
rect 210 131 228 139
rect 240 131 258 139
rect 270 131 288 139
rect 300 131 318 139
rect 330 131 348 139
rect 360 131 378 139
rect 390 131 408 139
rect 420 131 438 139
rect 450 131 468 139
rect 480 131 498 139
rect 510 131 528 139
rect 540 131 558 139
rect 60 129 68 131
rect 90 129 98 131
rect 120 129 128 131
rect 150 129 158 131
rect 180 129 188 131
rect 210 129 218 131
rect 240 129 248 131
rect 270 129 278 131
rect 300 129 308 131
rect 330 129 338 131
rect 360 129 368 131
rect 390 129 398 131
rect 420 129 428 131
rect 450 129 458 131
rect 480 129 488 131
rect 510 129 518 131
rect 540 129 548 131
rect 30 121 38 129
rect 50 121 68 129
rect 80 121 98 129
rect 110 121 128 129
rect 140 121 158 129
rect 170 121 188 129
rect 200 121 218 129
rect 230 121 248 129
rect 260 121 278 129
rect 290 121 308 129
rect 320 121 338 129
rect 350 121 368 129
rect 380 121 398 129
rect 410 121 428 129
rect 440 121 458 129
rect 470 121 488 129
rect 500 121 518 129
rect 530 121 548 129
rect 560 121 568 129
rect 60 119 68 121
rect 90 119 98 121
rect 120 119 128 121
rect 150 119 158 121
rect 180 119 188 121
rect 210 119 218 121
rect 240 119 248 121
rect 270 119 278 121
rect 300 119 308 121
rect 330 119 338 121
rect 360 119 368 121
rect 390 119 398 121
rect 420 119 428 121
rect 450 119 458 121
rect 480 119 488 121
rect 510 119 518 121
rect 540 119 548 121
rect 40 111 48 119
rect 60 111 78 119
rect 90 111 108 119
rect 120 111 138 119
rect 150 111 168 119
rect 180 111 198 119
rect 210 111 228 119
rect 240 111 258 119
rect 270 111 288 119
rect 300 111 318 119
rect 330 111 348 119
rect 360 111 378 119
rect 390 111 408 119
rect 420 111 438 119
rect 450 111 468 119
rect 480 111 498 119
rect 510 111 528 119
rect 540 111 558 119
rect 60 109 68 111
rect 90 109 98 111
rect 120 109 128 111
rect 150 109 158 111
rect 180 109 188 111
rect 210 109 218 111
rect 240 109 248 111
rect 270 109 278 111
rect 300 109 308 111
rect 330 109 338 111
rect 360 109 368 111
rect 390 109 398 111
rect 420 109 428 111
rect 450 109 458 111
rect 480 109 488 111
rect 510 109 518 111
rect 540 109 548 111
rect 30 101 38 109
rect 50 101 68 109
rect 80 101 98 109
rect 110 101 128 109
rect 140 101 158 109
rect 170 101 188 109
rect 200 101 218 109
rect 230 101 248 109
rect 260 101 278 109
rect 290 101 308 109
rect 320 101 338 109
rect 350 101 368 109
rect 380 101 398 109
rect 410 101 428 109
rect 440 101 458 109
rect 470 101 488 109
rect 500 101 518 109
rect 530 101 548 109
rect 560 101 568 109
rect 60 99 68 101
rect 90 99 98 101
rect 120 99 128 101
rect 150 99 158 101
rect 180 99 188 101
rect 210 99 218 101
rect 240 99 248 101
rect 270 99 278 101
rect 300 99 308 101
rect 330 99 338 101
rect 360 99 368 101
rect 390 99 398 101
rect 420 99 428 101
rect 450 99 458 101
rect 480 99 488 101
rect 510 99 518 101
rect 540 99 548 101
rect 40 91 48 99
rect 60 91 78 99
rect 90 91 108 99
rect 120 91 138 99
rect 150 91 168 99
rect 180 91 198 99
rect 210 91 228 99
rect 240 91 258 99
rect 270 91 288 99
rect 300 91 318 99
rect 330 91 348 99
rect 360 91 378 99
rect 390 91 408 99
rect 420 91 438 99
rect 450 91 468 99
rect 480 91 498 99
rect 510 91 528 99
rect 540 91 558 99
rect 60 89 68 91
rect 90 89 98 91
rect 120 89 128 91
rect 150 89 158 91
rect 180 89 188 91
rect 210 89 218 91
rect 240 89 248 91
rect 270 89 278 91
rect 300 89 308 91
rect 330 89 338 91
rect 360 89 368 91
rect 390 89 398 91
rect 420 89 428 91
rect 450 89 458 91
rect 480 89 488 91
rect 510 89 518 91
rect 540 89 548 91
rect 30 81 38 89
rect 50 81 68 89
rect 80 81 98 89
rect 110 81 128 89
rect 140 81 158 89
rect 170 81 188 89
rect 200 81 218 89
rect 230 81 248 89
rect 260 81 278 89
rect 290 81 308 89
rect 320 81 338 89
rect 350 81 368 89
rect 380 81 398 89
rect 410 81 428 89
rect 440 81 458 89
rect 470 81 488 89
rect 500 81 518 89
rect 530 81 548 89
rect 560 81 568 89
rect 60 79 68 81
rect 90 79 98 81
rect 120 79 128 81
rect 150 79 158 81
rect 180 79 188 81
rect 210 79 218 81
rect 240 79 248 81
rect 270 79 278 81
rect 300 79 308 81
rect 330 79 338 81
rect 360 79 368 81
rect 390 79 398 81
rect 420 79 428 81
rect 450 79 458 81
rect 480 79 488 81
rect 510 79 518 81
rect 540 79 548 81
rect 40 71 48 79
rect 60 71 78 79
rect 90 71 108 79
rect 120 71 138 79
rect 150 71 168 79
rect 180 71 198 79
rect 210 71 228 79
rect 240 71 258 79
rect 270 71 288 79
rect 300 71 318 79
rect 330 71 348 79
rect 360 71 378 79
rect 390 71 408 79
rect 420 71 438 79
rect 450 71 468 79
rect 480 71 498 79
rect 510 71 528 79
rect 540 71 558 79
rect 60 69 68 71
rect 90 69 98 71
rect 120 69 128 71
rect 150 69 158 71
rect 180 69 188 71
rect 210 69 218 71
rect 240 69 248 71
rect 270 69 278 71
rect 300 69 308 71
rect 330 69 338 71
rect 360 69 368 71
rect 390 69 398 71
rect 420 69 428 71
rect 450 69 458 71
rect 480 69 488 71
rect 510 69 518 71
rect 540 69 548 71
rect 30 61 38 69
rect 50 61 68 69
rect 80 61 98 69
rect 110 61 128 69
rect 140 61 158 69
rect 170 61 188 69
rect 200 61 218 69
rect 230 61 248 69
rect 260 61 278 69
rect 290 61 308 69
rect 320 61 338 69
rect 350 61 368 69
rect 380 61 398 69
rect 410 61 428 69
rect 440 61 458 69
rect 470 61 488 69
rect 500 61 518 69
rect 530 61 548 69
rect 560 61 568 69
rect 60 59 68 61
rect 90 59 98 61
rect 120 59 128 61
rect 150 59 158 61
rect 180 59 188 61
rect 210 59 218 61
rect 240 59 248 61
rect 270 59 278 61
rect 300 59 308 61
rect 330 59 338 61
rect 360 59 368 61
rect 390 59 398 61
rect 420 59 428 61
rect 450 59 458 61
rect 480 59 488 61
rect 510 59 518 61
rect 540 59 548 61
rect 40 51 48 59
rect 60 51 78 59
rect 90 51 108 59
rect 120 51 138 59
rect 150 51 168 59
rect 180 51 198 59
rect 210 51 228 59
rect 240 51 258 59
rect 270 51 288 59
rect 300 51 318 59
rect 330 51 348 59
rect 360 51 378 59
rect 390 51 408 59
rect 420 51 438 59
rect 450 51 468 59
rect 480 51 498 59
rect 510 51 528 59
rect 540 51 558 59
rect 60 49 68 51
rect 90 49 98 51
rect 120 49 128 51
rect 150 49 158 51
rect 180 49 188 51
rect 210 49 218 51
rect 240 49 248 51
rect 270 49 278 51
rect 300 49 308 51
rect 330 49 338 51
rect 360 49 368 51
rect 390 49 398 51
rect 420 49 428 51
rect 450 49 458 51
rect 480 49 488 51
rect 510 49 518 51
rect 540 49 548 51
rect 30 41 38 49
rect 50 41 68 49
rect 80 41 98 49
rect 110 41 128 49
rect 140 41 158 49
rect 170 41 188 49
rect 200 41 218 49
rect 230 41 248 49
rect 260 41 278 49
rect 290 41 308 49
rect 320 41 338 49
rect 350 41 368 49
rect 380 41 398 49
rect 410 41 428 49
rect 440 41 458 49
rect 470 41 488 49
rect 500 41 518 49
rect 530 41 548 49
rect 560 41 568 49
rect 60 39 68 41
rect 90 39 98 41
rect 120 39 128 41
rect 150 39 158 41
rect 180 39 188 41
rect 210 39 218 41
rect 240 39 248 41
rect 270 39 278 41
rect 300 39 308 41
rect 330 39 338 41
rect 360 39 368 41
rect 390 39 398 41
rect 420 39 428 41
rect 450 39 458 41
rect 480 39 488 41
rect 510 39 518 41
rect 540 39 548 41
rect 40 31 48 39
rect 60 31 78 39
rect 90 31 108 39
rect 120 31 138 39
rect 150 31 168 39
rect 180 31 198 39
rect 210 31 228 39
rect 240 31 258 39
rect 270 31 288 39
rect 300 31 318 39
rect 330 31 348 39
rect 360 31 378 39
rect 390 31 408 39
rect 420 31 438 39
rect 450 31 468 39
rect 480 31 498 39
rect 510 31 528 39
rect 540 31 558 39
<< nsubstratencontact >>
rect 51 1290 59 1298
rect 72 1294 80 1298
rect 520 1294 528 1298
rect 72 1290 90 1294
rect 41 1280 49 1288
rect 62 1281 70 1289
rect 82 1286 90 1290
rect 102 1286 110 1294
rect 122 1286 130 1294
rect 142 1286 150 1294
rect 162 1286 170 1294
rect 182 1286 190 1294
rect 202 1286 210 1294
rect 222 1286 230 1294
rect 370 1286 378 1294
rect 390 1286 398 1294
rect 410 1286 418 1294
rect 430 1286 438 1294
rect 450 1286 458 1294
rect 470 1286 478 1294
rect 490 1286 498 1294
rect 510 1290 528 1294
rect 541 1290 549 1298
rect 510 1286 518 1290
rect 51 1270 59 1278
rect 41 1260 49 1268
rect 92 1276 100 1284
rect 112 1276 120 1284
rect 132 1276 140 1284
rect 152 1276 160 1284
rect 172 1276 180 1284
rect 192 1276 200 1284
rect 212 1276 220 1284
rect 232 1276 240 1284
rect 51 1250 59 1258
rect 41 1240 49 1248
rect 51 1230 59 1238
rect 41 1220 49 1228
rect 51 1210 59 1218
rect 41 1200 49 1208
rect 51 1190 59 1198
rect 41 1180 49 1188
rect 51 1170 59 1178
rect 41 1160 49 1168
rect 51 1150 59 1158
rect 41 1140 49 1148
rect 51 1130 59 1138
rect 41 1120 49 1128
rect 51 1110 59 1118
rect 41 1100 49 1108
rect 51 1090 59 1098
rect 41 1080 49 1088
rect 51 1070 59 1078
rect 41 1060 49 1068
rect 51 1050 59 1058
rect 41 1040 49 1048
rect 51 1030 59 1038
rect 41 1020 49 1028
rect 51 1010 59 1018
rect 41 1000 49 1008
rect 51 990 59 998
rect 41 980 49 988
rect 51 970 59 978
rect 41 960 49 968
rect 51 950 59 958
rect 41 940 49 948
rect 51 930 59 938
rect 41 920 49 928
rect 51 910 59 918
rect 41 900 49 908
rect 360 1276 368 1284
rect 380 1276 388 1284
rect 400 1276 408 1284
rect 420 1276 428 1284
rect 440 1276 448 1284
rect 460 1276 468 1284
rect 480 1276 488 1284
rect 500 1276 508 1284
rect 530 1281 538 1289
rect 551 1280 559 1288
rect 541 1270 549 1278
rect 551 1260 559 1268
rect 286 1222 314 1230
rect 286 1202 314 1210
rect 286 1182 314 1190
rect 286 1094 314 1102
rect 286 1074 314 1082
rect 286 1054 314 1062
rect 286 964 314 972
rect 286 944 314 952
rect 286 924 314 932
rect 51 890 59 898
rect 41 880 49 888
rect 541 1250 549 1258
rect 551 1240 559 1248
rect 541 1230 549 1238
rect 551 1220 559 1228
rect 541 1210 549 1218
rect 551 1200 559 1208
rect 541 1190 549 1198
rect 551 1180 559 1188
rect 541 1170 549 1178
rect 551 1160 559 1168
rect 541 1150 549 1158
rect 551 1140 559 1148
rect 541 1130 549 1138
rect 551 1120 559 1128
rect 541 1110 549 1118
rect 551 1100 559 1108
rect 541 1090 549 1098
rect 551 1080 559 1088
rect 541 1070 549 1078
rect 551 1060 559 1068
rect 541 1050 549 1058
rect 551 1040 559 1048
rect 541 1030 549 1038
rect 551 1020 559 1028
rect 541 1010 549 1018
rect 551 1000 559 1008
rect 541 990 549 998
rect 551 980 559 988
rect 541 970 549 978
rect 551 960 559 968
rect 541 950 549 958
rect 551 940 559 948
rect 541 930 549 938
rect 551 920 559 928
rect 541 910 549 918
rect 551 900 559 908
rect 541 890 549 898
rect 62 873 240 883
rect 42 865 240 873
rect 360 873 538 883
rect 551 880 559 888
rect 360 865 558 873
rect 4 644 12 652
rect 24 644 42 652
rect 54 644 72 652
rect 84 644 102 652
rect 114 644 132 652
rect 144 644 162 652
rect 174 644 192 652
rect 34 642 42 644
rect 64 642 72 644
rect 94 642 102 644
rect 124 642 132 644
rect 154 642 162 644
rect 14 634 22 642
rect 34 634 52 642
rect 64 634 82 642
rect 94 634 112 642
rect 124 634 142 642
rect 154 634 172 642
rect 34 632 42 634
rect 64 632 72 634
rect 94 632 102 634
rect 124 632 132 634
rect 154 632 162 634
rect 184 632 192 644
rect 408 644 426 652
rect 438 644 456 652
rect 468 644 486 652
rect 498 644 516 652
rect 528 644 546 652
rect 558 644 576 652
rect 588 644 596 652
rect 286 634 314 642
rect 4 624 12 632
rect 24 624 42 632
rect 54 624 72 632
rect 84 624 102 632
rect 114 624 132 632
rect 144 624 162 632
rect 174 624 192 632
rect 34 622 42 624
rect 64 622 72 624
rect 94 622 102 624
rect 124 622 132 624
rect 154 622 162 624
rect 14 614 22 622
rect 34 614 52 622
rect 64 614 82 622
rect 94 614 112 622
rect 124 614 142 622
rect 154 614 172 622
rect 184 614 192 624
rect 408 632 416 644
rect 438 642 446 644
rect 468 642 476 644
rect 498 642 506 644
rect 528 642 536 644
rect 558 642 566 644
rect 428 634 446 642
rect 458 634 476 642
rect 488 634 506 642
rect 518 634 536 642
rect 548 634 566 642
rect 578 634 586 642
rect 438 632 446 634
rect 468 632 476 634
rect 498 632 506 634
rect 528 632 536 634
rect 558 632 566 634
rect 408 624 426 632
rect 438 624 456 632
rect 468 624 486 632
rect 498 624 516 632
rect 528 624 546 632
rect 558 624 576 632
rect 588 624 596 632
rect 286 614 314 622
rect 408 614 416 624
rect 438 622 446 624
rect 468 622 476 624
rect 498 622 506 624
rect 528 622 536 624
rect 558 622 566 624
rect 428 614 446 622
rect 458 614 476 622
rect 488 614 506 622
rect 518 614 536 622
rect 548 614 566 622
rect 578 614 586 622
rect 4 604 12 612
rect 24 604 32 612
rect 568 604 576 612
rect 588 604 596 612
rect 14 594 22 602
rect 34 594 52 602
rect 64 594 82 602
rect 94 594 112 602
rect 124 594 142 602
rect 154 594 172 602
rect 34 592 42 594
rect 64 592 72 594
rect 94 592 102 594
rect 124 592 132 594
rect 154 592 162 594
rect 184 592 192 602
rect 286 594 314 602
rect 4 584 12 592
rect 24 584 42 592
rect 54 584 72 592
rect 84 584 102 592
rect 34 582 42 584
rect 64 582 72 584
rect 94 582 102 584
rect 114 582 132 592
rect 144 582 162 592
rect 174 582 192 592
rect 408 592 416 602
rect 428 594 446 602
rect 458 594 476 602
rect 488 594 506 602
rect 518 594 536 602
rect 548 594 566 602
rect 578 594 586 602
rect 438 592 446 594
rect 468 592 476 594
rect 498 592 506 594
rect 528 592 536 594
rect 558 592 566 594
rect 14 574 22 582
rect 34 574 52 582
rect 64 574 82 582
rect 94 574 192 582
rect 34 572 42 574
rect 64 572 72 574
rect 94 572 102 574
rect 4 564 12 572
rect 24 564 42 572
rect 54 564 72 572
rect 84 564 102 572
rect 114 564 132 574
rect 144 564 162 574
rect 174 564 192 574
rect 286 566 314 584
rect 408 582 426 592
rect 438 582 456 592
rect 468 582 486 592
rect 498 584 516 592
rect 528 584 546 592
rect 558 584 576 592
rect 588 584 596 592
rect 498 582 506 584
rect 528 582 536 584
rect 558 582 566 584
rect 408 574 506 582
rect 518 574 536 582
rect 548 574 566 582
rect 578 574 586 582
rect 34 562 42 564
rect 64 562 72 564
rect 94 562 102 564
rect 124 562 132 564
rect 154 562 162 564
rect 14 554 22 562
rect 34 554 52 562
rect 64 554 82 562
rect 94 554 112 562
rect 124 554 142 562
rect 154 554 172 562
rect 34 552 42 554
rect 64 552 72 554
rect 94 552 102 554
rect 124 552 132 554
rect 154 552 162 554
rect 184 552 192 564
rect 408 564 426 574
rect 438 564 456 574
rect 468 564 486 574
rect 498 572 506 574
rect 528 572 536 574
rect 558 572 566 574
rect 498 564 516 572
rect 528 564 546 572
rect 558 564 576 572
rect 588 564 596 572
rect 4 544 12 552
rect 24 544 42 552
rect 54 544 72 552
rect 84 544 102 552
rect 114 544 132 552
rect 144 544 162 552
rect 174 544 192 552
rect 286 546 314 554
rect 408 552 416 564
rect 438 562 446 564
rect 468 562 476 564
rect 498 562 506 564
rect 528 562 536 564
rect 558 562 566 564
rect 428 554 446 562
rect 458 554 476 562
rect 488 554 506 562
rect 518 554 536 562
rect 548 554 566 562
rect 578 554 586 562
rect 438 552 446 554
rect 468 552 476 554
rect 498 552 506 554
rect 528 552 536 554
rect 558 552 566 554
rect 34 542 42 544
rect 64 542 72 544
rect 94 542 102 544
rect 124 542 132 544
rect 154 542 162 544
rect 14 534 22 542
rect 34 534 52 542
rect 64 534 82 542
rect 94 534 112 542
rect 124 534 142 542
rect 154 534 172 542
rect 34 532 42 534
rect 64 532 72 534
rect 94 532 102 534
rect 124 532 132 534
rect 154 532 162 534
rect 184 532 192 544
rect 408 544 426 552
rect 438 544 456 552
rect 468 544 486 552
rect 498 544 516 552
rect 528 544 546 552
rect 558 544 576 552
rect 588 544 596 552
rect 4 524 12 532
rect 24 524 42 532
rect 54 524 72 532
rect 84 524 102 532
rect 114 524 132 532
rect 144 524 162 532
rect 174 524 192 532
rect 286 526 314 534
rect 408 532 416 544
rect 438 542 446 544
rect 468 542 476 544
rect 498 542 506 544
rect 528 542 536 544
rect 558 542 566 544
rect 428 534 446 542
rect 458 534 476 542
rect 488 534 506 542
rect 518 534 536 542
rect 548 534 566 542
rect 578 534 586 542
rect 438 532 446 534
rect 468 532 476 534
rect 498 532 506 534
rect 528 532 536 534
rect 558 532 566 534
rect 408 524 426 532
rect 438 524 456 532
rect 468 524 486 532
rect 498 524 516 532
rect 528 524 546 532
rect 558 524 576 532
rect 588 524 596 532
rect 4 12 12 512
rect 24 508 32 516
rect 44 508 52 516
rect 64 508 72 516
rect 84 508 92 516
rect 104 508 112 516
rect 124 508 132 516
rect 144 508 152 516
rect 164 508 172 516
rect 184 508 192 516
rect 286 506 314 514
rect 408 508 416 516
rect 428 508 436 516
rect 448 508 456 516
rect 468 508 476 516
rect 488 508 496 516
rect 508 508 516 516
rect 528 508 536 516
rect 548 508 556 516
rect 568 508 576 516
rect 588 12 596 512
rect 4 4 192 12
rect 408 4 596 12
<< polysilicon >>
rect 62 1252 76 1258
rect 276 1252 280 1258
rect 62 914 64 1252
rect 72 1170 74 1252
rect 320 1252 324 1258
rect 524 1252 538 1258
rect 72 1164 76 1170
rect 276 1164 280 1170
rect 72 1130 74 1164
rect 72 1124 76 1130
rect 276 1124 280 1130
rect 72 1042 74 1124
rect 526 1170 528 1252
rect 320 1164 324 1170
rect 524 1164 528 1170
rect 526 1130 528 1164
rect 320 1124 324 1130
rect 524 1124 528 1130
rect 72 1036 76 1042
rect 276 1036 280 1042
rect 72 1000 74 1036
rect 72 994 76 1000
rect 276 994 280 1000
rect 72 914 74 994
rect 62 912 74 914
rect 526 1042 528 1124
rect 320 1036 324 1042
rect 524 1036 528 1042
rect 526 1000 528 1036
rect 320 994 324 1000
rect 524 994 528 1000
rect 62 906 76 912
rect 276 906 280 912
rect 526 914 528 994
rect 536 914 538 1252
rect 526 912 538 914
rect 320 906 324 912
rect 524 906 538 912
<< polycontact >>
rect 64 914 72 1252
rect 528 914 536 1252
<< metal1 >>
rect 124 1460 476 1480
rect 144 1440 456 1460
rect 164 1420 436 1440
rect 184 1400 416 1420
rect 204 1340 396 1400
rect 0 1338 600 1340
rect 0 840 2 1338
rect 260 1320 340 1338
rect 20 1318 580 1320
rect 20 846 22 1318
rect 204 1306 396 1318
rect 72 1298 240 1300
rect 41 1290 42 1298
rect 50 1290 51 1298
rect 59 1290 62 1298
rect 70 1290 72 1298
rect 80 1294 240 1298
rect 41 1289 72 1290
rect 41 1288 62 1289
rect 49 1287 62 1288
rect 49 1280 50 1287
rect 41 1279 50 1280
rect 58 1281 62 1287
rect 70 1282 72 1289
rect 80 1286 82 1290
rect 90 1286 92 1294
rect 100 1286 102 1294
rect 110 1286 112 1294
rect 120 1286 122 1294
rect 130 1286 132 1294
rect 140 1286 142 1294
rect 150 1286 152 1294
rect 160 1286 162 1294
rect 170 1286 172 1294
rect 180 1286 182 1294
rect 190 1286 192 1294
rect 200 1286 202 1294
rect 210 1286 212 1294
rect 220 1286 222 1294
rect 230 1286 232 1294
rect 80 1284 240 1286
rect 70 1281 82 1282
rect 58 1279 82 1281
rect 41 1278 82 1279
rect 41 1270 42 1278
rect 50 1270 51 1278
rect 59 1276 82 1278
rect 90 1276 92 1284
rect 100 1276 102 1284
rect 110 1276 112 1284
rect 120 1276 122 1284
rect 130 1276 132 1284
rect 140 1276 142 1284
rect 150 1276 152 1284
rect 160 1276 162 1284
rect 170 1276 172 1284
rect 180 1276 182 1284
rect 190 1276 192 1284
rect 200 1276 202 1284
rect 210 1276 212 1284
rect 220 1276 222 1284
rect 230 1276 232 1284
rect 59 1274 240 1276
rect 59 1270 82 1274
rect 41 1268 82 1270
rect 49 1267 82 1268
rect 49 1260 50 1267
rect 41 1259 50 1260
rect 58 1266 82 1267
rect 58 1259 240 1266
rect 41 1258 240 1259
rect 41 1250 42 1258
rect 50 1250 51 1258
rect 59 1252 240 1258
rect 59 1250 64 1252
rect 41 1248 64 1250
rect 49 1247 64 1248
rect 49 1240 50 1247
rect 41 1239 50 1240
rect 58 1239 64 1247
rect 41 1238 64 1239
rect 41 1230 42 1238
rect 50 1230 51 1238
rect 59 1230 64 1238
rect 41 1228 64 1230
rect 49 1227 64 1228
rect 49 1220 50 1227
rect 41 1219 50 1220
rect 58 1219 64 1227
rect 41 1218 64 1219
rect 41 1210 42 1218
rect 50 1210 51 1218
rect 59 1210 64 1218
rect 41 1208 64 1210
rect 49 1207 64 1208
rect 49 1200 50 1207
rect 41 1199 50 1200
rect 58 1199 64 1207
rect 41 1198 64 1199
rect 41 1190 42 1198
rect 50 1190 51 1198
rect 59 1190 64 1198
rect 41 1188 64 1190
rect 49 1187 64 1188
rect 49 1180 50 1187
rect 41 1179 50 1180
rect 58 1179 64 1187
rect 41 1178 64 1179
rect 41 1170 42 1178
rect 50 1170 51 1178
rect 59 1170 64 1178
rect 41 1168 64 1170
rect 49 1167 64 1168
rect 49 1160 50 1167
rect 41 1159 50 1160
rect 58 1159 64 1167
rect 41 1158 64 1159
rect 41 1150 42 1158
rect 50 1150 51 1158
rect 59 1150 64 1158
rect 41 1148 64 1150
rect 49 1147 64 1148
rect 49 1140 50 1147
rect 41 1139 50 1140
rect 58 1139 64 1147
rect 41 1138 64 1139
rect 41 1130 42 1138
rect 50 1130 51 1138
rect 59 1130 64 1138
rect 41 1128 64 1130
rect 49 1127 64 1128
rect 49 1120 50 1127
rect 41 1119 50 1120
rect 58 1119 64 1127
rect 41 1118 64 1119
rect 41 1110 42 1118
rect 50 1110 51 1118
rect 59 1110 64 1118
rect 41 1108 64 1110
rect 49 1107 64 1108
rect 49 1100 50 1107
rect 41 1099 50 1100
rect 58 1099 64 1107
rect 41 1098 64 1099
rect 41 1090 42 1098
rect 50 1090 51 1098
rect 59 1090 64 1098
rect 41 1088 64 1090
rect 49 1087 64 1088
rect 49 1080 50 1087
rect 41 1079 50 1080
rect 58 1079 64 1087
rect 41 1078 64 1079
rect 41 1070 42 1078
rect 50 1070 51 1078
rect 59 1070 64 1078
rect 41 1068 64 1070
rect 49 1067 64 1068
rect 49 1060 50 1067
rect 41 1059 50 1060
rect 58 1059 64 1067
rect 41 1058 64 1059
rect 41 1050 42 1058
rect 50 1050 51 1058
rect 59 1050 64 1058
rect 41 1048 64 1050
rect 49 1047 64 1048
rect 49 1040 50 1047
rect 41 1039 50 1040
rect 58 1039 64 1047
rect 41 1038 64 1039
rect 41 1030 42 1038
rect 50 1030 51 1038
rect 59 1030 64 1038
rect 41 1028 64 1030
rect 49 1027 64 1028
rect 49 1020 50 1027
rect 41 1019 50 1020
rect 58 1019 64 1027
rect 41 1018 64 1019
rect 41 1010 42 1018
rect 50 1010 51 1018
rect 59 1010 64 1018
rect 41 1008 64 1010
rect 49 1007 64 1008
rect 49 1000 50 1007
rect 41 999 50 1000
rect 58 999 64 1007
rect 41 998 64 999
rect 41 990 42 998
rect 50 990 51 998
rect 59 990 64 998
rect 41 988 64 990
rect 49 987 64 988
rect 49 980 50 987
rect 41 979 50 980
rect 58 979 64 987
rect 41 978 64 979
rect 41 970 42 978
rect 50 970 51 978
rect 59 970 64 978
rect 41 968 64 970
rect 49 967 64 968
rect 49 960 50 967
rect 41 959 50 960
rect 58 959 64 967
rect 41 958 64 959
rect 41 950 42 958
rect 50 950 51 958
rect 59 950 64 958
rect 41 948 64 950
rect 49 947 64 948
rect 49 940 50 947
rect 41 939 50 940
rect 58 939 64 947
rect 41 938 64 939
rect 41 930 42 938
rect 50 930 51 938
rect 59 930 64 938
rect 41 928 64 930
rect 49 927 64 928
rect 49 920 50 927
rect 41 919 50 920
rect 58 919 64 927
rect 41 918 64 919
rect 41 910 42 918
rect 50 910 51 918
rect 59 914 64 918
rect 72 1250 240 1252
rect 72 1172 78 1250
rect 236 1242 240 1250
rect 96 1180 102 1242
rect 246 1236 354 1306
rect 360 1298 528 1300
rect 360 1294 520 1298
rect 368 1286 370 1294
rect 378 1286 380 1294
rect 388 1286 390 1294
rect 398 1286 400 1294
rect 408 1286 410 1294
rect 418 1286 420 1294
rect 428 1286 430 1294
rect 438 1286 440 1294
rect 448 1286 450 1294
rect 458 1286 460 1294
rect 468 1286 470 1294
rect 478 1286 480 1294
rect 488 1286 490 1294
rect 498 1286 500 1294
rect 508 1286 510 1294
rect 528 1290 530 1298
rect 538 1290 541 1298
rect 549 1290 550 1298
rect 558 1290 559 1298
rect 518 1286 520 1290
rect 360 1284 520 1286
rect 528 1289 559 1290
rect 368 1276 370 1284
rect 378 1276 380 1284
rect 388 1276 390 1284
rect 398 1276 400 1284
rect 408 1276 410 1284
rect 418 1276 420 1284
rect 428 1276 430 1284
rect 438 1276 440 1284
rect 448 1276 450 1284
rect 458 1276 460 1284
rect 468 1276 470 1284
rect 478 1276 480 1284
rect 488 1276 490 1284
rect 498 1276 500 1284
rect 508 1276 510 1284
rect 528 1282 530 1289
rect 518 1281 530 1282
rect 538 1288 559 1289
rect 538 1287 551 1288
rect 538 1281 542 1287
rect 518 1279 542 1281
rect 550 1280 551 1287
rect 550 1279 559 1280
rect 518 1278 559 1279
rect 518 1276 541 1278
rect 360 1274 541 1276
rect 518 1270 541 1274
rect 549 1270 550 1278
rect 558 1270 559 1278
rect 518 1268 559 1270
rect 518 1267 551 1268
rect 518 1266 542 1267
rect 360 1259 542 1266
rect 550 1260 551 1267
rect 550 1259 559 1260
rect 360 1258 559 1259
rect 360 1252 541 1258
rect 360 1250 528 1252
rect 360 1242 364 1250
rect 112 1220 280 1236
rect 240 1202 280 1220
rect 112 1186 280 1202
rect 236 1172 240 1180
rect 72 1156 240 1172
rect 72 1138 82 1156
rect 72 1122 240 1138
rect 72 1044 78 1122
rect 236 1114 240 1122
rect 246 1176 280 1186
rect 286 1220 314 1222
rect 286 1212 290 1220
rect 298 1212 302 1220
rect 310 1212 314 1220
rect 286 1210 314 1212
rect 286 1200 314 1202
rect 286 1192 290 1200
rect 298 1192 302 1200
rect 310 1192 314 1200
rect 286 1190 314 1192
rect 320 1220 488 1236
rect 320 1202 360 1220
rect 320 1186 488 1202
rect 320 1176 354 1186
rect 498 1180 504 1242
rect 96 1052 102 1114
rect 246 1108 354 1176
rect 360 1172 364 1180
rect 522 1172 528 1250
rect 360 1156 528 1172
rect 518 1138 528 1156
rect 360 1122 528 1138
rect 360 1114 364 1122
rect 112 1092 280 1108
rect 240 1074 280 1092
rect 112 1058 280 1074
rect 236 1044 240 1052
rect 72 1028 240 1044
rect 72 1020 82 1028
rect 72 1016 240 1020
rect 72 1008 82 1016
rect 72 992 240 1008
rect 72 914 78 992
rect 236 984 240 992
rect 246 1048 280 1058
rect 286 1092 314 1094
rect 286 1084 290 1092
rect 298 1084 302 1092
rect 310 1084 314 1092
rect 286 1082 314 1084
rect 286 1072 314 1074
rect 286 1064 290 1072
rect 298 1064 302 1072
rect 310 1064 314 1072
rect 286 1062 314 1064
rect 320 1092 488 1108
rect 320 1074 360 1092
rect 320 1058 488 1074
rect 320 1048 354 1058
rect 498 1052 504 1114
rect 96 922 102 984
rect 246 978 354 1048
rect 360 1044 364 1052
rect 522 1044 528 1122
rect 360 1028 528 1044
rect 518 1020 528 1028
rect 360 1016 528 1020
rect 518 1008 528 1016
rect 360 992 528 1008
rect 360 984 364 992
rect 112 962 280 978
rect 240 944 280 962
rect 112 928 280 944
rect 236 914 240 922
rect 59 910 240 914
rect 41 908 240 910
rect 49 907 240 908
rect 49 900 50 907
rect 41 899 50 900
rect 58 899 240 907
rect 41 898 240 899
rect 41 890 42 898
rect 50 890 51 898
rect 59 890 82 898
rect 41 888 240 890
rect 49 880 50 888
rect 58 883 240 888
rect 58 880 62 883
rect 41 873 62 880
rect 41 865 42 873
rect 246 918 280 928
rect 286 962 314 964
rect 286 954 290 962
rect 298 954 302 962
rect 310 954 314 962
rect 286 952 314 954
rect 286 942 314 944
rect 286 934 290 942
rect 298 934 302 942
rect 310 934 314 942
rect 286 932 314 934
rect 320 962 488 978
rect 320 944 360 962
rect 320 928 488 944
rect 320 918 354 928
rect 498 922 504 984
rect 246 859 354 918
rect 360 914 364 922
rect 522 914 528 992
rect 536 1250 541 1252
rect 549 1250 550 1258
rect 558 1250 559 1258
rect 536 1248 559 1250
rect 536 1247 551 1248
rect 536 1239 542 1247
rect 550 1240 551 1247
rect 550 1239 559 1240
rect 536 1238 559 1239
rect 536 1230 541 1238
rect 549 1230 550 1238
rect 558 1230 559 1238
rect 536 1228 559 1230
rect 536 1227 551 1228
rect 536 1219 542 1227
rect 550 1220 551 1227
rect 550 1219 559 1220
rect 536 1218 559 1219
rect 536 1210 541 1218
rect 549 1210 550 1218
rect 558 1210 559 1218
rect 536 1208 559 1210
rect 536 1207 551 1208
rect 536 1199 542 1207
rect 550 1200 551 1207
rect 550 1199 559 1200
rect 536 1198 559 1199
rect 536 1190 541 1198
rect 549 1190 550 1198
rect 558 1190 559 1198
rect 536 1188 559 1190
rect 536 1187 551 1188
rect 536 1179 542 1187
rect 550 1180 551 1187
rect 550 1179 559 1180
rect 536 1178 559 1179
rect 536 1170 541 1178
rect 549 1170 550 1178
rect 558 1170 559 1178
rect 536 1168 559 1170
rect 536 1167 551 1168
rect 536 1159 542 1167
rect 550 1160 551 1167
rect 550 1159 559 1160
rect 536 1158 559 1159
rect 536 1150 541 1158
rect 549 1150 550 1158
rect 558 1150 559 1158
rect 536 1148 559 1150
rect 536 1147 551 1148
rect 536 1139 542 1147
rect 550 1140 551 1147
rect 550 1139 559 1140
rect 536 1138 559 1139
rect 536 1130 541 1138
rect 549 1130 550 1138
rect 558 1130 559 1138
rect 536 1128 559 1130
rect 536 1127 551 1128
rect 536 1119 542 1127
rect 550 1120 551 1127
rect 550 1119 559 1120
rect 536 1118 559 1119
rect 536 1110 541 1118
rect 549 1110 550 1118
rect 558 1110 559 1118
rect 536 1108 559 1110
rect 536 1107 551 1108
rect 536 1099 542 1107
rect 550 1100 551 1107
rect 550 1099 559 1100
rect 536 1098 559 1099
rect 536 1090 541 1098
rect 549 1090 550 1098
rect 558 1090 559 1098
rect 536 1088 559 1090
rect 536 1087 551 1088
rect 536 1079 542 1087
rect 550 1080 551 1087
rect 550 1079 559 1080
rect 536 1078 559 1079
rect 536 1070 541 1078
rect 549 1070 550 1078
rect 558 1070 559 1078
rect 536 1068 559 1070
rect 536 1067 551 1068
rect 536 1059 542 1067
rect 550 1060 551 1067
rect 550 1059 559 1060
rect 536 1058 559 1059
rect 536 1050 541 1058
rect 549 1050 550 1058
rect 558 1050 559 1058
rect 536 1048 559 1050
rect 536 1047 551 1048
rect 536 1039 542 1047
rect 550 1040 551 1047
rect 550 1039 559 1040
rect 536 1038 559 1039
rect 536 1030 541 1038
rect 549 1030 550 1038
rect 558 1030 559 1038
rect 536 1028 559 1030
rect 536 1027 551 1028
rect 536 1019 542 1027
rect 550 1020 551 1027
rect 550 1019 559 1020
rect 536 1018 559 1019
rect 536 1010 541 1018
rect 549 1010 550 1018
rect 558 1010 559 1018
rect 536 1008 559 1010
rect 536 1007 551 1008
rect 536 999 542 1007
rect 550 1000 551 1007
rect 550 999 559 1000
rect 536 998 559 999
rect 536 990 541 998
rect 549 990 550 998
rect 558 990 559 998
rect 536 988 559 990
rect 536 987 551 988
rect 536 979 542 987
rect 550 980 551 987
rect 550 979 559 980
rect 536 978 559 979
rect 536 970 541 978
rect 549 970 550 978
rect 558 970 559 978
rect 536 968 559 970
rect 536 967 551 968
rect 536 959 542 967
rect 550 960 551 967
rect 550 959 559 960
rect 536 958 559 959
rect 536 950 541 958
rect 549 950 550 958
rect 558 950 559 958
rect 536 948 559 950
rect 536 947 551 948
rect 536 939 542 947
rect 550 940 551 947
rect 550 939 559 940
rect 536 938 559 939
rect 536 930 541 938
rect 549 930 550 938
rect 558 930 559 938
rect 536 928 559 930
rect 536 927 551 928
rect 536 919 542 927
rect 550 920 551 927
rect 550 919 559 920
rect 536 918 559 919
rect 536 914 541 918
rect 360 910 541 914
rect 549 910 550 918
rect 558 910 559 918
rect 360 908 559 910
rect 360 907 551 908
rect 360 899 542 907
rect 550 900 551 907
rect 550 899 559 900
rect 360 898 559 899
rect 518 890 541 898
rect 549 890 550 898
rect 558 890 559 898
rect 360 888 559 890
rect 360 883 542 888
rect 538 880 542 883
rect 550 880 551 888
rect 538 873 559 880
rect 558 865 559 873
rect 204 846 396 859
rect 578 846 580 1318
rect 20 844 580 846
rect 20 840 24 844
rect 0 836 24 840
rect 0 828 4 836
rect 12 828 14 836
rect 22 828 24 836
rect 42 828 44 844
rect 52 828 54 844
rect 72 828 74 844
rect 82 828 84 844
rect 102 828 104 844
rect 112 828 114 844
rect 132 828 134 844
rect 142 828 144 844
rect 162 828 164 844
rect 172 828 174 844
rect 192 828 194 844
rect 202 828 204 844
rect 222 828 224 844
rect 232 828 234 844
rect 242 828 244 844
rect 262 828 264 844
rect 272 828 274 844
rect 282 828 286 844
rect 294 828 296 844
rect 304 828 306 844
rect 314 828 318 844
rect 326 828 328 844
rect 336 828 338 844
rect 356 828 358 844
rect 366 828 368 844
rect 376 828 378 844
rect 396 828 398 844
rect 406 828 408 844
rect 426 828 428 844
rect 436 828 438 844
rect 456 828 458 844
rect 466 828 468 844
rect 486 828 488 844
rect 496 828 498 844
rect 516 828 518 844
rect 526 828 528 844
rect 546 828 548 844
rect 556 828 558 844
rect 576 840 580 844
rect 598 840 600 1338
rect 576 836 600 840
rect 576 828 578 836
rect 586 828 588 836
rect 596 828 600 836
rect 0 826 34 828
rect 42 826 64 828
rect 72 826 94 828
rect 102 826 124 828
rect 132 826 154 828
rect 162 826 184 828
rect 192 826 214 828
rect 222 826 378 828
rect 386 826 408 828
rect 416 826 438 828
rect 446 826 468 828
rect 476 826 498 828
rect 506 826 528 828
rect 536 826 558 828
rect 566 826 600 828
rect 0 818 4 826
rect 12 818 14 826
rect 22 818 24 826
rect 32 818 34 826
rect 52 818 54 826
rect 62 818 64 826
rect 82 818 84 826
rect 92 818 94 826
rect 112 818 114 826
rect 122 818 124 826
rect 142 818 144 826
rect 152 818 154 826
rect 172 818 174 826
rect 182 818 184 826
rect 202 818 204 826
rect 212 818 214 826
rect 232 818 234 826
rect 242 818 244 826
rect 262 818 264 826
rect 272 818 274 826
rect 282 818 286 826
rect 294 818 296 826
rect 304 818 306 826
rect 314 818 318 826
rect 326 818 328 826
rect 336 818 338 826
rect 356 818 358 826
rect 366 818 368 826
rect 386 818 388 826
rect 396 818 398 826
rect 416 818 418 826
rect 426 818 428 826
rect 446 818 448 826
rect 456 818 458 826
rect 476 818 478 826
rect 486 818 488 826
rect 506 818 508 826
rect 516 818 518 826
rect 536 818 538 826
rect 546 818 548 826
rect 566 818 568 826
rect 576 818 578 826
rect 586 818 588 826
rect 596 818 600 826
rect 0 816 34 818
rect 42 816 64 818
rect 72 816 94 818
rect 102 816 124 818
rect 132 816 154 818
rect 162 816 184 818
rect 192 816 214 818
rect 222 816 378 818
rect 386 816 408 818
rect 416 816 438 818
rect 446 816 468 818
rect 476 816 498 818
rect 506 816 528 818
rect 536 816 558 818
rect 566 816 600 818
rect 0 808 4 816
rect 12 808 14 816
rect 22 808 24 816
rect 42 808 44 816
rect 52 808 54 816
rect 72 808 74 816
rect 82 808 84 816
rect 102 808 104 816
rect 112 808 114 816
rect 132 808 134 816
rect 142 808 144 816
rect 162 808 164 816
rect 172 808 174 816
rect 192 808 194 816
rect 202 808 204 816
rect 222 808 224 816
rect 232 808 234 816
rect 242 808 244 816
rect 262 808 264 816
rect 272 808 276 816
rect 284 808 286 816
rect 294 808 296 816
rect 304 808 306 816
rect 314 808 316 816
rect 324 808 328 816
rect 336 808 338 816
rect 356 808 358 816
rect 366 808 368 816
rect 376 808 378 816
rect 396 808 398 816
rect 406 808 408 816
rect 426 808 428 816
rect 436 808 438 816
rect 456 808 458 816
rect 466 808 468 816
rect 486 808 488 816
rect 496 808 498 816
rect 516 808 518 816
rect 526 808 528 816
rect 546 808 548 816
rect 556 808 558 816
rect 576 808 578 816
rect 586 808 588 816
rect 596 808 600 816
rect 0 806 34 808
rect 42 806 64 808
rect 72 806 94 808
rect 102 806 124 808
rect 132 806 154 808
rect 162 806 184 808
rect 192 806 214 808
rect 222 806 378 808
rect 386 806 408 808
rect 416 806 438 808
rect 446 806 468 808
rect 476 806 498 808
rect 506 806 528 808
rect 536 806 558 808
rect 566 806 600 808
rect 0 798 4 806
rect 12 798 14 806
rect 22 798 24 806
rect 32 798 34 806
rect 52 798 54 806
rect 62 798 64 806
rect 82 798 84 806
rect 92 798 94 806
rect 112 798 114 806
rect 122 798 124 806
rect 142 798 144 806
rect 152 798 154 806
rect 172 798 174 806
rect 182 798 184 806
rect 202 798 204 806
rect 212 798 214 806
rect 232 798 234 806
rect 242 798 244 806
rect 262 798 264 806
rect 272 798 274 806
rect 282 798 286 806
rect 294 798 296 806
rect 304 798 306 806
rect 314 798 318 806
rect 326 798 328 806
rect 336 798 338 806
rect 356 798 358 806
rect 366 798 368 806
rect 386 798 388 806
rect 396 798 398 806
rect 416 798 418 806
rect 426 798 428 806
rect 446 798 448 806
rect 456 798 458 806
rect 476 798 478 806
rect 486 798 488 806
rect 506 798 508 806
rect 516 798 518 806
rect 536 798 538 806
rect 546 798 548 806
rect 566 798 568 806
rect 576 798 578 806
rect 586 798 588 806
rect 596 798 600 806
rect 0 796 34 798
rect 42 796 64 798
rect 72 796 94 798
rect 102 796 124 798
rect 132 796 154 798
rect 162 796 184 798
rect 192 796 214 798
rect 222 796 378 798
rect 386 796 408 798
rect 416 796 438 798
rect 446 796 468 798
rect 476 796 498 798
rect 506 796 528 798
rect 536 796 558 798
rect 566 796 600 798
rect 0 788 4 796
rect 12 788 14 796
rect 22 788 24 796
rect 42 788 44 796
rect 52 788 54 796
rect 72 788 74 796
rect 82 788 84 796
rect 102 788 104 796
rect 112 788 114 796
rect 132 788 134 796
rect 142 788 144 796
rect 162 788 164 796
rect 172 788 174 796
rect 192 788 194 796
rect 202 788 204 796
rect 222 788 224 796
rect 232 788 234 796
rect 242 788 244 796
rect 262 788 264 796
rect 272 788 276 796
rect 284 788 286 796
rect 294 788 296 796
rect 304 788 306 796
rect 314 788 316 796
rect 324 788 328 796
rect 336 788 338 796
rect 356 788 358 796
rect 366 788 368 796
rect 376 788 378 796
rect 396 788 398 796
rect 406 788 408 796
rect 426 788 428 796
rect 436 788 438 796
rect 456 788 458 796
rect 466 788 468 796
rect 486 788 488 796
rect 496 788 498 796
rect 516 788 518 796
rect 526 788 528 796
rect 546 788 548 796
rect 556 788 558 796
rect 576 788 578 796
rect 586 788 588 796
rect 596 788 600 796
rect 0 786 34 788
rect 42 786 64 788
rect 72 786 94 788
rect 102 786 124 788
rect 132 786 154 788
rect 162 786 184 788
rect 192 786 214 788
rect 222 786 378 788
rect 386 786 408 788
rect 416 786 438 788
rect 446 786 468 788
rect 476 786 498 788
rect 506 786 528 788
rect 536 786 558 788
rect 566 786 600 788
rect 0 778 4 786
rect 12 778 14 786
rect 22 778 24 786
rect 32 778 34 786
rect 52 778 54 786
rect 62 778 64 786
rect 82 778 84 786
rect 92 778 94 786
rect 0 776 34 778
rect 42 776 64 778
rect 72 776 94 778
rect 112 778 114 786
rect 122 778 124 786
rect 112 776 124 778
rect 142 778 144 786
rect 152 778 154 786
rect 142 776 154 778
rect 172 778 174 786
rect 182 778 184 786
rect 172 776 184 778
rect 202 778 204 786
rect 212 778 214 786
rect 202 776 214 778
rect 232 778 234 786
rect 242 778 244 786
rect 232 776 244 778
rect 262 778 264 786
rect 272 778 274 786
rect 262 776 274 778
rect 282 778 286 786
rect 294 778 296 786
rect 282 776 296 778
rect 0 768 4 776
rect 12 768 14 776
rect 22 768 24 776
rect 42 768 44 776
rect 52 768 54 776
rect 72 768 74 776
rect 82 768 84 776
rect 292 768 296 776
rect 0 766 34 768
rect 42 766 64 768
rect 72 766 94 768
rect 0 758 4 766
rect 12 758 14 766
rect 22 758 24 766
rect 32 758 34 766
rect 52 758 54 766
rect 62 758 64 766
rect 82 758 84 766
rect 92 758 94 766
rect 112 766 124 768
rect 112 758 114 766
rect 122 758 124 766
rect 142 766 154 768
rect 142 758 144 766
rect 152 758 154 766
rect 172 766 184 768
rect 172 758 174 766
rect 182 758 184 766
rect 202 766 214 768
rect 202 758 204 766
rect 212 758 214 766
rect 232 766 244 768
rect 232 758 234 766
rect 242 758 244 766
rect 262 766 274 768
rect 262 758 264 766
rect 272 758 274 766
rect 282 766 296 768
rect 282 758 286 766
rect 294 758 296 766
rect 304 778 306 786
rect 314 778 318 786
rect 304 776 318 778
rect 326 778 328 786
rect 336 778 338 786
rect 326 776 338 778
rect 356 778 358 786
rect 366 778 368 786
rect 356 776 368 778
rect 386 778 388 786
rect 396 778 398 786
rect 386 776 398 778
rect 416 778 418 786
rect 426 778 428 786
rect 416 776 428 778
rect 446 778 448 786
rect 456 778 458 786
rect 446 776 458 778
rect 476 778 478 786
rect 486 778 488 786
rect 476 776 488 778
rect 506 778 508 786
rect 516 778 518 786
rect 536 778 538 786
rect 546 778 548 786
rect 566 778 568 786
rect 576 778 578 786
rect 586 778 588 786
rect 596 778 600 786
rect 506 776 528 778
rect 536 776 558 778
rect 566 776 600 778
rect 304 768 308 776
rect 516 768 518 776
rect 526 768 528 776
rect 546 768 548 776
rect 556 768 558 776
rect 576 768 578 776
rect 586 768 588 776
rect 596 768 600 776
rect 304 766 318 768
rect 304 758 306 766
rect 314 758 318 766
rect 326 766 338 768
rect 326 758 328 766
rect 336 758 338 766
rect 356 766 368 768
rect 356 758 358 766
rect 366 758 368 766
rect 386 766 398 768
rect 386 758 388 766
rect 396 758 398 766
rect 416 766 428 768
rect 416 758 418 766
rect 426 758 428 766
rect 446 766 458 768
rect 446 758 448 766
rect 456 758 458 766
rect 476 766 488 768
rect 476 758 478 766
rect 486 758 488 766
rect 506 766 528 768
rect 536 766 558 768
rect 566 766 600 768
rect 506 758 508 766
rect 516 758 518 766
rect 536 758 538 766
rect 546 758 548 766
rect 566 758 568 766
rect 576 758 578 766
rect 586 758 588 766
rect 596 758 600 766
rect 0 756 34 758
rect 42 756 64 758
rect 72 756 94 758
rect 102 756 124 758
rect 132 756 154 758
rect 162 756 184 758
rect 192 756 214 758
rect 222 756 378 758
rect 386 756 408 758
rect 416 756 438 758
rect 446 756 468 758
rect 476 756 498 758
rect 506 756 528 758
rect 536 756 558 758
rect 566 756 600 758
rect 0 748 4 756
rect 12 748 14 756
rect 22 748 24 756
rect 42 748 44 756
rect 52 748 54 756
rect 72 748 74 756
rect 82 748 84 756
rect 102 748 104 756
rect 112 748 114 756
rect 132 748 134 756
rect 142 748 144 756
rect 162 748 164 756
rect 172 748 174 756
rect 192 748 194 756
rect 202 748 204 756
rect 222 748 224 756
rect 232 748 234 756
rect 242 748 244 756
rect 262 748 264 756
rect 272 748 274 756
rect 282 748 286 756
rect 294 748 296 756
rect 304 748 306 756
rect 314 748 318 756
rect 326 748 328 756
rect 336 748 338 756
rect 356 748 358 756
rect 366 748 368 756
rect 376 748 378 756
rect 396 748 398 756
rect 406 748 408 756
rect 426 748 428 756
rect 436 748 438 756
rect 456 748 458 756
rect 466 748 468 756
rect 486 748 488 756
rect 496 748 498 756
rect 516 748 518 756
rect 526 748 528 756
rect 546 748 548 756
rect 556 748 558 756
rect 576 748 578 756
rect 586 748 588 756
rect 596 748 600 756
rect 0 746 34 748
rect 42 746 64 748
rect 72 746 94 748
rect 102 746 124 748
rect 132 746 154 748
rect 162 746 184 748
rect 192 746 214 748
rect 222 746 378 748
rect 386 746 408 748
rect 416 746 438 748
rect 446 746 468 748
rect 476 746 498 748
rect 506 746 528 748
rect 536 746 558 748
rect 566 746 600 748
rect 0 738 4 746
rect 12 738 14 746
rect 22 738 24 746
rect 32 738 34 746
rect 52 738 54 746
rect 62 738 64 746
rect 82 738 84 746
rect 92 738 94 746
rect 112 738 114 746
rect 122 738 124 746
rect 142 738 144 746
rect 152 738 154 746
rect 172 738 174 746
rect 182 738 184 746
rect 202 738 204 746
rect 212 738 214 746
rect 232 738 234 746
rect 242 738 244 746
rect 262 738 264 746
rect 272 738 274 746
rect 282 738 286 746
rect 294 738 296 746
rect 304 738 306 746
rect 314 738 318 746
rect 326 738 328 746
rect 336 738 338 746
rect 356 738 358 746
rect 366 738 368 746
rect 386 738 388 746
rect 396 738 398 746
rect 416 738 418 746
rect 426 738 428 746
rect 446 738 448 746
rect 456 738 458 746
rect 476 738 478 746
rect 486 738 488 746
rect 506 738 508 746
rect 516 738 518 746
rect 536 738 538 746
rect 546 738 548 746
rect 566 738 568 746
rect 576 738 578 746
rect 586 738 588 746
rect 596 738 600 746
rect 0 737 214 738
rect 0 736 42 737
rect 0 728 4 736
rect 12 728 14 736
rect 22 728 24 736
rect 32 728 42 736
rect 0 727 42 728
rect 204 727 214 737
rect 0 726 214 727
rect 222 736 378 738
rect 222 728 224 736
rect 232 728 234 736
rect 242 728 244 736
rect 262 728 276 736
rect 284 728 286 736
rect 294 728 296 736
rect 304 728 306 736
rect 314 728 316 736
rect 324 728 338 736
rect 356 728 358 736
rect 366 728 368 736
rect 376 728 378 736
rect 222 726 378 728
rect 386 728 396 738
rect 560 736 600 738
rect 560 728 568 736
rect 576 728 578 736
rect 586 728 588 736
rect 596 728 600 736
rect 386 726 600 728
rect 0 718 4 726
rect 12 718 14 726
rect 22 718 24 726
rect 32 718 34 726
rect 52 718 54 726
rect 62 718 64 726
rect 82 718 84 726
rect 92 718 94 726
rect 112 718 114 726
rect 122 718 124 726
rect 142 718 144 726
rect 152 718 154 726
rect 172 718 174 726
rect 182 718 184 726
rect 202 718 204 726
rect 212 718 214 726
rect 232 718 234 726
rect 242 718 244 726
rect 262 718 264 726
rect 272 718 286 726
rect 294 718 296 726
rect 304 718 306 726
rect 314 718 328 726
rect 336 718 338 726
rect 356 718 358 726
rect 366 718 368 726
rect 386 718 388 726
rect 396 718 398 726
rect 416 718 418 726
rect 426 718 428 726
rect 446 718 448 726
rect 456 718 458 726
rect 476 718 478 726
rect 486 718 488 726
rect 506 718 508 726
rect 516 718 518 726
rect 536 718 538 726
rect 546 718 548 726
rect 566 718 568 726
rect 576 718 578 726
rect 586 718 588 726
rect 596 718 600 726
rect 0 716 34 718
rect 42 716 64 718
rect 72 716 94 718
rect 102 716 124 718
rect 132 716 154 718
rect 162 716 184 718
rect 192 716 214 718
rect 222 716 378 718
rect 386 716 408 718
rect 416 716 438 718
rect 446 716 468 718
rect 476 716 498 718
rect 506 716 528 718
rect 536 716 558 718
rect 566 716 600 718
rect 0 708 4 716
rect 12 708 14 716
rect 22 708 24 716
rect 42 708 44 716
rect 52 708 54 716
rect 72 708 74 716
rect 82 708 84 716
rect 102 708 104 716
rect 112 708 114 716
rect 132 708 134 716
rect 142 708 144 716
rect 162 708 164 716
rect 172 708 174 716
rect 192 708 194 716
rect 202 708 204 716
rect 222 708 224 716
rect 232 708 234 716
rect 242 708 244 716
rect 262 708 264 716
rect 272 708 276 716
rect 284 708 286 716
rect 294 708 296 716
rect 304 708 306 716
rect 314 708 316 716
rect 324 708 328 716
rect 336 708 338 716
rect 356 708 358 716
rect 366 708 368 716
rect 376 708 378 716
rect 396 708 398 716
rect 406 708 408 716
rect 426 708 428 716
rect 436 708 438 716
rect 456 708 458 716
rect 466 708 468 716
rect 486 708 488 716
rect 496 708 498 716
rect 516 708 518 716
rect 526 708 528 716
rect 546 708 548 716
rect 556 708 558 716
rect 576 708 578 716
rect 586 708 588 716
rect 596 708 600 716
rect 0 706 34 708
rect 42 706 64 708
rect 72 706 94 708
rect 102 706 124 708
rect 132 706 154 708
rect 162 706 184 708
rect 192 706 214 708
rect 222 706 378 708
rect 386 706 408 708
rect 416 706 438 708
rect 446 706 468 708
rect 476 706 498 708
rect 506 706 528 708
rect 536 706 558 708
rect 566 706 600 708
rect 0 698 4 706
rect 12 698 14 706
rect 22 698 24 706
rect 32 698 34 706
rect 52 698 54 706
rect 62 698 64 706
rect 82 698 84 706
rect 92 698 94 706
rect 112 698 114 706
rect 122 698 124 706
rect 142 698 144 706
rect 152 698 154 706
rect 172 698 174 706
rect 182 698 184 706
rect 202 698 204 706
rect 212 698 214 706
rect 232 698 234 706
rect 242 698 244 706
rect 262 698 264 706
rect 272 698 274 706
rect 282 698 286 706
rect 294 698 296 706
rect 304 698 306 706
rect 314 698 318 706
rect 326 698 328 706
rect 336 698 338 706
rect 356 698 358 706
rect 366 698 368 706
rect 386 698 388 706
rect 396 698 398 706
rect 416 698 418 706
rect 426 698 428 706
rect 446 698 448 706
rect 456 698 458 706
rect 476 698 478 706
rect 486 698 488 706
rect 506 698 508 706
rect 516 698 518 706
rect 536 698 538 706
rect 546 698 548 706
rect 566 698 568 706
rect 576 698 578 706
rect 586 698 588 706
rect 596 698 600 706
rect 0 696 34 698
rect 42 696 64 698
rect 72 696 94 698
rect 102 696 124 698
rect 132 696 154 698
rect 162 696 184 698
rect 192 696 214 698
rect 222 697 378 698
rect 222 696 286 697
rect 0 688 4 696
rect 12 688 14 696
rect 22 688 24 696
rect 42 688 44 696
rect 52 688 54 696
rect 72 688 74 696
rect 82 688 84 696
rect 102 688 104 696
rect 112 688 114 696
rect 132 688 134 696
rect 142 688 144 696
rect 162 688 164 696
rect 172 688 174 696
rect 192 688 194 696
rect 202 688 204 696
rect 222 688 224 696
rect 232 688 234 696
rect 242 688 244 696
rect 262 688 274 696
rect 282 689 286 696
rect 294 689 296 697
rect 304 689 306 697
rect 314 696 378 697
rect 386 696 408 698
rect 416 696 438 698
rect 446 696 468 698
rect 476 696 498 698
rect 506 696 528 698
rect 536 696 558 698
rect 566 696 600 698
rect 314 689 318 696
rect 282 688 318 689
rect 326 688 338 696
rect 356 688 358 696
rect 366 688 368 696
rect 376 688 378 696
rect 396 688 398 696
rect 406 688 408 696
rect 426 688 428 696
rect 436 688 438 696
rect 456 688 458 696
rect 466 688 468 696
rect 486 688 488 696
rect 496 688 498 696
rect 516 688 518 696
rect 526 688 528 696
rect 546 688 548 696
rect 556 688 558 696
rect 576 688 578 696
rect 586 688 588 696
rect 596 688 600 696
rect 204 658 396 688
rect 0 644 4 652
rect 12 644 14 652
rect 22 644 24 652
rect 42 644 44 652
rect 52 644 54 652
rect 72 644 74 652
rect 82 644 84 652
rect 102 644 104 652
rect 112 644 114 652
rect 132 644 134 652
rect 142 644 144 652
rect 162 644 164 652
rect 172 644 174 652
rect 0 642 34 644
rect 42 642 64 644
rect 72 642 94 644
rect 102 642 124 644
rect 132 642 154 644
rect 162 642 184 644
rect 0 634 4 642
rect 12 634 14 642
rect 22 634 24 642
rect 32 634 34 642
rect 52 634 54 642
rect 62 634 64 642
rect 82 634 84 642
rect 92 634 94 642
rect 112 634 114 642
rect 122 634 124 642
rect 142 634 144 642
rect 152 634 154 642
rect 172 634 174 642
rect 182 634 184 642
rect 0 632 34 634
rect 42 632 64 634
rect 72 632 94 634
rect 102 632 124 634
rect 132 632 154 634
rect 162 632 184 634
rect 0 624 4 632
rect 12 624 14 632
rect 22 624 24 632
rect 42 624 44 632
rect 52 624 54 632
rect 72 624 74 632
rect 82 624 84 632
rect 102 624 104 632
rect 112 624 114 632
rect 132 624 134 632
rect 142 624 144 632
rect 162 624 164 632
rect 172 624 174 632
rect 0 622 34 624
rect 42 622 64 624
rect 72 622 94 624
rect 102 622 124 624
rect 132 622 154 624
rect 162 622 184 624
rect 0 614 4 622
rect 12 614 14 622
rect 22 614 24 622
rect 32 614 34 622
rect 52 614 54 622
rect 62 614 64 622
rect 82 614 84 622
rect 92 614 94 622
rect 112 614 114 622
rect 122 614 124 622
rect 142 614 144 622
rect 152 614 154 622
rect 172 614 174 622
rect 182 614 184 622
rect 192 614 198 652
rect 0 612 198 614
rect 0 604 4 612
rect 12 604 14 612
rect 22 604 24 612
rect 32 604 40 612
rect 0 602 40 604
rect 0 594 4 602
rect 12 594 14 602
rect 22 594 24 602
rect 32 594 34 602
rect 52 594 54 602
rect 62 594 64 602
rect 82 594 84 602
rect 92 594 94 602
rect 112 594 114 602
rect 122 594 124 602
rect 142 594 144 602
rect 152 594 154 602
rect 172 594 174 602
rect 182 594 184 602
rect 0 592 34 594
rect 42 592 64 594
rect 72 592 94 594
rect 102 592 124 594
rect 132 592 154 594
rect 162 592 184 594
rect 0 584 4 592
rect 12 584 14 592
rect 22 584 24 592
rect 42 584 44 592
rect 52 584 54 592
rect 72 584 74 592
rect 82 584 84 592
rect 102 584 104 592
rect 112 584 114 592
rect 0 582 34 584
rect 42 582 64 584
rect 72 582 94 584
rect 102 582 114 584
rect 132 584 134 592
rect 142 584 144 592
rect 132 582 144 584
rect 162 584 164 592
rect 172 584 174 592
rect 162 582 174 584
rect 0 574 4 582
rect 12 574 14 582
rect 22 574 24 582
rect 32 574 34 582
rect 52 574 54 582
rect 62 574 64 582
rect 82 574 84 582
rect 92 574 94 582
rect 0 572 34 574
rect 42 572 64 574
rect 72 572 94 574
rect 102 572 114 574
rect 0 564 4 572
rect 12 564 14 572
rect 22 564 24 572
rect 42 564 44 572
rect 52 564 54 572
rect 72 564 74 572
rect 82 564 84 572
rect 102 564 104 572
rect 112 564 114 572
rect 132 572 144 574
rect 132 564 134 572
rect 142 564 144 572
rect 162 572 174 574
rect 162 564 164 572
rect 172 564 174 572
rect 0 562 34 564
rect 42 562 64 564
rect 72 562 94 564
rect 102 562 124 564
rect 132 562 154 564
rect 162 562 184 564
rect 0 554 4 562
rect 12 554 14 562
rect 22 554 24 562
rect 32 554 34 562
rect 52 554 54 562
rect 62 554 64 562
rect 82 554 84 562
rect 92 554 94 562
rect 112 554 114 562
rect 122 554 124 562
rect 142 554 144 562
rect 152 554 154 562
rect 172 554 174 562
rect 182 554 184 562
rect 0 552 34 554
rect 42 552 64 554
rect 72 552 94 554
rect 102 552 124 554
rect 132 552 154 554
rect 162 552 184 554
rect 0 544 4 552
rect 12 544 14 552
rect 22 544 24 552
rect 42 544 44 552
rect 52 544 54 552
rect 72 544 74 552
rect 82 544 84 552
rect 102 544 104 552
rect 112 544 114 552
rect 132 544 134 552
rect 142 544 144 552
rect 162 544 164 552
rect 172 544 174 552
rect 0 542 34 544
rect 42 542 64 544
rect 72 542 94 544
rect 102 542 124 544
rect 132 542 154 544
rect 162 542 184 544
rect 0 534 4 542
rect 12 534 14 542
rect 22 534 24 542
rect 32 534 34 542
rect 52 534 54 542
rect 62 534 64 542
rect 82 534 84 542
rect 92 534 94 542
rect 112 534 114 542
rect 122 534 124 542
rect 142 534 144 542
rect 152 534 154 542
rect 172 534 174 542
rect 182 534 184 542
rect 0 532 34 534
rect 42 532 64 534
rect 72 532 94 534
rect 102 532 124 534
rect 132 532 154 534
rect 162 532 184 534
rect 0 524 4 532
rect 12 524 14 532
rect 22 524 24 532
rect 42 524 44 532
rect 52 524 54 532
rect 72 524 74 532
rect 82 524 84 532
rect 102 524 104 532
rect 112 524 114 532
rect 132 524 134 532
rect 142 524 144 532
rect 162 524 164 532
rect 172 524 174 532
rect 192 524 198 602
rect 0 516 198 524
rect 0 512 14 516
rect 0 4 4 512
rect 12 508 14 512
rect 22 508 24 516
rect 32 508 34 516
rect 42 508 44 516
rect 52 508 54 516
rect 62 508 64 516
rect 72 508 74 516
rect 82 508 84 516
rect 92 508 94 516
rect 102 508 104 516
rect 112 508 114 516
rect 122 508 124 516
rect 132 508 134 516
rect 142 508 144 516
rect 152 508 154 516
rect 162 508 164 516
rect 172 508 174 516
rect 182 508 184 516
rect 192 508 198 516
rect 12 506 198 508
rect 12 14 14 506
rect 204 492 280 658
rect 286 644 290 652
rect 298 644 302 652
rect 310 644 314 652
rect 286 642 314 644
rect 286 632 314 634
rect 286 624 290 632
rect 298 624 302 632
rect 310 624 314 632
rect 286 622 314 624
rect 286 612 314 614
rect 286 604 290 612
rect 298 604 302 612
rect 310 604 314 612
rect 286 602 314 604
rect 286 586 290 594
rect 298 586 302 594
rect 310 586 314 594
rect 286 584 314 586
rect 286 564 314 566
rect 286 556 290 564
rect 298 556 302 564
rect 310 556 314 564
rect 286 554 314 556
rect 286 544 314 546
rect 286 536 290 544
rect 298 536 302 544
rect 310 536 314 544
rect 286 534 314 536
rect 286 524 314 526
rect 286 516 290 524
rect 298 516 302 524
rect 310 516 314 524
rect 286 514 314 516
rect 286 504 314 506
rect 320 492 396 658
rect 402 614 408 652
rect 426 644 428 652
rect 436 644 438 652
rect 456 644 458 652
rect 466 644 468 652
rect 486 644 488 652
rect 496 644 498 652
rect 516 644 518 652
rect 526 644 528 652
rect 546 644 548 652
rect 556 644 558 652
rect 576 644 578 652
rect 586 644 588 652
rect 596 644 600 652
rect 416 642 438 644
rect 446 642 468 644
rect 476 642 498 644
rect 506 642 528 644
rect 536 642 558 644
rect 566 642 600 644
rect 416 634 418 642
rect 426 634 428 642
rect 446 634 448 642
rect 456 634 458 642
rect 476 634 478 642
rect 486 634 488 642
rect 506 634 508 642
rect 516 634 518 642
rect 536 634 538 642
rect 546 634 548 642
rect 566 634 568 642
rect 576 634 578 642
rect 586 634 588 642
rect 596 634 600 642
rect 416 632 438 634
rect 446 632 468 634
rect 476 632 498 634
rect 506 632 528 634
rect 536 632 558 634
rect 566 632 600 634
rect 426 624 428 632
rect 436 624 438 632
rect 456 624 458 632
rect 466 624 468 632
rect 486 624 488 632
rect 496 624 498 632
rect 516 624 518 632
rect 526 624 528 632
rect 546 624 548 632
rect 556 624 558 632
rect 576 624 578 632
rect 586 624 588 632
rect 596 624 600 632
rect 416 622 438 624
rect 446 622 468 624
rect 476 622 498 624
rect 506 622 528 624
rect 536 622 558 624
rect 566 622 600 624
rect 416 614 418 622
rect 426 614 428 622
rect 446 614 448 622
rect 456 614 458 622
rect 476 614 478 622
rect 486 614 488 622
rect 506 614 508 622
rect 516 614 518 622
rect 536 614 538 622
rect 546 614 548 622
rect 566 614 568 622
rect 576 614 578 622
rect 586 614 588 622
rect 596 614 600 622
rect 402 612 600 614
rect 560 604 568 612
rect 576 604 578 612
rect 586 604 588 612
rect 596 604 600 612
rect 560 602 600 604
rect 402 524 408 602
rect 416 594 418 602
rect 426 594 428 602
rect 446 594 448 602
rect 456 594 458 602
rect 476 594 478 602
rect 486 594 488 602
rect 506 594 508 602
rect 516 594 518 602
rect 536 594 538 602
rect 546 594 548 602
rect 566 594 568 602
rect 576 594 578 602
rect 586 594 588 602
rect 596 594 600 602
rect 416 592 438 594
rect 446 592 468 594
rect 476 592 498 594
rect 506 592 528 594
rect 536 592 558 594
rect 566 592 600 594
rect 426 584 428 592
rect 436 584 438 592
rect 426 582 438 584
rect 456 584 458 592
rect 466 584 468 592
rect 456 582 468 584
rect 486 584 488 592
rect 496 584 498 592
rect 516 584 518 592
rect 526 584 528 592
rect 546 584 548 592
rect 556 584 558 592
rect 576 584 578 592
rect 586 584 588 592
rect 596 584 600 592
rect 486 582 498 584
rect 506 582 528 584
rect 536 582 558 584
rect 566 582 600 584
rect 506 574 508 582
rect 516 574 518 582
rect 536 574 538 582
rect 546 574 548 582
rect 566 574 568 582
rect 576 574 578 582
rect 586 574 588 582
rect 596 574 600 582
rect 426 572 438 574
rect 426 564 428 572
rect 436 564 438 572
rect 456 572 468 574
rect 456 564 458 572
rect 466 564 468 572
rect 486 572 498 574
rect 506 572 528 574
rect 536 572 558 574
rect 566 572 600 574
rect 486 564 488 572
rect 496 564 498 572
rect 516 564 518 572
rect 526 564 528 572
rect 546 564 548 572
rect 556 564 558 572
rect 576 564 578 572
rect 586 564 588 572
rect 596 564 600 572
rect 416 562 438 564
rect 446 562 468 564
rect 476 562 498 564
rect 506 562 528 564
rect 536 562 558 564
rect 566 562 600 564
rect 416 554 418 562
rect 426 554 428 562
rect 446 554 448 562
rect 456 554 458 562
rect 476 554 478 562
rect 486 554 488 562
rect 506 554 508 562
rect 516 554 518 562
rect 536 554 538 562
rect 546 554 548 562
rect 566 554 568 562
rect 576 554 578 562
rect 586 554 588 562
rect 596 554 600 562
rect 416 552 438 554
rect 446 552 468 554
rect 476 552 498 554
rect 506 552 528 554
rect 536 552 558 554
rect 566 552 600 554
rect 426 544 428 552
rect 436 544 438 552
rect 456 544 458 552
rect 466 544 468 552
rect 486 544 488 552
rect 496 544 498 552
rect 516 544 518 552
rect 526 544 528 552
rect 546 544 548 552
rect 556 544 558 552
rect 576 544 578 552
rect 586 544 588 552
rect 596 544 600 552
rect 416 542 438 544
rect 446 542 468 544
rect 476 542 498 544
rect 506 542 528 544
rect 536 542 558 544
rect 566 542 600 544
rect 416 534 418 542
rect 426 534 428 542
rect 446 534 448 542
rect 456 534 458 542
rect 476 534 478 542
rect 486 534 488 542
rect 506 534 508 542
rect 516 534 518 542
rect 536 534 538 542
rect 546 534 548 542
rect 566 534 568 542
rect 576 534 578 542
rect 586 534 588 542
rect 596 534 600 542
rect 416 532 438 534
rect 446 532 468 534
rect 476 532 498 534
rect 506 532 528 534
rect 536 532 558 534
rect 566 532 600 534
rect 426 524 428 532
rect 436 524 438 532
rect 456 524 458 532
rect 466 524 468 532
rect 486 524 488 532
rect 496 524 498 532
rect 516 524 518 532
rect 526 524 528 532
rect 546 524 548 532
rect 556 524 558 532
rect 576 524 578 532
rect 586 524 588 532
rect 596 524 600 532
rect 402 516 600 524
rect 402 508 408 516
rect 416 508 418 516
rect 426 508 428 516
rect 436 508 438 516
rect 446 508 448 516
rect 456 508 458 516
rect 466 508 468 516
rect 476 508 478 516
rect 486 508 488 516
rect 496 508 498 516
rect 506 508 508 516
rect 516 508 518 516
rect 526 508 528 516
rect 536 508 538 516
rect 546 508 548 516
rect 556 508 558 516
rect 566 508 568 516
rect 576 508 578 516
rect 586 512 600 516
rect 586 508 588 512
rect 402 506 588 508
rect 204 490 396 492
rect 30 489 570 490
rect 568 461 570 489
rect 30 459 40 461
rect 38 451 40 459
rect 48 459 60 461
rect 48 451 50 459
rect 58 451 60 459
rect 78 459 90 461
rect 78 451 80 459
rect 88 451 90 459
rect 108 459 120 461
rect 108 451 110 459
rect 118 451 120 459
rect 138 459 150 461
rect 138 451 140 459
rect 148 451 150 459
rect 168 459 180 461
rect 168 451 170 459
rect 178 451 180 459
rect 198 459 210 461
rect 198 451 200 459
rect 208 451 210 459
rect 228 459 240 461
rect 228 451 230 459
rect 238 451 240 459
rect 258 459 270 461
rect 258 451 260 459
rect 268 451 270 459
rect 288 459 300 461
rect 288 451 290 459
rect 298 451 300 459
rect 318 459 330 461
rect 318 451 320 459
rect 328 451 330 459
rect 348 459 360 461
rect 348 451 350 459
rect 358 451 360 459
rect 378 459 390 461
rect 378 451 380 459
rect 388 451 390 459
rect 408 459 420 461
rect 408 451 410 459
rect 418 451 420 459
rect 438 459 450 461
rect 438 451 440 459
rect 448 451 450 459
rect 468 459 480 461
rect 468 451 470 459
rect 478 451 480 459
rect 498 459 510 461
rect 498 451 500 459
rect 508 451 510 459
rect 528 459 540 461
rect 528 451 530 459
rect 538 451 540 459
rect 558 459 570 461
rect 558 451 560 459
rect 568 451 570 459
rect 30 449 60 451
rect 68 449 90 451
rect 98 449 120 451
rect 128 449 150 451
rect 158 449 180 451
rect 188 449 210 451
rect 218 449 240 451
rect 248 449 270 451
rect 278 449 300 451
rect 308 449 330 451
rect 338 449 360 451
rect 368 449 390 451
rect 398 449 420 451
rect 428 449 450 451
rect 458 449 480 451
rect 488 449 510 451
rect 518 449 540 451
rect 548 449 570 451
rect 38 441 40 449
rect 48 441 50 449
rect 68 441 70 449
rect 78 441 80 449
rect 98 441 100 449
rect 108 441 110 449
rect 128 441 130 449
rect 138 441 140 449
rect 158 441 160 449
rect 168 441 170 449
rect 188 441 190 449
rect 198 441 200 449
rect 218 441 220 449
rect 228 441 230 449
rect 248 441 250 449
rect 258 441 260 449
rect 278 441 280 449
rect 288 441 290 449
rect 308 441 310 449
rect 318 441 320 449
rect 338 441 340 449
rect 348 441 350 449
rect 368 441 370 449
rect 378 441 380 449
rect 398 441 400 449
rect 408 441 410 449
rect 428 441 430 449
rect 438 441 440 449
rect 458 441 460 449
rect 468 441 470 449
rect 488 441 490 449
rect 498 441 500 449
rect 518 441 520 449
rect 528 441 530 449
rect 548 441 550 449
rect 558 441 560 449
rect 568 441 570 449
rect 30 439 60 441
rect 68 439 90 441
rect 98 439 120 441
rect 128 439 150 441
rect 158 439 180 441
rect 188 439 210 441
rect 218 439 240 441
rect 248 439 270 441
rect 278 439 300 441
rect 308 439 330 441
rect 338 439 360 441
rect 368 439 390 441
rect 398 439 420 441
rect 428 439 450 441
rect 458 439 480 441
rect 488 439 510 441
rect 518 439 540 441
rect 548 439 570 441
rect 38 431 40 439
rect 48 431 50 439
rect 58 431 60 439
rect 78 431 80 439
rect 88 431 90 439
rect 108 431 110 439
rect 118 431 120 439
rect 138 431 140 439
rect 148 431 150 439
rect 168 431 170 439
rect 178 431 180 439
rect 198 431 200 439
rect 208 431 210 439
rect 228 431 230 439
rect 238 431 240 439
rect 258 431 260 439
rect 268 431 270 439
rect 288 431 290 439
rect 298 431 300 439
rect 318 431 320 439
rect 328 431 330 439
rect 348 431 350 439
rect 358 431 360 439
rect 378 431 380 439
rect 388 431 390 439
rect 408 431 410 439
rect 418 431 420 439
rect 438 431 440 439
rect 448 431 450 439
rect 468 431 470 439
rect 478 431 480 439
rect 498 431 500 439
rect 508 431 510 439
rect 528 431 530 439
rect 538 431 540 439
rect 558 431 560 439
rect 568 431 570 439
rect 30 429 60 431
rect 68 429 90 431
rect 98 429 120 431
rect 128 429 150 431
rect 158 429 180 431
rect 188 429 210 431
rect 218 429 240 431
rect 248 429 270 431
rect 278 429 300 431
rect 308 429 330 431
rect 338 429 360 431
rect 368 429 390 431
rect 398 429 420 431
rect 428 429 450 431
rect 458 429 480 431
rect 488 429 510 431
rect 518 429 540 431
rect 548 429 570 431
rect 38 421 40 429
rect 48 421 50 429
rect 68 421 70 429
rect 78 421 80 429
rect 98 421 100 429
rect 108 421 110 429
rect 128 421 130 429
rect 138 421 140 429
rect 158 421 160 429
rect 168 421 170 429
rect 188 421 190 429
rect 198 421 200 429
rect 218 421 220 429
rect 228 421 230 429
rect 248 421 250 429
rect 258 421 260 429
rect 278 421 280 429
rect 288 421 290 429
rect 308 421 310 429
rect 318 421 320 429
rect 338 421 340 429
rect 348 421 350 429
rect 368 421 370 429
rect 378 421 380 429
rect 398 421 400 429
rect 408 421 410 429
rect 428 421 430 429
rect 438 421 440 429
rect 458 421 460 429
rect 468 421 470 429
rect 488 421 490 429
rect 498 421 500 429
rect 518 421 520 429
rect 528 421 530 429
rect 548 421 550 429
rect 558 421 560 429
rect 568 421 570 429
rect 30 419 60 421
rect 68 419 90 421
rect 98 419 120 421
rect 128 419 150 421
rect 158 419 180 421
rect 188 419 210 421
rect 218 419 240 421
rect 248 419 270 421
rect 278 419 300 421
rect 308 419 330 421
rect 338 419 360 421
rect 368 419 390 421
rect 398 419 420 421
rect 428 419 450 421
rect 458 419 480 421
rect 488 419 510 421
rect 518 419 540 421
rect 548 419 570 421
rect 38 411 40 419
rect 48 411 50 419
rect 58 411 60 419
rect 78 411 80 419
rect 88 411 90 419
rect 108 411 110 419
rect 118 411 120 419
rect 138 411 140 419
rect 148 411 150 419
rect 168 411 170 419
rect 178 411 180 419
rect 198 411 200 419
rect 208 411 210 419
rect 228 411 230 419
rect 238 411 240 419
rect 258 411 260 419
rect 268 411 270 419
rect 288 411 290 419
rect 298 411 300 419
rect 318 411 320 419
rect 328 411 330 419
rect 348 411 350 419
rect 358 411 360 419
rect 378 411 380 419
rect 388 411 390 419
rect 408 411 410 419
rect 418 411 420 419
rect 438 411 440 419
rect 448 411 450 419
rect 468 411 470 419
rect 478 411 480 419
rect 498 411 500 419
rect 508 411 510 419
rect 528 411 530 419
rect 538 411 540 419
rect 558 411 560 419
rect 568 411 570 419
rect 30 409 60 411
rect 68 409 90 411
rect 98 409 120 411
rect 128 409 150 411
rect 158 409 180 411
rect 188 409 210 411
rect 218 409 240 411
rect 248 409 270 411
rect 278 409 300 411
rect 308 409 330 411
rect 338 409 360 411
rect 368 409 390 411
rect 398 409 420 411
rect 428 409 450 411
rect 458 409 480 411
rect 488 409 510 411
rect 518 409 540 411
rect 548 409 570 411
rect 38 401 40 409
rect 48 401 50 409
rect 68 401 70 409
rect 78 401 80 409
rect 98 401 100 409
rect 108 401 110 409
rect 128 401 130 409
rect 138 401 140 409
rect 158 401 160 409
rect 168 401 170 409
rect 188 401 190 409
rect 198 401 200 409
rect 218 401 220 409
rect 228 401 230 409
rect 248 401 250 409
rect 258 401 260 409
rect 278 401 280 409
rect 288 401 290 409
rect 308 401 310 409
rect 318 401 320 409
rect 338 401 340 409
rect 348 401 350 409
rect 368 401 370 409
rect 378 401 380 409
rect 398 401 400 409
rect 408 401 410 409
rect 428 401 430 409
rect 438 401 440 409
rect 458 401 460 409
rect 468 401 470 409
rect 488 401 490 409
rect 498 401 500 409
rect 518 401 520 409
rect 528 401 530 409
rect 548 401 550 409
rect 558 401 560 409
rect 568 401 570 409
rect 30 399 60 401
rect 68 399 90 401
rect 98 399 120 401
rect 128 399 150 401
rect 158 399 180 401
rect 188 399 210 401
rect 218 399 240 401
rect 248 399 270 401
rect 278 399 300 401
rect 308 399 330 401
rect 338 399 360 401
rect 368 399 390 401
rect 398 399 420 401
rect 428 399 450 401
rect 458 399 480 401
rect 488 399 510 401
rect 518 399 540 401
rect 548 399 570 401
rect 38 371 40 399
rect 48 371 50 399
rect 58 371 60 399
rect 78 371 80 399
rect 88 371 90 399
rect 108 391 110 399
rect 118 391 120 399
rect 138 391 140 399
rect 148 391 150 399
rect 168 391 170 399
rect 178 391 180 399
rect 198 391 200 399
rect 208 391 210 399
rect 228 391 230 399
rect 238 391 240 399
rect 258 391 260 399
rect 268 391 270 399
rect 288 391 290 399
rect 298 391 300 399
rect 318 391 320 399
rect 328 391 330 399
rect 348 391 350 399
rect 358 391 360 399
rect 378 391 380 399
rect 388 391 390 399
rect 408 391 410 399
rect 418 391 420 399
rect 438 391 440 399
rect 448 391 450 399
rect 468 391 470 399
rect 478 391 480 399
rect 498 391 500 399
rect 98 390 500 391
rect 98 380 100 390
rect 204 380 396 390
rect 98 379 500 380
rect 108 371 110 379
rect 118 371 120 379
rect 138 371 140 379
rect 148 371 150 379
rect 168 371 170 379
rect 178 371 180 379
rect 198 371 200 379
rect 208 371 210 379
rect 228 371 230 379
rect 238 371 240 379
rect 258 371 260 379
rect 268 371 270 379
rect 288 371 290 379
rect 298 371 300 379
rect 318 371 320 379
rect 328 371 330 379
rect 348 371 350 379
rect 358 371 360 379
rect 378 371 380 379
rect 388 371 390 379
rect 408 371 410 379
rect 418 371 420 379
rect 438 371 440 379
rect 448 371 450 379
rect 468 371 470 379
rect 478 371 480 379
rect 498 371 500 379
rect 508 371 510 399
rect 528 391 530 399
rect 538 391 540 399
rect 558 391 560 399
rect 568 391 570 399
rect 518 389 540 391
rect 548 389 570 391
rect 518 381 520 389
rect 528 381 530 389
rect 548 381 550 389
rect 558 381 560 389
rect 568 381 570 389
rect 518 379 540 381
rect 548 379 570 381
rect 528 371 530 379
rect 538 371 540 379
rect 558 371 560 379
rect 568 371 570 379
rect 30 369 60 371
rect 68 369 90 371
rect 98 369 120 371
rect 128 369 150 371
rect 158 369 180 371
rect 188 369 210 371
rect 218 369 240 371
rect 248 369 270 371
rect 278 369 300 371
rect 308 369 330 371
rect 338 369 360 371
rect 368 369 390 371
rect 398 369 420 371
rect 428 369 450 371
rect 458 369 480 371
rect 488 369 510 371
rect 518 369 540 371
rect 548 369 570 371
rect 38 361 40 369
rect 48 361 50 369
rect 68 361 70 369
rect 78 361 80 369
rect 98 361 100 369
rect 108 361 110 369
rect 128 361 130 369
rect 138 361 140 369
rect 158 361 160 369
rect 168 361 170 369
rect 188 361 190 369
rect 198 361 200 369
rect 218 361 220 369
rect 228 361 230 369
rect 248 361 250 369
rect 258 361 260 369
rect 278 361 280 369
rect 288 361 290 369
rect 308 361 310 369
rect 318 361 320 369
rect 338 361 340 369
rect 348 361 350 369
rect 368 361 370 369
rect 378 361 380 369
rect 398 361 400 369
rect 408 361 410 369
rect 428 361 430 369
rect 438 361 440 369
rect 458 361 460 369
rect 468 361 470 369
rect 488 361 490 369
rect 498 361 500 369
rect 518 361 520 369
rect 528 361 530 369
rect 548 361 550 369
rect 558 361 560 369
rect 568 361 570 369
rect 30 359 60 361
rect 68 359 90 361
rect 98 359 120 361
rect 128 359 150 361
rect 158 359 180 361
rect 188 359 210 361
rect 218 359 240 361
rect 248 359 270 361
rect 278 359 300 361
rect 308 359 330 361
rect 338 359 360 361
rect 368 359 390 361
rect 398 359 420 361
rect 428 359 450 361
rect 458 359 480 361
rect 488 359 510 361
rect 518 359 540 361
rect 548 359 570 361
rect 38 351 40 359
rect 48 351 50 359
rect 58 351 60 359
rect 78 351 80 359
rect 88 351 90 359
rect 108 351 110 359
rect 118 351 120 359
rect 138 351 140 359
rect 148 351 150 359
rect 168 351 170 359
rect 178 351 180 359
rect 198 351 200 359
rect 208 351 210 359
rect 228 351 230 359
rect 238 351 240 359
rect 258 351 260 359
rect 268 351 270 359
rect 288 351 290 359
rect 298 351 300 359
rect 318 351 320 359
rect 328 351 330 359
rect 348 351 350 359
rect 358 351 360 359
rect 378 351 380 359
rect 388 351 390 359
rect 408 351 410 359
rect 418 351 420 359
rect 438 351 440 359
rect 448 351 450 359
rect 468 351 470 359
rect 478 351 480 359
rect 498 351 500 359
rect 508 351 510 359
rect 528 351 530 359
rect 538 351 540 359
rect 558 351 560 359
rect 568 351 570 359
rect 30 349 60 351
rect 68 349 90 351
rect 98 349 120 351
rect 128 349 150 351
rect 158 349 180 351
rect 188 349 210 351
rect 218 349 240 351
rect 248 349 270 351
rect 278 349 300 351
rect 308 349 330 351
rect 338 349 360 351
rect 368 349 390 351
rect 398 349 420 351
rect 428 349 450 351
rect 458 349 480 351
rect 488 349 510 351
rect 518 349 540 351
rect 548 349 570 351
rect 38 341 40 349
rect 48 341 50 349
rect 68 341 70 349
rect 78 341 80 349
rect 98 341 100 349
rect 108 341 110 349
rect 128 341 130 349
rect 138 341 140 349
rect 158 341 160 349
rect 168 341 170 349
rect 188 341 190 349
rect 198 341 200 349
rect 218 341 220 349
rect 228 341 230 349
rect 248 341 250 349
rect 258 341 260 349
rect 278 341 280 349
rect 288 341 290 349
rect 308 341 310 349
rect 318 341 320 349
rect 338 341 340 349
rect 348 341 350 349
rect 368 341 370 349
rect 378 341 380 349
rect 398 341 400 349
rect 408 341 410 349
rect 428 341 430 349
rect 438 341 440 349
rect 458 341 460 349
rect 468 341 470 349
rect 488 341 490 349
rect 498 341 500 349
rect 518 341 520 349
rect 528 341 530 349
rect 548 341 550 349
rect 558 341 560 349
rect 568 341 570 349
rect 30 339 60 341
rect 68 339 90 341
rect 98 339 120 341
rect 128 339 150 341
rect 158 339 180 341
rect 188 339 210 341
rect 218 339 240 341
rect 248 339 270 341
rect 278 339 300 341
rect 308 339 330 341
rect 338 339 360 341
rect 368 339 390 341
rect 398 339 420 341
rect 428 339 450 341
rect 458 339 480 341
rect 488 339 510 341
rect 518 339 540 341
rect 548 339 570 341
rect 38 331 40 339
rect 48 331 50 339
rect 58 331 60 339
rect 78 331 80 339
rect 88 331 90 339
rect 108 331 110 339
rect 118 331 120 339
rect 138 331 140 339
rect 148 331 150 339
rect 168 331 170 339
rect 178 331 180 339
rect 198 331 200 339
rect 208 331 210 339
rect 228 331 230 339
rect 238 331 240 339
rect 258 331 260 339
rect 268 331 270 339
rect 288 331 290 339
rect 298 331 300 339
rect 318 331 320 339
rect 328 331 330 339
rect 348 331 350 339
rect 358 331 360 339
rect 378 331 380 339
rect 388 331 390 339
rect 408 331 410 339
rect 418 331 420 339
rect 438 331 440 339
rect 448 331 450 339
rect 468 331 470 339
rect 478 331 480 339
rect 498 331 500 339
rect 508 331 510 339
rect 528 331 530 339
rect 538 331 540 339
rect 558 331 560 339
rect 568 331 570 339
rect 30 329 60 331
rect 68 329 90 331
rect 98 329 120 331
rect 128 329 150 331
rect 158 329 180 331
rect 188 329 210 331
rect 218 329 240 331
rect 248 329 270 331
rect 278 329 300 331
rect 308 329 330 331
rect 338 329 360 331
rect 368 329 390 331
rect 398 329 420 331
rect 428 329 450 331
rect 458 329 480 331
rect 488 329 510 331
rect 518 329 540 331
rect 548 329 570 331
rect 38 321 40 329
rect 48 321 50 329
rect 68 321 70 329
rect 78 321 80 329
rect 98 321 100 329
rect 108 321 110 329
rect 128 321 130 329
rect 138 321 140 329
rect 158 321 160 329
rect 168 321 170 329
rect 188 321 190 329
rect 198 321 200 329
rect 218 321 220 329
rect 228 321 230 329
rect 248 321 250 329
rect 258 321 260 329
rect 278 321 280 329
rect 288 321 290 329
rect 308 321 310 329
rect 318 321 320 329
rect 338 321 340 329
rect 348 321 350 329
rect 368 321 370 329
rect 378 321 380 329
rect 398 321 400 329
rect 408 321 410 329
rect 428 321 430 329
rect 438 321 440 329
rect 458 321 460 329
rect 468 321 470 329
rect 488 321 490 329
rect 498 321 500 329
rect 518 321 520 329
rect 528 321 530 329
rect 548 321 550 329
rect 558 321 560 329
rect 568 321 570 329
rect 30 319 60 321
rect 68 319 90 321
rect 98 319 120 321
rect 128 319 150 321
rect 158 319 180 321
rect 188 319 210 321
rect 218 319 240 321
rect 248 319 270 321
rect 278 319 300 321
rect 308 319 330 321
rect 338 319 360 321
rect 368 319 390 321
rect 398 319 420 321
rect 428 319 450 321
rect 458 319 480 321
rect 488 319 510 321
rect 518 319 540 321
rect 548 319 570 321
rect 38 311 40 319
rect 48 311 50 319
rect 58 311 60 319
rect 78 311 80 319
rect 88 311 90 319
rect 108 311 110 319
rect 118 311 120 319
rect 138 311 140 319
rect 148 311 150 319
rect 168 311 170 319
rect 178 311 180 319
rect 198 311 200 319
rect 208 311 210 319
rect 228 311 230 319
rect 238 311 240 319
rect 258 311 260 319
rect 268 311 270 319
rect 288 311 290 319
rect 298 311 300 319
rect 318 311 320 319
rect 328 311 330 319
rect 348 311 350 319
rect 358 311 360 319
rect 378 311 380 319
rect 388 311 390 319
rect 408 311 410 319
rect 418 311 420 319
rect 438 311 440 319
rect 448 311 450 319
rect 468 311 470 319
rect 478 311 480 319
rect 498 311 500 319
rect 508 311 510 319
rect 528 311 530 319
rect 538 311 540 319
rect 558 311 560 319
rect 568 311 570 319
rect 30 309 60 311
rect 68 309 510 311
rect 518 309 540 311
rect 548 309 570 311
rect 38 301 40 309
rect 48 301 50 309
rect 68 301 70 309
rect 78 301 80 309
rect 88 301 90 309
rect 98 301 500 309
rect 518 301 520 309
rect 528 301 530 309
rect 548 301 550 309
rect 558 301 560 309
rect 568 301 570 309
rect 30 299 60 301
rect 68 299 510 301
rect 518 299 540 301
rect 548 299 570 301
rect 38 291 40 299
rect 48 291 50 299
rect 58 291 60 299
rect 78 291 80 299
rect 88 291 90 299
rect 108 291 110 299
rect 118 291 120 299
rect 138 291 140 299
rect 148 291 150 299
rect 168 291 170 299
rect 178 291 180 299
rect 198 291 200 299
rect 208 291 210 299
rect 228 291 230 299
rect 238 291 240 299
rect 258 291 260 299
rect 268 291 270 299
rect 288 291 290 299
rect 298 291 300 299
rect 318 291 320 299
rect 328 291 330 299
rect 348 291 350 299
rect 358 291 360 299
rect 378 291 380 299
rect 388 291 390 299
rect 408 291 410 299
rect 418 291 420 299
rect 438 291 440 299
rect 448 291 450 299
rect 468 291 470 299
rect 478 291 480 299
rect 498 291 500 299
rect 508 291 510 299
rect 528 291 530 299
rect 538 291 540 299
rect 558 291 560 299
rect 568 291 570 299
rect 30 289 60 291
rect 68 289 90 291
rect 98 289 120 291
rect 128 289 150 291
rect 158 289 180 291
rect 188 289 210 291
rect 218 289 240 291
rect 248 289 270 291
rect 278 289 300 291
rect 308 289 330 291
rect 338 289 360 291
rect 368 289 390 291
rect 398 289 420 291
rect 428 289 450 291
rect 458 289 480 291
rect 488 289 510 291
rect 518 289 540 291
rect 548 289 570 291
rect 38 281 40 289
rect 48 281 50 289
rect 68 281 70 289
rect 78 281 80 289
rect 98 281 100 289
rect 108 281 110 289
rect 128 281 130 289
rect 138 281 140 289
rect 158 281 160 289
rect 168 281 170 289
rect 188 281 190 289
rect 198 281 200 289
rect 218 281 220 289
rect 228 281 230 289
rect 248 281 250 289
rect 258 281 260 289
rect 278 281 280 289
rect 288 281 290 289
rect 308 281 310 289
rect 318 281 320 289
rect 338 281 340 289
rect 348 281 350 289
rect 368 281 370 289
rect 378 281 380 289
rect 398 281 400 289
rect 408 281 410 289
rect 428 281 430 289
rect 438 281 440 289
rect 458 281 460 289
rect 468 281 470 289
rect 488 281 490 289
rect 498 281 500 289
rect 518 281 520 289
rect 528 281 530 289
rect 548 281 550 289
rect 558 281 560 289
rect 568 281 570 289
rect 30 279 60 281
rect 68 279 90 281
rect 98 279 120 281
rect 128 279 150 281
rect 158 279 180 281
rect 188 279 210 281
rect 218 279 240 281
rect 248 279 270 281
rect 278 279 300 281
rect 308 279 330 281
rect 338 279 360 281
rect 368 279 390 281
rect 398 279 420 281
rect 428 279 450 281
rect 458 279 480 281
rect 488 279 510 281
rect 518 279 540 281
rect 548 279 570 281
rect 38 271 40 279
rect 48 271 50 279
rect 58 271 60 279
rect 78 271 80 279
rect 88 271 90 279
rect 108 271 110 279
rect 118 271 120 279
rect 138 271 140 279
rect 148 271 150 279
rect 168 271 170 279
rect 178 271 180 279
rect 198 271 200 279
rect 208 271 210 279
rect 228 271 230 279
rect 238 271 240 279
rect 258 271 260 279
rect 268 271 270 279
rect 288 271 290 279
rect 298 271 300 279
rect 318 271 320 279
rect 328 271 330 279
rect 348 271 350 279
rect 358 271 360 279
rect 378 271 380 279
rect 388 271 390 279
rect 408 271 410 279
rect 418 271 420 279
rect 438 271 440 279
rect 448 271 450 279
rect 468 271 470 279
rect 478 271 480 279
rect 498 271 500 279
rect 508 271 510 279
rect 528 271 530 279
rect 538 271 540 279
rect 558 271 560 279
rect 568 271 570 279
rect 30 269 60 271
rect 68 269 90 271
rect 98 269 120 271
rect 128 269 150 271
rect 158 269 180 271
rect 188 269 210 271
rect 218 269 240 271
rect 248 269 270 271
rect 278 269 300 271
rect 308 269 330 271
rect 338 269 360 271
rect 368 269 390 271
rect 398 269 420 271
rect 428 269 450 271
rect 458 269 480 271
rect 488 269 510 271
rect 518 269 540 271
rect 548 269 570 271
rect 38 261 40 269
rect 48 261 50 269
rect 68 261 70 269
rect 78 261 80 269
rect 98 261 100 269
rect 108 261 110 269
rect 128 261 130 269
rect 138 261 140 269
rect 158 261 160 269
rect 168 261 170 269
rect 188 261 190 269
rect 198 261 200 269
rect 218 261 220 269
rect 228 261 230 269
rect 248 261 250 269
rect 258 261 260 269
rect 278 261 280 269
rect 288 261 290 269
rect 308 261 310 269
rect 318 261 320 269
rect 338 261 340 269
rect 348 261 350 269
rect 368 261 370 269
rect 378 261 380 269
rect 398 261 400 269
rect 408 261 410 269
rect 428 261 430 269
rect 438 261 440 269
rect 458 261 460 269
rect 468 261 470 269
rect 488 261 490 269
rect 498 261 500 269
rect 518 261 520 269
rect 528 261 530 269
rect 548 261 550 269
rect 558 261 560 269
rect 568 261 570 269
rect 30 259 60 261
rect 68 259 90 261
rect 98 259 120 261
rect 128 259 150 261
rect 158 259 180 261
rect 188 259 210 261
rect 218 259 240 261
rect 248 259 270 261
rect 278 259 300 261
rect 308 259 330 261
rect 338 259 360 261
rect 368 259 390 261
rect 398 259 420 261
rect 428 259 450 261
rect 458 259 480 261
rect 488 259 510 261
rect 518 259 540 261
rect 548 259 570 261
rect 38 251 40 259
rect 48 251 50 259
rect 58 251 60 259
rect 78 251 80 259
rect 88 251 90 259
rect 108 251 110 259
rect 118 251 120 259
rect 138 251 140 259
rect 148 251 150 259
rect 168 251 170 259
rect 178 251 180 259
rect 198 251 200 259
rect 208 251 210 259
rect 228 251 230 259
rect 238 251 240 259
rect 258 251 260 259
rect 268 251 270 259
rect 288 251 290 259
rect 298 251 300 259
rect 318 251 320 259
rect 328 251 330 259
rect 348 251 350 259
rect 358 251 360 259
rect 378 251 380 259
rect 388 251 390 259
rect 408 251 410 259
rect 418 251 420 259
rect 438 251 440 259
rect 448 251 450 259
rect 468 251 470 259
rect 478 251 480 259
rect 498 251 500 259
rect 508 251 510 259
rect 528 251 530 259
rect 538 251 540 259
rect 558 251 560 259
rect 568 251 570 259
rect 30 249 60 251
rect 68 249 90 251
rect 98 249 120 251
rect 128 249 150 251
rect 158 249 180 251
rect 188 249 210 251
rect 218 249 240 251
rect 248 249 270 251
rect 278 249 300 251
rect 308 249 330 251
rect 338 249 360 251
rect 368 249 390 251
rect 398 249 420 251
rect 428 249 450 251
rect 458 249 480 251
rect 488 249 510 251
rect 518 249 540 251
rect 548 249 570 251
rect 38 241 40 249
rect 48 241 50 249
rect 30 239 60 241
rect 38 231 40 239
rect 48 231 50 239
rect 58 231 60 239
rect 30 229 60 231
rect 38 221 40 229
rect 48 221 50 229
rect 68 221 70 249
rect 78 221 80 249
rect 98 241 100 249
rect 108 241 110 249
rect 128 241 130 249
rect 138 241 140 249
rect 158 241 160 249
rect 168 241 170 249
rect 188 241 190 249
rect 198 241 200 249
rect 218 241 220 249
rect 228 241 230 249
rect 248 241 250 249
rect 258 241 260 249
rect 278 241 280 249
rect 288 241 290 249
rect 308 241 310 249
rect 318 241 320 249
rect 338 241 340 249
rect 348 241 350 249
rect 368 241 370 249
rect 378 241 380 249
rect 398 241 400 249
rect 408 241 410 249
rect 428 241 430 249
rect 438 241 440 249
rect 458 241 460 249
rect 468 241 470 249
rect 488 241 490 249
rect 498 241 500 249
rect 518 241 520 249
rect 528 241 530 249
rect 548 241 550 249
rect 558 241 560 249
rect 568 241 570 249
rect 88 240 500 241
rect 88 230 100 240
rect 204 230 396 240
rect 88 229 500 230
rect 508 239 540 241
rect 548 239 570 241
rect 508 231 510 239
rect 518 231 520 239
rect 528 231 530 239
rect 538 231 540 239
rect 558 231 560 239
rect 568 231 570 239
rect 508 229 540 231
rect 548 229 570 231
rect 98 221 100 229
rect 108 221 110 229
rect 128 221 130 229
rect 138 221 140 229
rect 158 221 160 229
rect 168 221 170 229
rect 188 221 190 229
rect 198 221 200 229
rect 218 221 220 229
rect 228 221 230 229
rect 248 221 250 229
rect 258 221 260 229
rect 278 221 280 229
rect 288 221 290 229
rect 308 221 310 229
rect 318 221 320 229
rect 338 221 340 229
rect 348 221 350 229
rect 368 221 370 229
rect 378 221 380 229
rect 398 221 400 229
rect 408 221 410 229
rect 428 221 430 229
rect 438 221 440 229
rect 458 221 460 229
rect 468 221 470 229
rect 488 221 490 229
rect 498 221 500 229
rect 518 221 520 229
rect 528 221 530 229
rect 548 221 550 229
rect 558 221 560 229
rect 568 221 570 229
rect 30 219 60 221
rect 68 219 90 221
rect 98 219 120 221
rect 128 219 150 221
rect 158 219 180 221
rect 188 219 210 221
rect 218 219 240 221
rect 248 219 270 221
rect 278 219 300 221
rect 308 219 330 221
rect 338 219 360 221
rect 368 219 390 221
rect 398 219 420 221
rect 428 219 450 221
rect 458 219 480 221
rect 488 219 510 221
rect 518 219 540 221
rect 548 219 570 221
rect 38 211 40 219
rect 48 211 50 219
rect 58 211 60 219
rect 78 211 80 219
rect 88 211 90 219
rect 108 211 110 219
rect 118 211 120 219
rect 138 211 140 219
rect 148 211 150 219
rect 168 211 170 219
rect 178 211 180 219
rect 198 211 200 219
rect 208 211 210 219
rect 228 211 230 219
rect 238 211 240 219
rect 258 211 260 219
rect 268 211 270 219
rect 288 211 290 219
rect 298 211 300 219
rect 318 211 320 219
rect 328 211 330 219
rect 348 211 350 219
rect 358 211 360 219
rect 378 211 380 219
rect 388 211 390 219
rect 408 211 410 219
rect 418 211 420 219
rect 438 211 440 219
rect 448 211 450 219
rect 468 211 470 219
rect 478 211 480 219
rect 498 211 500 219
rect 508 211 510 219
rect 528 211 530 219
rect 538 211 540 219
rect 558 211 560 219
rect 568 211 570 219
rect 30 209 60 211
rect 68 209 90 211
rect 98 209 120 211
rect 128 209 150 211
rect 158 209 180 211
rect 188 209 210 211
rect 218 209 240 211
rect 248 209 270 211
rect 278 209 300 211
rect 308 209 330 211
rect 338 209 360 211
rect 368 209 390 211
rect 398 209 420 211
rect 428 209 450 211
rect 458 209 480 211
rect 488 209 510 211
rect 518 209 540 211
rect 548 209 570 211
rect 38 201 40 209
rect 48 201 50 209
rect 68 201 70 209
rect 78 201 80 209
rect 98 201 100 209
rect 108 201 110 209
rect 128 201 130 209
rect 138 201 140 209
rect 158 201 160 209
rect 168 201 170 209
rect 188 201 190 209
rect 198 201 200 209
rect 218 201 220 209
rect 228 201 230 209
rect 248 201 250 209
rect 258 201 260 209
rect 278 201 280 209
rect 288 201 290 209
rect 308 201 310 209
rect 318 201 320 209
rect 338 201 340 209
rect 348 201 350 209
rect 368 201 370 209
rect 378 201 380 209
rect 398 201 400 209
rect 408 201 410 209
rect 428 201 430 209
rect 438 201 440 209
rect 458 201 460 209
rect 468 201 470 209
rect 488 201 490 209
rect 498 201 500 209
rect 518 201 520 209
rect 528 201 530 209
rect 548 201 550 209
rect 558 201 560 209
rect 568 201 570 209
rect 30 199 60 201
rect 68 199 90 201
rect 98 199 120 201
rect 128 199 150 201
rect 158 199 180 201
rect 188 199 210 201
rect 218 199 240 201
rect 248 199 270 201
rect 278 199 300 201
rect 308 199 330 201
rect 338 199 360 201
rect 368 199 390 201
rect 398 199 420 201
rect 428 199 450 201
rect 458 199 480 201
rect 488 199 510 201
rect 518 199 540 201
rect 548 199 570 201
rect 38 191 40 199
rect 48 191 50 199
rect 58 191 60 199
rect 78 191 80 199
rect 88 191 90 199
rect 108 191 110 199
rect 118 191 120 199
rect 138 191 140 199
rect 148 191 150 199
rect 168 191 170 199
rect 178 191 180 199
rect 198 191 200 199
rect 208 191 210 199
rect 228 191 230 199
rect 238 191 240 199
rect 258 191 260 199
rect 268 191 270 199
rect 288 191 290 199
rect 298 191 300 199
rect 318 191 320 199
rect 328 191 330 199
rect 348 191 350 199
rect 358 191 360 199
rect 378 191 380 199
rect 388 191 390 199
rect 408 191 410 199
rect 418 191 420 199
rect 438 191 440 199
rect 448 191 450 199
rect 468 191 470 199
rect 478 191 480 199
rect 498 191 500 199
rect 508 191 510 199
rect 528 191 530 199
rect 538 191 540 199
rect 558 191 560 199
rect 568 191 570 199
rect 30 189 60 191
rect 68 189 90 191
rect 98 189 120 191
rect 128 189 150 191
rect 158 189 180 191
rect 188 189 210 191
rect 218 189 240 191
rect 248 189 270 191
rect 278 189 300 191
rect 308 189 330 191
rect 338 189 360 191
rect 368 189 390 191
rect 398 189 420 191
rect 428 189 450 191
rect 458 189 480 191
rect 488 189 510 191
rect 518 189 540 191
rect 548 189 570 191
rect 38 181 40 189
rect 48 181 50 189
rect 68 181 70 189
rect 78 181 80 189
rect 98 181 100 189
rect 108 181 110 189
rect 128 181 130 189
rect 138 181 140 189
rect 158 181 160 189
rect 168 181 170 189
rect 188 181 190 189
rect 198 181 200 189
rect 218 181 220 189
rect 228 181 230 189
rect 248 181 250 189
rect 258 181 260 189
rect 278 181 280 189
rect 288 181 290 189
rect 308 181 310 189
rect 318 181 320 189
rect 338 181 340 189
rect 348 181 350 189
rect 368 181 370 189
rect 378 181 380 189
rect 398 181 400 189
rect 408 181 410 189
rect 428 181 430 189
rect 438 181 440 189
rect 458 181 460 189
rect 468 181 470 189
rect 488 181 490 189
rect 498 181 500 189
rect 518 181 520 189
rect 528 181 530 189
rect 548 181 550 189
rect 558 181 560 189
rect 568 181 570 189
rect 30 179 60 181
rect 68 179 90 181
rect 98 179 120 181
rect 128 179 150 181
rect 158 179 180 181
rect 188 179 210 181
rect 218 179 240 181
rect 248 179 270 181
rect 278 179 300 181
rect 308 179 330 181
rect 338 179 360 181
rect 368 179 390 181
rect 398 179 420 181
rect 428 179 450 181
rect 458 179 480 181
rect 488 179 510 181
rect 518 179 540 181
rect 548 179 570 181
rect 38 171 40 179
rect 48 171 50 179
rect 58 171 60 179
rect 78 171 80 179
rect 88 171 90 179
rect 108 171 110 179
rect 118 171 120 179
rect 138 171 140 179
rect 148 171 150 179
rect 168 171 170 179
rect 178 171 180 179
rect 198 171 200 179
rect 208 171 210 179
rect 228 171 230 179
rect 238 171 240 179
rect 258 171 260 179
rect 268 171 270 179
rect 288 171 290 179
rect 298 171 300 179
rect 318 171 320 179
rect 328 171 330 179
rect 348 171 350 179
rect 358 171 360 179
rect 378 171 380 179
rect 388 171 390 179
rect 408 171 410 179
rect 418 171 420 179
rect 438 171 440 179
rect 448 171 450 179
rect 468 171 470 179
rect 478 171 480 179
rect 498 171 500 179
rect 508 171 510 179
rect 528 171 530 179
rect 538 171 540 179
rect 558 171 560 179
rect 568 171 570 179
rect 30 169 60 171
rect 68 169 90 171
rect 98 169 120 171
rect 128 169 150 171
rect 158 169 180 171
rect 188 169 210 171
rect 218 169 240 171
rect 248 169 270 171
rect 278 169 300 171
rect 308 169 330 171
rect 338 169 360 171
rect 368 169 390 171
rect 398 169 420 171
rect 428 169 450 171
rect 458 169 480 171
rect 488 169 510 171
rect 518 169 540 171
rect 548 169 570 171
rect 38 161 40 169
rect 48 161 50 169
rect 68 161 70 169
rect 78 161 80 169
rect 98 161 100 169
rect 108 161 110 169
rect 128 161 130 169
rect 138 161 140 169
rect 158 161 160 169
rect 168 161 170 169
rect 188 161 190 169
rect 198 161 200 169
rect 218 161 220 169
rect 228 161 230 169
rect 248 161 250 169
rect 258 161 260 169
rect 278 161 280 169
rect 288 161 290 169
rect 308 161 310 169
rect 318 161 320 169
rect 338 161 340 169
rect 348 161 350 169
rect 368 161 370 169
rect 378 161 380 169
rect 398 161 400 169
rect 408 161 410 169
rect 428 161 430 169
rect 438 161 440 169
rect 458 161 460 169
rect 468 161 470 169
rect 488 161 490 169
rect 498 161 500 169
rect 518 161 520 169
rect 528 161 530 169
rect 548 161 550 169
rect 558 161 560 169
rect 568 161 570 169
rect 30 159 60 161
rect 68 159 90 161
rect 38 151 40 159
rect 48 151 50 159
rect 58 151 60 159
rect 78 151 80 159
rect 88 151 90 159
rect 30 149 60 151
rect 68 149 90 151
rect 98 149 500 161
rect 508 159 540 161
rect 548 159 570 161
rect 508 151 510 159
rect 518 151 520 159
rect 528 151 530 159
rect 538 151 540 159
rect 558 151 560 159
rect 568 151 570 159
rect 508 149 540 151
rect 548 149 570 151
rect 38 141 40 149
rect 48 141 50 149
rect 68 141 70 149
rect 78 141 80 149
rect 98 141 100 149
rect 108 141 110 149
rect 128 141 130 149
rect 138 141 140 149
rect 158 141 160 149
rect 168 141 170 149
rect 188 141 190 149
rect 198 141 200 149
rect 218 141 220 149
rect 228 141 230 149
rect 248 141 250 149
rect 258 141 260 149
rect 278 141 280 149
rect 288 141 290 149
rect 308 141 310 149
rect 318 141 320 149
rect 338 141 340 149
rect 348 141 350 149
rect 368 141 370 149
rect 378 141 380 149
rect 398 141 400 149
rect 408 141 410 149
rect 428 141 430 149
rect 438 141 440 149
rect 458 141 460 149
rect 468 141 470 149
rect 488 141 490 149
rect 498 141 500 149
rect 518 141 520 149
rect 528 141 530 149
rect 548 141 550 149
rect 558 141 560 149
rect 568 141 570 149
rect 30 139 60 141
rect 68 139 90 141
rect 98 139 120 141
rect 128 139 150 141
rect 158 139 180 141
rect 188 139 210 141
rect 218 139 240 141
rect 248 139 270 141
rect 278 139 300 141
rect 308 139 330 141
rect 338 139 360 141
rect 368 139 390 141
rect 398 139 420 141
rect 428 139 450 141
rect 458 139 480 141
rect 488 139 510 141
rect 518 139 540 141
rect 548 139 570 141
rect 38 131 40 139
rect 48 131 50 139
rect 58 131 60 139
rect 78 131 80 139
rect 88 131 90 139
rect 108 131 110 139
rect 118 131 120 139
rect 138 131 140 139
rect 148 131 150 139
rect 168 131 170 139
rect 178 131 180 139
rect 198 131 200 139
rect 208 131 210 139
rect 228 131 230 139
rect 238 131 240 139
rect 258 131 260 139
rect 268 131 270 139
rect 288 131 290 139
rect 298 131 300 139
rect 318 131 320 139
rect 328 131 330 139
rect 348 131 350 139
rect 358 131 360 139
rect 378 131 380 139
rect 388 131 390 139
rect 408 131 410 139
rect 418 131 420 139
rect 438 131 440 139
rect 448 131 450 139
rect 468 131 470 139
rect 478 131 480 139
rect 498 131 500 139
rect 508 131 510 139
rect 528 131 530 139
rect 538 131 540 139
rect 558 131 560 139
rect 568 131 570 139
rect 30 129 60 131
rect 68 129 90 131
rect 98 129 120 131
rect 128 129 150 131
rect 158 129 180 131
rect 188 129 210 131
rect 218 129 240 131
rect 248 129 270 131
rect 278 129 300 131
rect 308 129 330 131
rect 338 129 360 131
rect 368 129 390 131
rect 398 129 420 131
rect 428 129 450 131
rect 458 129 480 131
rect 488 129 510 131
rect 518 129 540 131
rect 548 129 570 131
rect 38 121 40 129
rect 48 121 50 129
rect 68 121 70 129
rect 78 121 80 129
rect 98 121 100 129
rect 108 121 110 129
rect 128 121 130 129
rect 138 121 140 129
rect 158 121 160 129
rect 168 121 170 129
rect 188 121 190 129
rect 198 121 200 129
rect 218 121 220 129
rect 228 121 230 129
rect 248 121 250 129
rect 258 121 260 129
rect 278 121 280 129
rect 288 121 290 129
rect 308 121 310 129
rect 318 121 320 129
rect 338 121 340 129
rect 348 121 350 129
rect 368 121 370 129
rect 378 121 380 129
rect 398 121 400 129
rect 408 121 410 129
rect 428 121 430 129
rect 438 121 440 129
rect 458 121 460 129
rect 468 121 470 129
rect 488 121 490 129
rect 498 121 500 129
rect 518 121 520 129
rect 528 121 530 129
rect 548 121 550 129
rect 558 121 560 129
rect 568 121 570 129
rect 30 119 60 121
rect 68 119 90 121
rect 98 119 120 121
rect 128 119 150 121
rect 158 119 180 121
rect 188 119 210 121
rect 218 119 240 121
rect 248 119 270 121
rect 278 119 300 121
rect 308 119 330 121
rect 338 119 360 121
rect 368 119 390 121
rect 398 119 420 121
rect 428 119 450 121
rect 458 119 480 121
rect 488 119 510 121
rect 518 119 540 121
rect 548 119 570 121
rect 38 111 40 119
rect 48 111 50 119
rect 58 111 60 119
rect 78 111 80 119
rect 88 111 90 119
rect 108 111 110 119
rect 118 111 120 119
rect 138 111 140 119
rect 148 111 150 119
rect 168 111 170 119
rect 178 111 180 119
rect 198 111 200 119
rect 208 111 210 119
rect 228 111 230 119
rect 238 111 240 119
rect 258 111 260 119
rect 268 111 270 119
rect 288 111 290 119
rect 298 111 300 119
rect 318 111 320 119
rect 328 111 330 119
rect 348 111 350 119
rect 358 111 360 119
rect 378 111 380 119
rect 388 111 390 119
rect 408 111 410 119
rect 418 111 420 119
rect 438 111 440 119
rect 448 111 450 119
rect 468 111 470 119
rect 478 111 480 119
rect 498 111 500 119
rect 508 111 510 119
rect 528 111 530 119
rect 538 111 540 119
rect 558 111 560 119
rect 568 111 570 119
rect 30 109 60 111
rect 68 109 90 111
rect 98 109 120 111
rect 128 109 150 111
rect 158 109 180 111
rect 188 109 210 111
rect 218 109 240 111
rect 248 109 270 111
rect 278 109 300 111
rect 308 109 330 111
rect 338 109 360 111
rect 368 109 390 111
rect 398 109 420 111
rect 428 109 450 111
rect 458 109 480 111
rect 488 109 510 111
rect 518 109 540 111
rect 548 109 570 111
rect 38 101 40 109
rect 48 101 50 109
rect 68 101 70 109
rect 78 101 80 109
rect 98 101 100 109
rect 108 101 110 109
rect 128 101 130 109
rect 138 101 140 109
rect 158 101 160 109
rect 168 101 170 109
rect 188 101 190 109
rect 198 101 200 109
rect 218 101 220 109
rect 228 101 230 109
rect 248 101 250 109
rect 258 101 260 109
rect 278 101 280 109
rect 288 101 290 109
rect 308 101 310 109
rect 318 101 320 109
rect 338 101 340 109
rect 348 101 350 109
rect 368 101 370 109
rect 378 101 380 109
rect 398 101 400 109
rect 408 101 410 109
rect 428 101 430 109
rect 438 101 440 109
rect 458 101 460 109
rect 468 101 470 109
rect 488 101 490 109
rect 498 101 500 109
rect 518 101 520 109
rect 528 101 530 109
rect 548 101 550 109
rect 558 101 560 109
rect 568 101 570 109
rect 30 99 60 101
rect 68 99 90 101
rect 98 99 120 101
rect 128 99 150 101
rect 158 99 180 101
rect 188 99 210 101
rect 218 99 240 101
rect 248 99 270 101
rect 278 99 300 101
rect 308 99 330 101
rect 338 99 360 101
rect 368 99 390 101
rect 398 99 420 101
rect 428 99 450 101
rect 458 99 480 101
rect 488 99 510 101
rect 518 99 540 101
rect 548 99 570 101
rect 38 91 40 99
rect 48 91 50 99
rect 58 91 60 99
rect 78 91 80 99
rect 88 91 90 99
rect 108 91 110 99
rect 118 91 120 99
rect 138 91 140 99
rect 148 91 150 99
rect 168 91 170 99
rect 178 91 180 99
rect 198 91 200 99
rect 208 91 210 99
rect 228 91 230 99
rect 238 91 240 99
rect 258 91 260 99
rect 268 91 270 99
rect 288 91 290 99
rect 298 91 300 99
rect 318 91 320 99
rect 328 91 330 99
rect 348 91 350 99
rect 358 91 360 99
rect 378 91 380 99
rect 388 91 390 99
rect 408 91 410 99
rect 418 91 420 99
rect 438 91 440 99
rect 448 91 450 99
rect 468 91 470 99
rect 478 91 480 99
rect 498 91 500 99
rect 508 91 510 99
rect 528 91 530 99
rect 538 91 540 99
rect 558 91 560 99
rect 568 91 570 99
rect 30 89 60 91
rect 68 89 90 91
rect 98 89 120 91
rect 128 89 150 91
rect 158 89 180 91
rect 188 89 210 91
rect 218 89 240 91
rect 248 89 270 91
rect 278 89 300 91
rect 308 89 330 91
rect 338 89 360 91
rect 368 89 390 91
rect 398 89 420 91
rect 428 89 450 91
rect 458 89 480 91
rect 488 89 510 91
rect 518 89 540 91
rect 548 89 570 91
rect 38 81 40 89
rect 48 81 50 89
rect 68 81 70 89
rect 78 81 80 89
rect 98 81 100 89
rect 108 81 110 89
rect 128 81 130 89
rect 138 81 140 89
rect 158 81 160 89
rect 168 81 170 89
rect 188 81 190 89
rect 198 81 200 89
rect 218 81 220 89
rect 228 81 230 89
rect 248 81 250 89
rect 258 81 260 89
rect 278 81 280 89
rect 288 81 290 89
rect 308 81 310 89
rect 318 81 320 89
rect 338 81 340 89
rect 348 81 350 89
rect 368 81 370 89
rect 378 81 380 89
rect 398 81 400 89
rect 408 81 410 89
rect 428 81 430 89
rect 438 81 440 89
rect 458 81 460 89
rect 468 81 470 89
rect 488 81 490 89
rect 498 81 500 89
rect 518 81 520 89
rect 528 81 530 89
rect 548 81 550 89
rect 558 81 560 89
rect 568 81 570 89
rect 30 79 60 81
rect 68 79 90 81
rect 98 79 120 81
rect 128 79 150 81
rect 158 79 180 81
rect 188 79 210 81
rect 218 79 240 81
rect 248 79 270 81
rect 278 79 300 81
rect 308 79 330 81
rect 338 79 360 81
rect 368 79 390 81
rect 398 79 420 81
rect 428 79 450 81
rect 458 79 480 81
rect 488 79 510 81
rect 518 79 540 81
rect 548 79 570 81
rect 38 71 40 79
rect 48 71 50 79
rect 58 71 60 79
rect 78 71 80 79
rect 88 71 90 79
rect 108 71 110 79
rect 118 71 120 79
rect 138 71 140 79
rect 148 71 150 79
rect 168 71 170 79
rect 178 71 180 79
rect 198 71 200 79
rect 208 71 210 79
rect 228 71 230 79
rect 238 71 240 79
rect 258 71 260 79
rect 268 71 270 79
rect 288 71 290 79
rect 298 71 300 79
rect 318 71 320 79
rect 328 71 330 79
rect 348 71 350 79
rect 358 71 360 79
rect 378 71 380 79
rect 388 71 390 79
rect 408 71 410 79
rect 418 71 420 79
rect 438 71 440 79
rect 448 71 450 79
rect 468 71 470 79
rect 478 71 480 79
rect 498 71 500 79
rect 508 71 510 79
rect 528 71 530 79
rect 538 71 540 79
rect 558 71 560 79
rect 568 71 570 79
rect 30 69 60 71
rect 68 69 90 71
rect 98 69 120 71
rect 128 69 150 71
rect 158 69 180 71
rect 188 69 210 71
rect 218 69 240 71
rect 248 69 270 71
rect 278 69 300 71
rect 308 69 330 71
rect 338 69 360 71
rect 368 69 390 71
rect 398 69 420 71
rect 428 69 450 71
rect 458 69 480 71
rect 488 69 510 71
rect 518 69 540 71
rect 548 69 570 71
rect 38 61 40 69
rect 48 61 50 69
rect 68 61 70 69
rect 78 61 80 69
rect 98 61 100 69
rect 108 61 110 69
rect 128 61 130 69
rect 138 61 140 69
rect 158 61 160 69
rect 168 61 170 69
rect 188 61 190 69
rect 198 61 200 69
rect 218 61 220 69
rect 228 61 230 69
rect 248 61 250 69
rect 258 61 260 69
rect 278 61 280 69
rect 288 61 290 69
rect 308 61 310 69
rect 318 61 320 69
rect 338 61 340 69
rect 348 61 350 69
rect 368 61 370 69
rect 378 61 380 69
rect 398 61 400 69
rect 408 61 410 69
rect 428 61 430 69
rect 438 61 440 69
rect 458 61 460 69
rect 468 61 470 69
rect 488 61 490 69
rect 498 61 500 69
rect 518 61 520 69
rect 528 61 530 69
rect 548 61 550 69
rect 558 61 560 69
rect 568 61 570 69
rect 30 59 60 61
rect 68 59 90 61
rect 98 59 120 61
rect 128 59 150 61
rect 158 59 180 61
rect 188 59 210 61
rect 218 59 240 61
rect 248 59 270 61
rect 278 59 300 61
rect 308 59 330 61
rect 338 59 360 61
rect 368 59 390 61
rect 398 59 420 61
rect 428 59 450 61
rect 458 59 480 61
rect 488 59 510 61
rect 518 59 540 61
rect 548 59 570 61
rect 38 51 40 59
rect 48 51 50 59
rect 58 51 60 59
rect 78 51 80 59
rect 88 51 90 59
rect 108 51 110 59
rect 118 51 120 59
rect 138 51 140 59
rect 148 51 150 59
rect 168 51 170 59
rect 178 51 180 59
rect 198 51 200 59
rect 208 51 210 59
rect 228 51 230 59
rect 238 51 240 59
rect 258 51 260 59
rect 268 51 270 59
rect 288 51 290 59
rect 298 51 300 59
rect 318 51 320 59
rect 328 51 330 59
rect 348 51 350 59
rect 358 51 360 59
rect 378 51 380 59
rect 388 51 390 59
rect 408 51 410 59
rect 418 51 420 59
rect 438 51 440 59
rect 448 51 450 59
rect 468 51 470 59
rect 478 51 480 59
rect 498 51 500 59
rect 508 51 510 59
rect 528 51 530 59
rect 538 51 540 59
rect 558 51 560 59
rect 568 51 570 59
rect 30 49 60 51
rect 68 49 90 51
rect 98 49 120 51
rect 128 49 150 51
rect 158 49 180 51
rect 188 49 210 51
rect 218 49 240 51
rect 248 49 270 51
rect 278 49 300 51
rect 308 49 330 51
rect 338 49 360 51
rect 368 49 390 51
rect 398 49 420 51
rect 428 49 450 51
rect 458 49 480 51
rect 488 49 510 51
rect 518 49 540 51
rect 548 49 570 51
rect 38 41 40 49
rect 48 41 50 49
rect 68 41 70 49
rect 78 41 80 49
rect 98 41 100 49
rect 108 41 110 49
rect 128 41 130 49
rect 138 41 140 49
rect 158 41 160 49
rect 168 41 170 49
rect 188 41 190 49
rect 198 41 200 49
rect 218 41 220 49
rect 228 41 230 49
rect 248 41 250 49
rect 258 41 260 49
rect 278 41 280 49
rect 288 41 290 49
rect 308 41 310 49
rect 318 41 320 49
rect 338 41 340 49
rect 348 41 350 49
rect 368 41 370 49
rect 378 41 380 49
rect 398 41 400 49
rect 408 41 410 49
rect 428 41 430 49
rect 438 41 440 49
rect 458 41 460 49
rect 468 41 470 49
rect 488 41 490 49
rect 498 41 500 49
rect 518 41 520 49
rect 528 41 530 49
rect 548 41 550 49
rect 558 41 560 49
rect 568 41 570 49
rect 30 39 60 41
rect 68 39 90 41
rect 98 39 120 41
rect 128 39 150 41
rect 158 39 180 41
rect 188 39 210 41
rect 218 39 240 41
rect 248 39 270 41
rect 278 39 300 41
rect 308 39 330 41
rect 338 39 360 41
rect 368 39 390 41
rect 398 39 420 41
rect 428 39 450 41
rect 458 39 480 41
rect 488 39 510 41
rect 518 39 540 41
rect 548 39 570 41
rect 38 31 40 39
rect 48 31 50 39
rect 58 31 60 39
rect 78 31 80 39
rect 88 31 90 39
rect 108 31 110 39
rect 118 31 120 39
rect 138 31 140 39
rect 148 31 150 39
rect 168 31 170 39
rect 178 31 180 39
rect 198 31 200 39
rect 208 31 210 39
rect 228 31 230 39
rect 238 31 240 39
rect 258 31 260 39
rect 268 31 270 39
rect 288 31 290 39
rect 298 31 300 39
rect 318 31 320 39
rect 328 31 330 39
rect 348 31 350 39
rect 358 31 360 39
rect 378 31 380 39
rect 388 31 390 39
rect 408 31 410 39
rect 418 31 420 39
rect 438 31 440 39
rect 448 31 450 39
rect 468 31 470 39
rect 478 31 480 39
rect 498 31 500 39
rect 508 31 510 39
rect 528 31 530 39
rect 538 31 540 39
rect 558 31 560 39
rect 568 31 570 39
rect 30 30 570 31
rect 12 12 198 14
rect 192 4 198 12
rect 0 2 198 4
rect 204 12 396 30
rect 586 14 588 506
rect 204 4 206 12
rect 394 4 396 12
rect 204 0 396 4
rect 402 12 588 14
rect 402 4 408 12
rect 596 4 600 512
rect 402 2 600 4
<< m2contact >>
rect 42 1290 50 1298
rect 62 1290 70 1298
rect 50 1279 58 1287
rect 72 1284 80 1290
rect 92 1286 100 1294
rect 112 1286 120 1294
rect 132 1286 140 1294
rect 152 1286 160 1294
rect 172 1286 180 1294
rect 192 1286 200 1294
rect 212 1286 220 1294
rect 232 1286 240 1294
rect 72 1282 90 1284
rect 42 1270 50 1278
rect 82 1276 90 1282
rect 102 1276 110 1284
rect 122 1276 130 1284
rect 142 1276 150 1284
rect 162 1276 170 1284
rect 182 1276 190 1284
rect 202 1276 210 1284
rect 222 1276 230 1284
rect 50 1259 58 1267
rect 42 1250 50 1258
rect 50 1239 58 1247
rect 42 1230 50 1238
rect 50 1219 58 1227
rect 42 1210 50 1218
rect 50 1199 58 1207
rect 42 1190 50 1198
rect 50 1179 58 1187
rect 42 1170 50 1178
rect 50 1159 58 1167
rect 42 1150 50 1158
rect 50 1139 58 1147
rect 42 1130 50 1138
rect 50 1119 58 1127
rect 42 1110 50 1118
rect 50 1099 58 1107
rect 42 1090 50 1098
rect 50 1079 58 1087
rect 42 1070 50 1078
rect 50 1059 58 1067
rect 42 1050 50 1058
rect 50 1039 58 1047
rect 42 1030 50 1038
rect 50 1019 58 1027
rect 42 1010 50 1018
rect 50 999 58 1007
rect 42 990 50 998
rect 50 979 58 987
rect 42 970 50 978
rect 50 959 58 967
rect 42 950 50 958
rect 50 939 58 947
rect 42 930 50 938
rect 50 919 58 927
rect 42 910 50 918
rect 78 1242 236 1250
rect 78 1180 96 1242
rect 360 1286 368 1294
rect 380 1286 388 1294
rect 400 1286 408 1294
rect 420 1286 428 1294
rect 440 1286 448 1294
rect 460 1286 468 1294
rect 480 1286 488 1294
rect 500 1286 508 1294
rect 530 1290 538 1298
rect 550 1290 558 1298
rect 520 1284 528 1290
rect 370 1276 378 1284
rect 390 1276 398 1284
rect 410 1276 418 1284
rect 430 1276 438 1284
rect 450 1276 458 1284
rect 470 1276 478 1284
rect 490 1276 498 1284
rect 510 1282 528 1284
rect 510 1276 518 1282
rect 542 1279 550 1287
rect 550 1270 558 1278
rect 542 1259 550 1267
rect 364 1242 522 1250
rect 78 1172 236 1180
rect 78 1114 236 1122
rect 290 1212 298 1220
rect 302 1212 310 1220
rect 290 1192 298 1200
rect 302 1192 310 1200
rect 504 1180 522 1242
rect 78 1052 96 1114
rect 364 1172 522 1180
rect 364 1114 522 1122
rect 78 1044 236 1052
rect 78 984 236 992
rect 290 1084 298 1092
rect 302 1084 310 1092
rect 290 1064 298 1072
rect 302 1064 310 1072
rect 504 1052 522 1114
rect 78 922 96 984
rect 364 1044 522 1052
rect 364 984 522 992
rect 78 914 236 922
rect 50 899 58 907
rect 42 890 50 898
rect 50 880 58 888
rect 290 954 298 962
rect 302 954 310 962
rect 290 934 298 942
rect 302 934 310 942
rect 504 922 522 984
rect 364 914 522 922
rect 550 1250 558 1258
rect 542 1239 550 1247
rect 550 1230 558 1238
rect 542 1219 550 1227
rect 550 1210 558 1218
rect 542 1199 550 1207
rect 550 1190 558 1198
rect 542 1179 550 1187
rect 550 1170 558 1178
rect 542 1159 550 1167
rect 550 1150 558 1158
rect 542 1139 550 1147
rect 550 1130 558 1138
rect 542 1119 550 1127
rect 550 1110 558 1118
rect 542 1099 550 1107
rect 550 1090 558 1098
rect 542 1079 550 1087
rect 550 1070 558 1078
rect 542 1059 550 1067
rect 550 1050 558 1058
rect 542 1039 550 1047
rect 550 1030 558 1038
rect 542 1019 550 1027
rect 550 1010 558 1018
rect 542 999 550 1007
rect 550 990 558 998
rect 542 979 550 987
rect 550 970 558 978
rect 542 959 550 967
rect 550 950 558 958
rect 542 939 550 947
rect 550 930 558 938
rect 542 919 550 927
rect 550 910 558 918
rect 542 899 550 907
rect 550 890 558 898
rect 542 880 550 888
rect 24 836 42 844
rect 14 828 22 836
rect 44 828 52 836
rect 54 836 72 844
rect 74 828 82 836
rect 84 836 102 844
rect 104 828 112 836
rect 114 836 132 844
rect 134 828 142 836
rect 144 836 162 844
rect 164 828 172 836
rect 174 836 192 844
rect 194 828 202 836
rect 204 836 222 844
rect 224 828 232 836
rect 234 836 242 844
rect 244 828 262 836
rect 264 836 272 844
rect 274 828 282 836
rect 286 836 294 844
rect 296 828 304 836
rect 306 836 314 844
rect 318 828 326 836
rect 328 836 336 844
rect 338 828 356 836
rect 358 836 366 844
rect 368 828 376 836
rect 378 836 396 844
rect 398 828 406 836
rect 408 836 426 844
rect 428 828 436 836
rect 438 836 456 844
rect 458 828 466 836
rect 468 836 486 844
rect 488 828 496 836
rect 498 836 516 844
rect 518 828 526 836
rect 528 836 546 844
rect 548 828 556 836
rect 558 836 576 844
rect 578 828 586 836
rect 4 818 12 826
rect 24 818 32 826
rect 54 818 62 826
rect 84 818 92 826
rect 114 818 122 826
rect 144 818 152 826
rect 174 818 182 826
rect 204 818 212 826
rect 234 818 242 826
rect 264 818 272 826
rect 286 818 294 826
rect 306 818 314 826
rect 328 818 336 826
rect 358 818 366 826
rect 388 818 396 826
rect 418 818 426 826
rect 448 818 456 826
rect 478 818 486 826
rect 508 818 516 826
rect 538 818 546 826
rect 568 818 576 826
rect 588 818 596 826
rect 14 808 22 816
rect 44 808 52 816
rect 74 808 82 816
rect 104 808 112 816
rect 134 808 142 816
rect 164 808 172 816
rect 194 808 202 816
rect 224 808 232 816
rect 244 808 262 816
rect 276 808 284 816
rect 296 808 304 816
rect 316 808 324 816
rect 338 808 356 816
rect 368 808 376 816
rect 398 808 406 816
rect 428 808 436 816
rect 458 808 466 816
rect 488 808 496 816
rect 518 808 526 816
rect 548 808 556 816
rect 578 808 586 816
rect 4 798 12 806
rect 24 798 32 806
rect 54 798 62 806
rect 84 798 92 806
rect 114 798 122 806
rect 144 798 152 806
rect 174 798 182 806
rect 204 798 212 806
rect 234 798 242 806
rect 264 798 272 806
rect 286 798 294 806
rect 306 798 314 806
rect 328 798 336 806
rect 358 798 366 806
rect 388 798 396 806
rect 418 798 426 806
rect 448 798 456 806
rect 478 798 486 806
rect 508 798 516 806
rect 538 798 546 806
rect 568 798 576 806
rect 588 798 596 806
rect 14 788 22 796
rect 44 788 52 796
rect 74 788 82 796
rect 104 788 112 796
rect 134 788 142 796
rect 164 788 172 796
rect 194 788 202 796
rect 224 788 232 796
rect 244 788 262 796
rect 276 788 284 796
rect 296 788 304 796
rect 316 788 324 796
rect 338 788 356 796
rect 368 788 376 796
rect 398 788 406 796
rect 428 788 436 796
rect 458 788 466 796
rect 488 788 496 796
rect 518 788 526 796
rect 548 788 556 796
rect 578 788 586 796
rect 4 778 12 786
rect 24 778 32 786
rect 54 778 62 786
rect 84 778 92 786
rect 114 778 122 786
rect 144 778 152 786
rect 174 778 182 786
rect 204 778 212 786
rect 234 778 242 786
rect 264 778 272 786
rect 286 778 294 786
rect 14 768 22 776
rect 44 768 52 776
rect 74 768 82 776
rect 4 758 12 766
rect 24 758 32 766
rect 54 758 62 766
rect 84 758 92 766
rect 114 758 122 766
rect 144 758 152 766
rect 174 758 182 766
rect 204 758 212 766
rect 234 758 242 766
rect 264 758 272 766
rect 286 758 294 766
rect 306 778 314 786
rect 328 778 336 786
rect 358 778 366 786
rect 388 778 396 786
rect 418 778 426 786
rect 448 778 456 786
rect 478 778 486 786
rect 508 778 516 786
rect 538 778 546 786
rect 568 778 576 786
rect 588 778 596 786
rect 518 768 526 776
rect 548 768 556 776
rect 578 768 586 776
rect 306 758 314 766
rect 328 758 336 766
rect 358 758 366 766
rect 388 758 396 766
rect 418 758 426 766
rect 448 758 456 766
rect 478 758 486 766
rect 508 758 516 766
rect 538 758 546 766
rect 568 758 576 766
rect 588 758 596 766
rect 14 748 22 756
rect 44 748 52 756
rect 74 748 82 756
rect 104 748 112 756
rect 134 748 142 756
rect 164 748 172 756
rect 194 748 202 756
rect 224 748 232 756
rect 244 748 262 756
rect 274 748 282 756
rect 296 748 304 756
rect 318 748 326 756
rect 338 748 356 756
rect 368 748 376 756
rect 398 748 406 756
rect 428 748 436 756
rect 458 748 466 756
rect 488 748 496 756
rect 518 748 526 756
rect 548 748 556 756
rect 578 748 586 756
rect 4 738 12 746
rect 24 738 32 746
rect 54 738 62 746
rect 84 738 92 746
rect 114 738 122 746
rect 144 738 152 746
rect 174 738 182 746
rect 204 738 212 746
rect 234 738 242 746
rect 264 738 272 746
rect 286 738 294 746
rect 306 738 314 746
rect 328 738 336 746
rect 358 738 366 746
rect 388 738 396 746
rect 418 738 426 746
rect 448 738 456 746
rect 478 738 486 746
rect 508 738 516 746
rect 538 738 546 746
rect 568 738 576 746
rect 588 738 596 746
rect 14 728 22 736
rect 224 728 232 736
rect 244 728 262 736
rect 276 728 284 736
rect 296 728 304 736
rect 316 728 324 736
rect 338 728 356 736
rect 368 728 376 736
rect 578 728 586 736
rect 4 718 12 726
rect 24 718 32 726
rect 54 718 62 726
rect 84 718 92 726
rect 114 718 122 726
rect 144 718 152 726
rect 174 718 182 726
rect 204 718 212 726
rect 234 718 242 726
rect 264 718 272 726
rect 286 718 294 726
rect 306 718 314 726
rect 328 718 336 726
rect 358 718 366 726
rect 388 718 396 726
rect 418 718 426 726
rect 448 718 456 726
rect 478 718 486 726
rect 508 718 516 726
rect 538 718 546 726
rect 568 718 576 726
rect 588 718 596 726
rect 14 708 22 716
rect 44 708 52 716
rect 74 708 82 716
rect 104 708 112 716
rect 134 708 142 716
rect 164 708 172 716
rect 194 708 202 716
rect 224 708 232 716
rect 244 708 262 716
rect 276 708 284 716
rect 296 708 304 716
rect 316 708 324 716
rect 338 708 356 716
rect 368 708 376 716
rect 398 708 406 716
rect 428 708 436 716
rect 458 708 466 716
rect 488 708 496 716
rect 518 708 526 716
rect 548 708 556 716
rect 578 708 586 716
rect 4 698 12 706
rect 24 698 32 706
rect 54 698 62 706
rect 84 698 92 706
rect 114 698 122 706
rect 144 698 152 706
rect 174 698 182 706
rect 204 698 212 706
rect 234 698 242 706
rect 264 698 272 706
rect 286 698 294 706
rect 306 698 314 706
rect 328 698 336 706
rect 358 698 366 706
rect 388 698 396 706
rect 418 698 426 706
rect 448 698 456 706
rect 478 698 486 706
rect 508 698 516 706
rect 538 698 546 706
rect 568 698 576 706
rect 588 698 596 706
rect 14 688 22 696
rect 44 688 52 696
rect 74 688 82 696
rect 104 688 112 696
rect 134 688 142 696
rect 164 688 172 696
rect 194 688 202 696
rect 224 688 232 696
rect 244 688 262 696
rect 274 688 282 696
rect 296 689 304 697
rect 318 688 326 696
rect 338 688 356 696
rect 368 688 376 696
rect 398 688 406 696
rect 428 688 436 696
rect 458 688 466 696
rect 488 688 496 696
rect 518 688 526 696
rect 548 688 556 696
rect 578 688 586 696
rect 14 644 22 652
rect 44 644 52 652
rect 74 644 82 652
rect 104 644 112 652
rect 134 644 142 652
rect 164 644 172 652
rect 4 634 12 642
rect 24 634 32 642
rect 54 634 62 642
rect 84 634 92 642
rect 114 634 122 642
rect 144 634 152 642
rect 174 634 182 642
rect 14 624 22 632
rect 44 624 52 632
rect 74 624 82 632
rect 104 624 112 632
rect 134 624 142 632
rect 164 624 172 632
rect 4 614 12 622
rect 24 614 32 622
rect 54 614 62 622
rect 84 614 92 622
rect 114 614 122 622
rect 144 614 152 622
rect 174 614 182 622
rect 14 604 22 612
rect 4 594 12 602
rect 24 594 32 602
rect 54 594 62 602
rect 84 594 92 602
rect 114 594 122 602
rect 144 594 152 602
rect 174 594 182 602
rect 14 584 22 592
rect 44 584 52 592
rect 74 584 82 592
rect 104 584 112 592
rect 134 584 142 592
rect 164 584 172 592
rect 4 574 12 582
rect 24 574 32 582
rect 54 574 62 582
rect 84 574 92 582
rect 14 564 22 572
rect 44 564 52 572
rect 74 564 82 572
rect 104 564 112 572
rect 134 564 142 572
rect 164 564 172 572
rect 4 554 12 562
rect 24 554 32 562
rect 54 554 62 562
rect 84 554 92 562
rect 114 554 122 562
rect 144 554 152 562
rect 174 554 182 562
rect 14 544 22 552
rect 44 544 52 552
rect 74 544 82 552
rect 104 544 112 552
rect 134 544 142 552
rect 164 544 172 552
rect 4 534 12 542
rect 24 534 32 542
rect 54 534 62 542
rect 84 534 92 542
rect 114 534 122 542
rect 144 534 152 542
rect 174 534 182 542
rect 14 524 22 532
rect 44 524 52 532
rect 74 524 82 532
rect 104 524 112 532
rect 134 524 142 532
rect 164 524 172 532
rect 14 508 22 516
rect 34 508 42 516
rect 54 508 62 516
rect 74 508 82 516
rect 94 508 102 516
rect 114 508 122 516
rect 134 508 142 516
rect 154 508 162 516
rect 174 508 182 516
rect 290 644 298 652
rect 302 644 310 652
rect 290 624 298 632
rect 302 624 310 632
rect 290 604 298 612
rect 302 604 310 612
rect 290 586 298 594
rect 302 586 310 594
rect 290 556 298 564
rect 302 556 310 564
rect 290 536 298 544
rect 302 536 310 544
rect 290 516 298 524
rect 302 516 310 524
rect 428 644 436 652
rect 458 644 466 652
rect 488 644 496 652
rect 518 644 526 652
rect 548 644 556 652
rect 578 644 586 652
rect 418 634 426 642
rect 448 634 456 642
rect 478 634 486 642
rect 508 634 516 642
rect 538 634 546 642
rect 568 634 576 642
rect 588 634 596 642
rect 428 624 436 632
rect 458 624 466 632
rect 488 624 496 632
rect 518 624 526 632
rect 548 624 556 632
rect 578 624 586 632
rect 418 614 426 622
rect 448 614 456 622
rect 478 614 486 622
rect 508 614 516 622
rect 538 614 546 622
rect 568 614 576 622
rect 588 614 596 622
rect 578 604 586 612
rect 418 594 426 602
rect 448 594 456 602
rect 478 594 486 602
rect 508 594 516 602
rect 538 594 546 602
rect 568 594 576 602
rect 588 594 596 602
rect 428 584 436 592
rect 458 584 466 592
rect 488 584 496 592
rect 518 584 526 592
rect 548 584 556 592
rect 578 584 586 592
rect 508 574 516 582
rect 538 574 546 582
rect 568 574 576 582
rect 588 574 596 582
rect 428 564 436 572
rect 458 564 466 572
rect 488 564 496 572
rect 518 564 526 572
rect 548 564 556 572
rect 578 564 586 572
rect 418 554 426 562
rect 448 554 456 562
rect 478 554 486 562
rect 508 554 516 562
rect 538 554 546 562
rect 568 554 576 562
rect 588 554 596 562
rect 428 544 436 552
rect 458 544 466 552
rect 488 544 496 552
rect 518 544 526 552
rect 548 544 556 552
rect 578 544 586 552
rect 418 534 426 542
rect 448 534 456 542
rect 478 534 486 542
rect 508 534 516 542
rect 538 534 546 542
rect 568 534 576 542
rect 588 534 596 542
rect 428 524 436 532
rect 458 524 466 532
rect 488 524 496 532
rect 518 524 526 532
rect 548 524 556 532
rect 578 524 586 532
rect 418 508 426 516
rect 438 508 446 516
rect 458 508 466 516
rect 478 508 486 516
rect 498 508 506 516
rect 518 508 526 516
rect 538 508 546 516
rect 558 508 566 516
rect 578 508 586 516
rect 30 451 38 459
rect 50 451 58 459
rect 80 451 88 459
rect 110 451 118 459
rect 140 451 148 459
rect 170 451 178 459
rect 200 451 208 459
rect 230 451 238 459
rect 260 451 268 459
rect 290 451 298 459
rect 320 451 328 459
rect 350 451 358 459
rect 380 451 388 459
rect 410 451 418 459
rect 440 451 448 459
rect 470 451 478 459
rect 500 451 508 459
rect 530 451 538 459
rect 560 451 568 459
rect 40 441 48 449
rect 70 441 78 449
rect 100 441 108 449
rect 130 441 138 449
rect 160 441 168 449
rect 190 441 198 449
rect 220 441 228 449
rect 250 441 258 449
rect 280 441 288 449
rect 310 441 318 449
rect 340 441 348 449
rect 370 441 378 449
rect 400 441 408 449
rect 430 441 438 449
rect 460 441 468 449
rect 490 441 498 449
rect 520 441 528 449
rect 550 441 558 449
rect 30 431 38 439
rect 50 431 58 439
rect 80 431 88 439
rect 110 431 118 439
rect 140 431 148 439
rect 170 431 178 439
rect 200 431 208 439
rect 230 431 238 439
rect 260 431 268 439
rect 290 431 298 439
rect 320 431 328 439
rect 350 431 358 439
rect 380 431 388 439
rect 410 431 418 439
rect 440 431 448 439
rect 470 431 478 439
rect 500 431 508 439
rect 530 431 538 439
rect 560 431 568 439
rect 40 421 48 429
rect 70 421 78 429
rect 100 421 108 429
rect 130 421 138 429
rect 160 421 168 429
rect 190 421 198 429
rect 220 421 228 429
rect 250 421 258 429
rect 280 421 288 429
rect 310 421 318 429
rect 340 421 348 429
rect 370 421 378 429
rect 400 421 408 429
rect 430 421 438 429
rect 460 421 468 429
rect 490 421 498 429
rect 520 421 528 429
rect 550 421 558 429
rect 30 411 38 419
rect 50 411 58 419
rect 80 411 88 419
rect 110 411 118 419
rect 140 411 148 419
rect 170 411 178 419
rect 200 411 208 419
rect 230 411 238 419
rect 260 411 268 419
rect 290 411 298 419
rect 320 411 328 419
rect 350 411 358 419
rect 380 411 388 419
rect 410 411 418 419
rect 440 411 448 419
rect 470 411 478 419
rect 500 411 508 419
rect 530 411 538 419
rect 560 411 568 419
rect 40 401 48 409
rect 70 401 78 409
rect 100 401 108 409
rect 130 401 138 409
rect 160 401 168 409
rect 190 401 198 409
rect 220 401 228 409
rect 250 401 258 409
rect 280 401 288 409
rect 310 401 318 409
rect 340 401 348 409
rect 370 401 378 409
rect 400 401 408 409
rect 430 401 438 409
rect 460 401 468 409
rect 490 401 498 409
rect 520 401 528 409
rect 550 401 558 409
rect 30 371 38 399
rect 50 371 58 399
rect 80 371 88 399
rect 110 391 118 399
rect 140 391 148 399
rect 170 391 178 399
rect 200 391 208 399
rect 230 391 238 399
rect 260 391 268 399
rect 290 391 298 399
rect 320 391 328 399
rect 350 391 358 399
rect 380 391 388 399
rect 410 391 418 399
rect 440 391 448 399
rect 470 391 478 399
rect 110 371 118 379
rect 140 371 148 379
rect 170 371 178 379
rect 200 371 208 379
rect 230 371 238 379
rect 260 371 268 379
rect 290 371 298 379
rect 320 371 328 379
rect 350 371 358 379
rect 380 371 388 379
rect 410 371 418 379
rect 440 371 448 379
rect 470 371 478 379
rect 500 371 508 399
rect 530 391 538 399
rect 560 391 568 399
rect 520 381 528 389
rect 550 381 558 389
rect 530 371 538 379
rect 560 371 568 379
rect 40 361 48 369
rect 70 361 78 369
rect 100 361 108 369
rect 130 361 138 369
rect 160 361 168 369
rect 190 361 198 369
rect 220 361 228 369
rect 250 361 258 369
rect 280 361 288 369
rect 310 361 318 369
rect 340 361 348 369
rect 370 361 378 369
rect 400 361 408 369
rect 430 361 438 369
rect 460 361 468 369
rect 490 361 498 369
rect 520 361 528 369
rect 550 361 558 369
rect 30 351 38 359
rect 50 351 58 359
rect 80 351 88 359
rect 110 351 118 359
rect 140 351 148 359
rect 170 351 178 359
rect 200 351 208 359
rect 230 351 238 359
rect 260 351 268 359
rect 290 351 298 359
rect 320 351 328 359
rect 350 351 358 359
rect 380 351 388 359
rect 410 351 418 359
rect 440 351 448 359
rect 470 351 478 359
rect 500 351 508 359
rect 530 351 538 359
rect 560 351 568 359
rect 40 341 48 349
rect 70 341 78 349
rect 100 341 108 349
rect 130 341 138 349
rect 160 341 168 349
rect 190 341 198 349
rect 220 341 228 349
rect 250 341 258 349
rect 280 341 288 349
rect 310 341 318 349
rect 340 341 348 349
rect 370 341 378 349
rect 400 341 408 349
rect 430 341 438 349
rect 460 341 468 349
rect 490 341 498 349
rect 520 341 528 349
rect 550 341 558 349
rect 30 331 38 339
rect 50 331 58 339
rect 80 331 88 339
rect 110 331 118 339
rect 140 331 148 339
rect 170 331 178 339
rect 200 331 208 339
rect 230 331 238 339
rect 260 331 268 339
rect 290 331 298 339
rect 320 331 328 339
rect 350 331 358 339
rect 380 331 388 339
rect 410 331 418 339
rect 440 331 448 339
rect 470 331 478 339
rect 500 331 508 339
rect 530 331 538 339
rect 560 331 568 339
rect 40 321 48 329
rect 70 321 78 329
rect 100 321 108 329
rect 130 321 138 329
rect 160 321 168 329
rect 190 321 198 329
rect 220 321 228 329
rect 250 321 258 329
rect 280 321 288 329
rect 310 321 318 329
rect 340 321 348 329
rect 370 321 378 329
rect 400 321 408 329
rect 430 321 438 329
rect 460 321 468 329
rect 490 321 498 329
rect 520 321 528 329
rect 550 321 558 329
rect 30 311 38 319
rect 50 311 58 319
rect 80 311 88 319
rect 110 311 118 319
rect 140 311 148 319
rect 170 311 178 319
rect 200 311 208 319
rect 230 311 238 319
rect 260 311 268 319
rect 290 311 298 319
rect 320 311 328 319
rect 350 311 358 319
rect 380 311 388 319
rect 410 311 418 319
rect 440 311 448 319
rect 470 311 478 319
rect 500 311 508 319
rect 530 311 538 319
rect 560 311 568 319
rect 40 301 48 309
rect 70 301 78 309
rect 90 301 98 309
rect 520 301 528 309
rect 550 301 558 309
rect 30 291 38 299
rect 50 291 58 299
rect 80 291 88 299
rect 110 291 118 299
rect 140 291 148 299
rect 170 291 178 299
rect 200 291 208 299
rect 230 291 238 299
rect 260 291 268 299
rect 290 291 298 299
rect 320 291 328 299
rect 350 291 358 299
rect 380 291 388 299
rect 410 291 418 299
rect 440 291 448 299
rect 470 291 478 299
rect 500 291 508 299
rect 530 291 538 299
rect 560 291 568 299
rect 40 281 48 289
rect 70 281 78 289
rect 100 281 108 289
rect 130 281 138 289
rect 160 281 168 289
rect 190 281 198 289
rect 220 281 228 289
rect 250 281 258 289
rect 280 281 288 289
rect 310 281 318 289
rect 340 281 348 289
rect 370 281 378 289
rect 400 281 408 289
rect 430 281 438 289
rect 460 281 468 289
rect 490 281 498 289
rect 520 281 528 289
rect 550 281 558 289
rect 30 271 38 279
rect 50 271 58 279
rect 80 271 88 279
rect 110 271 118 279
rect 140 271 148 279
rect 170 271 178 279
rect 200 271 208 279
rect 230 271 238 279
rect 260 271 268 279
rect 290 271 298 279
rect 320 271 328 279
rect 350 271 358 279
rect 380 271 388 279
rect 410 271 418 279
rect 440 271 448 279
rect 470 271 478 279
rect 500 271 508 279
rect 530 271 538 279
rect 560 271 568 279
rect 40 261 48 269
rect 70 261 78 269
rect 100 261 108 269
rect 130 261 138 269
rect 160 261 168 269
rect 190 261 198 269
rect 220 261 228 269
rect 250 261 258 269
rect 280 261 288 269
rect 310 261 318 269
rect 340 261 348 269
rect 370 261 378 269
rect 400 261 408 269
rect 430 261 438 269
rect 460 261 468 269
rect 490 261 498 269
rect 520 261 528 269
rect 550 261 558 269
rect 30 251 38 259
rect 50 251 58 259
rect 80 251 88 259
rect 110 251 118 259
rect 140 251 148 259
rect 170 251 178 259
rect 200 251 208 259
rect 230 251 238 259
rect 260 251 268 259
rect 290 251 298 259
rect 320 251 328 259
rect 350 251 358 259
rect 380 251 388 259
rect 410 251 418 259
rect 440 251 448 259
rect 470 251 478 259
rect 500 251 508 259
rect 530 251 538 259
rect 560 251 568 259
rect 40 241 48 249
rect 30 231 38 239
rect 50 231 58 239
rect 40 221 48 229
rect 70 221 78 249
rect 100 241 108 249
rect 130 241 138 249
rect 160 241 168 249
rect 190 241 198 249
rect 220 241 228 249
rect 250 241 258 249
rect 280 241 288 249
rect 310 241 318 249
rect 340 241 348 249
rect 370 241 378 249
rect 400 241 408 249
rect 430 241 438 249
rect 460 241 468 249
rect 490 241 498 249
rect 520 241 528 249
rect 550 241 558 249
rect 510 231 518 239
rect 530 231 538 239
rect 560 231 568 239
rect 100 221 108 229
rect 130 221 138 229
rect 160 221 168 229
rect 190 221 198 229
rect 220 221 228 229
rect 250 221 258 229
rect 280 221 288 229
rect 310 221 318 229
rect 340 221 348 229
rect 370 221 378 229
rect 400 221 408 229
rect 430 221 438 229
rect 460 221 468 229
rect 490 221 498 229
rect 520 221 528 229
rect 550 221 558 229
rect 30 211 38 219
rect 50 211 58 219
rect 80 211 88 219
rect 110 211 118 219
rect 140 211 148 219
rect 170 211 178 219
rect 200 211 208 219
rect 230 211 238 219
rect 260 211 268 219
rect 290 211 298 219
rect 320 211 328 219
rect 350 211 358 219
rect 380 211 388 219
rect 410 211 418 219
rect 440 211 448 219
rect 470 211 478 219
rect 500 211 508 219
rect 530 211 538 219
rect 560 211 568 219
rect 40 201 48 209
rect 70 201 78 209
rect 100 201 108 209
rect 130 201 138 209
rect 160 201 168 209
rect 190 201 198 209
rect 220 201 228 209
rect 250 201 258 209
rect 280 201 288 209
rect 310 201 318 209
rect 340 201 348 209
rect 370 201 378 209
rect 400 201 408 209
rect 430 201 438 209
rect 460 201 468 209
rect 490 201 498 209
rect 520 201 528 209
rect 550 201 558 209
rect 30 191 38 199
rect 50 191 58 199
rect 80 191 88 199
rect 110 191 118 199
rect 140 191 148 199
rect 170 191 178 199
rect 200 191 208 199
rect 230 191 238 199
rect 260 191 268 199
rect 290 191 298 199
rect 320 191 328 199
rect 350 191 358 199
rect 380 191 388 199
rect 410 191 418 199
rect 440 191 448 199
rect 470 191 478 199
rect 500 191 508 199
rect 530 191 538 199
rect 560 191 568 199
rect 40 181 48 189
rect 70 181 78 189
rect 100 181 108 189
rect 130 181 138 189
rect 160 181 168 189
rect 190 181 198 189
rect 220 181 228 189
rect 250 181 258 189
rect 280 181 288 189
rect 310 181 318 189
rect 340 181 348 189
rect 370 181 378 189
rect 400 181 408 189
rect 430 181 438 189
rect 460 181 468 189
rect 490 181 498 189
rect 520 181 528 189
rect 550 181 558 189
rect 30 171 38 179
rect 50 171 58 179
rect 80 171 88 179
rect 110 171 118 179
rect 140 171 148 179
rect 170 171 178 179
rect 200 171 208 179
rect 230 171 238 179
rect 260 171 268 179
rect 290 171 298 179
rect 320 171 328 179
rect 350 171 358 179
rect 380 171 388 179
rect 410 171 418 179
rect 440 171 448 179
rect 470 171 478 179
rect 500 171 508 179
rect 530 171 538 179
rect 560 171 568 179
rect 40 161 48 169
rect 70 161 78 169
rect 100 161 108 169
rect 130 161 138 169
rect 160 161 168 169
rect 190 161 198 169
rect 220 161 228 169
rect 250 161 258 169
rect 280 161 288 169
rect 310 161 318 169
rect 340 161 348 169
rect 370 161 378 169
rect 400 161 408 169
rect 430 161 438 169
rect 460 161 468 169
rect 490 161 498 169
rect 520 161 528 169
rect 550 161 558 169
rect 30 151 38 159
rect 50 151 58 159
rect 80 151 88 159
rect 510 151 518 159
rect 530 151 538 159
rect 560 151 568 159
rect 40 141 48 149
rect 70 141 78 149
rect 100 141 108 149
rect 130 141 138 149
rect 160 141 168 149
rect 190 141 198 149
rect 220 141 228 149
rect 250 141 258 149
rect 280 141 288 149
rect 310 141 318 149
rect 340 141 348 149
rect 370 141 378 149
rect 400 141 408 149
rect 430 141 438 149
rect 460 141 468 149
rect 490 141 498 149
rect 520 141 528 149
rect 550 141 558 149
rect 30 131 38 139
rect 50 131 58 139
rect 80 131 88 139
rect 110 131 118 139
rect 140 131 148 139
rect 170 131 178 139
rect 200 131 208 139
rect 230 131 238 139
rect 260 131 268 139
rect 290 131 298 139
rect 320 131 328 139
rect 350 131 358 139
rect 380 131 388 139
rect 410 131 418 139
rect 440 131 448 139
rect 470 131 478 139
rect 500 131 508 139
rect 530 131 538 139
rect 560 131 568 139
rect 40 121 48 129
rect 70 121 78 129
rect 100 121 108 129
rect 130 121 138 129
rect 160 121 168 129
rect 190 121 198 129
rect 220 121 228 129
rect 250 121 258 129
rect 280 121 288 129
rect 310 121 318 129
rect 340 121 348 129
rect 370 121 378 129
rect 400 121 408 129
rect 430 121 438 129
rect 460 121 468 129
rect 490 121 498 129
rect 520 121 528 129
rect 550 121 558 129
rect 30 111 38 119
rect 50 111 58 119
rect 80 111 88 119
rect 110 111 118 119
rect 140 111 148 119
rect 170 111 178 119
rect 200 111 208 119
rect 230 111 238 119
rect 260 111 268 119
rect 290 111 298 119
rect 320 111 328 119
rect 350 111 358 119
rect 380 111 388 119
rect 410 111 418 119
rect 440 111 448 119
rect 470 111 478 119
rect 500 111 508 119
rect 530 111 538 119
rect 560 111 568 119
rect 40 101 48 109
rect 70 101 78 109
rect 100 101 108 109
rect 130 101 138 109
rect 160 101 168 109
rect 190 101 198 109
rect 220 101 228 109
rect 250 101 258 109
rect 280 101 288 109
rect 310 101 318 109
rect 340 101 348 109
rect 370 101 378 109
rect 400 101 408 109
rect 430 101 438 109
rect 460 101 468 109
rect 490 101 498 109
rect 520 101 528 109
rect 550 101 558 109
rect 30 91 38 99
rect 50 91 58 99
rect 80 91 88 99
rect 110 91 118 99
rect 140 91 148 99
rect 170 91 178 99
rect 200 91 208 99
rect 230 91 238 99
rect 260 91 268 99
rect 290 91 298 99
rect 320 91 328 99
rect 350 91 358 99
rect 380 91 388 99
rect 410 91 418 99
rect 440 91 448 99
rect 470 91 478 99
rect 500 91 508 99
rect 530 91 538 99
rect 560 91 568 99
rect 40 81 48 89
rect 70 81 78 89
rect 100 81 108 89
rect 130 81 138 89
rect 160 81 168 89
rect 190 81 198 89
rect 220 81 228 89
rect 250 81 258 89
rect 280 81 288 89
rect 310 81 318 89
rect 340 81 348 89
rect 370 81 378 89
rect 400 81 408 89
rect 430 81 438 89
rect 460 81 468 89
rect 490 81 498 89
rect 520 81 528 89
rect 550 81 558 89
rect 30 71 38 79
rect 50 71 58 79
rect 80 71 88 79
rect 110 71 118 79
rect 140 71 148 79
rect 170 71 178 79
rect 200 71 208 79
rect 230 71 238 79
rect 260 71 268 79
rect 290 71 298 79
rect 320 71 328 79
rect 350 71 358 79
rect 380 71 388 79
rect 410 71 418 79
rect 440 71 448 79
rect 470 71 478 79
rect 500 71 508 79
rect 530 71 538 79
rect 560 71 568 79
rect 40 61 48 69
rect 70 61 78 69
rect 100 61 108 69
rect 130 61 138 69
rect 160 61 168 69
rect 190 61 198 69
rect 220 61 228 69
rect 250 61 258 69
rect 280 61 288 69
rect 310 61 318 69
rect 340 61 348 69
rect 370 61 378 69
rect 400 61 408 69
rect 430 61 438 69
rect 460 61 468 69
rect 490 61 498 69
rect 520 61 528 69
rect 550 61 558 69
rect 30 51 38 59
rect 50 51 58 59
rect 80 51 88 59
rect 110 51 118 59
rect 140 51 148 59
rect 170 51 178 59
rect 200 51 208 59
rect 230 51 238 59
rect 260 51 268 59
rect 290 51 298 59
rect 320 51 328 59
rect 350 51 358 59
rect 380 51 388 59
rect 410 51 418 59
rect 440 51 448 59
rect 470 51 478 59
rect 500 51 508 59
rect 530 51 538 59
rect 560 51 568 59
rect 40 41 48 49
rect 70 41 78 49
rect 100 41 108 49
rect 130 41 138 49
rect 160 41 168 49
rect 190 41 198 49
rect 220 41 228 49
rect 250 41 258 49
rect 280 41 288 49
rect 310 41 318 49
rect 340 41 348 49
rect 370 41 378 49
rect 400 41 408 49
rect 430 41 438 49
rect 460 41 468 49
rect 490 41 498 49
rect 520 41 528 49
rect 550 41 558 49
rect 30 31 38 39
rect 50 31 58 39
rect 80 31 88 39
rect 110 31 118 39
rect 140 31 148 39
rect 170 31 178 39
rect 200 31 208 39
rect 230 31 238 39
rect 260 31 268 39
rect 290 31 298 39
rect 320 31 328 39
rect 350 31 358 39
rect 380 31 388 39
rect 410 31 418 39
rect 440 31 448 39
rect 470 31 478 39
rect 500 31 508 39
rect 530 31 538 39
rect 560 31 568 39
rect 206 4 394 12
<< metal2 >>
rect 0 1298 600 1340
rect 0 1290 42 1298
rect 50 1290 62 1298
rect 70 1294 530 1298
rect 70 1290 92 1294
rect 0 1287 72 1290
rect 0 1279 50 1287
rect 58 1282 72 1287
rect 80 1286 92 1290
rect 100 1286 112 1294
rect 120 1286 132 1294
rect 140 1286 152 1294
rect 160 1286 172 1294
rect 180 1286 192 1294
rect 200 1286 212 1294
rect 220 1286 232 1294
rect 240 1286 360 1294
rect 368 1286 380 1294
rect 388 1286 400 1294
rect 408 1286 420 1294
rect 428 1286 440 1294
rect 448 1286 460 1294
rect 468 1286 480 1294
rect 488 1286 500 1294
rect 508 1290 530 1294
rect 538 1290 550 1298
rect 558 1290 600 1298
rect 508 1286 520 1290
rect 80 1284 520 1286
rect 528 1287 600 1290
rect 58 1279 82 1282
rect 0 1278 82 1279
rect 0 1270 42 1278
rect 50 1276 82 1278
rect 90 1276 102 1284
rect 110 1276 122 1284
rect 130 1276 142 1284
rect 150 1276 162 1284
rect 170 1276 182 1284
rect 190 1276 202 1284
rect 210 1276 222 1284
rect 230 1276 370 1284
rect 378 1276 390 1284
rect 398 1276 410 1284
rect 418 1276 430 1284
rect 438 1276 450 1284
rect 458 1276 470 1284
rect 478 1276 490 1284
rect 498 1276 510 1284
rect 528 1282 542 1287
rect 518 1279 542 1282
rect 550 1279 600 1287
rect 518 1278 600 1279
rect 518 1276 550 1278
rect 50 1270 550 1276
rect 558 1270 600 1278
rect 0 1267 600 1270
rect 0 1259 50 1267
rect 58 1259 542 1267
rect 550 1259 600 1267
rect 0 1258 600 1259
rect 0 1250 42 1258
rect 50 1250 550 1258
rect 558 1250 600 1258
rect 0 1247 78 1250
rect 0 1239 50 1247
rect 58 1239 78 1247
rect 236 1242 364 1250
rect 522 1247 600 1250
rect 0 1238 78 1239
rect 0 1230 42 1238
rect 50 1230 78 1238
rect 0 1227 78 1230
rect 0 1219 50 1227
rect 58 1219 78 1227
rect 0 1218 78 1219
rect 0 1210 42 1218
rect 50 1210 78 1218
rect 0 1207 78 1210
rect 0 1199 50 1207
rect 58 1199 78 1207
rect 0 1198 78 1199
rect 0 1190 42 1198
rect 50 1190 78 1198
rect 0 1187 78 1190
rect 0 1179 50 1187
rect 58 1179 78 1187
rect 96 1220 504 1242
rect 96 1212 290 1220
rect 298 1212 302 1220
rect 310 1212 504 1220
rect 96 1200 504 1212
rect 96 1192 290 1200
rect 298 1192 302 1200
rect 310 1192 504 1200
rect 96 1190 504 1192
rect 96 1180 100 1190
rect 500 1180 504 1190
rect 522 1239 542 1247
rect 550 1239 600 1247
rect 522 1238 600 1239
rect 522 1230 550 1238
rect 558 1230 600 1238
rect 522 1227 600 1230
rect 522 1219 542 1227
rect 550 1219 600 1227
rect 522 1218 600 1219
rect 522 1210 550 1218
rect 558 1210 600 1218
rect 522 1207 600 1210
rect 522 1199 542 1207
rect 550 1199 600 1207
rect 522 1198 600 1199
rect 522 1190 550 1198
rect 558 1190 600 1198
rect 522 1187 600 1190
rect 0 1178 78 1179
rect 0 1170 42 1178
rect 50 1172 78 1178
rect 236 1172 364 1180
rect 522 1179 542 1187
rect 550 1179 600 1187
rect 522 1178 600 1179
rect 522 1172 550 1178
rect 50 1170 550 1172
rect 558 1170 600 1178
rect 0 1167 600 1170
rect 0 1159 50 1167
rect 58 1159 542 1167
rect 550 1159 600 1167
rect 0 1158 600 1159
rect 0 1150 42 1158
rect 50 1150 550 1158
rect 558 1150 600 1158
rect 0 1147 600 1150
rect 0 1139 50 1147
rect 58 1139 542 1147
rect 550 1139 600 1147
rect 0 1138 600 1139
rect 0 1130 42 1138
rect 50 1130 550 1138
rect 558 1130 600 1138
rect 0 1127 600 1130
rect 0 1119 50 1127
rect 58 1122 542 1127
rect 58 1119 78 1122
rect 0 1118 78 1119
rect 0 1110 42 1118
rect 50 1110 78 1118
rect 236 1114 364 1122
rect 522 1119 542 1122
rect 550 1119 600 1127
rect 522 1118 600 1119
rect 0 1107 78 1110
rect 0 1099 50 1107
rect 58 1099 78 1107
rect 0 1098 78 1099
rect 0 1090 42 1098
rect 50 1090 78 1098
rect 0 1087 78 1090
rect 0 1079 50 1087
rect 58 1079 78 1087
rect 0 1078 78 1079
rect 0 1070 42 1078
rect 50 1070 78 1078
rect 0 1067 78 1070
rect 0 1059 50 1067
rect 58 1059 78 1067
rect 0 1058 78 1059
rect 0 1050 42 1058
rect 50 1050 78 1058
rect 96 1092 504 1114
rect 96 1084 290 1092
rect 298 1084 302 1092
rect 310 1084 504 1092
rect 96 1072 504 1084
rect 96 1064 290 1072
rect 298 1064 302 1072
rect 310 1064 504 1072
rect 96 1052 504 1064
rect 522 1110 550 1118
rect 558 1110 600 1118
rect 522 1107 600 1110
rect 522 1099 542 1107
rect 550 1099 600 1107
rect 522 1098 600 1099
rect 522 1090 550 1098
rect 558 1090 600 1098
rect 522 1087 600 1090
rect 522 1079 542 1087
rect 550 1079 600 1087
rect 522 1078 600 1079
rect 522 1070 550 1078
rect 558 1070 600 1078
rect 522 1067 600 1070
rect 522 1059 542 1067
rect 550 1059 600 1067
rect 522 1058 600 1059
rect 0 1047 78 1050
rect 0 1039 50 1047
rect 58 1044 78 1047
rect 236 1044 364 1052
rect 522 1050 550 1058
rect 558 1050 600 1058
rect 522 1047 600 1050
rect 522 1044 542 1047
rect 58 1040 542 1044
rect 58 1039 100 1040
rect 0 1038 100 1039
rect 0 1030 42 1038
rect 50 1030 100 1038
rect 500 1039 542 1040
rect 550 1039 600 1047
rect 500 1038 600 1039
rect 500 1030 550 1038
rect 558 1030 600 1038
rect 0 1027 600 1030
rect 0 1019 50 1027
rect 58 1019 542 1027
rect 550 1019 600 1027
rect 0 1018 600 1019
rect 0 1010 42 1018
rect 50 1010 550 1018
rect 558 1010 600 1018
rect 0 1007 600 1010
rect 0 999 50 1007
rect 58 999 542 1007
rect 550 999 600 1007
rect 0 998 600 999
rect 0 990 42 998
rect 50 992 550 998
rect 50 990 78 992
rect 0 987 78 990
rect 0 979 50 987
rect 58 979 78 987
rect 236 984 364 992
rect 522 990 550 992
rect 558 990 600 998
rect 522 987 600 990
rect 0 978 78 979
rect 0 970 42 978
rect 50 970 78 978
rect 0 967 78 970
rect 0 959 50 967
rect 58 959 78 967
rect 0 958 78 959
rect 0 950 42 958
rect 50 950 78 958
rect 0 947 78 950
rect 0 939 50 947
rect 58 939 78 947
rect 0 938 78 939
rect 0 930 42 938
rect 50 930 78 938
rect 0 927 78 930
rect 0 919 50 927
rect 58 919 78 927
rect 96 962 504 984
rect 96 954 290 962
rect 298 954 302 962
rect 310 954 504 962
rect 96 942 504 954
rect 96 934 290 942
rect 298 934 302 942
rect 310 934 504 942
rect 96 922 504 934
rect 522 979 542 987
rect 550 979 600 987
rect 522 978 600 979
rect 522 970 550 978
rect 558 970 600 978
rect 522 967 600 970
rect 522 959 542 967
rect 550 959 600 967
rect 522 958 600 959
rect 522 950 550 958
rect 558 950 600 958
rect 522 947 600 950
rect 522 939 542 947
rect 550 939 600 947
rect 522 938 600 939
rect 522 930 550 938
rect 558 930 600 938
rect 522 927 600 930
rect 0 918 78 919
rect 0 910 42 918
rect 50 914 78 918
rect 236 914 364 922
rect 522 919 542 927
rect 550 919 600 927
rect 522 918 600 919
rect 522 914 550 918
rect 50 910 550 914
rect 558 910 600 918
rect 0 907 600 910
rect 0 899 50 907
rect 58 899 542 907
rect 550 899 600 907
rect 0 898 600 899
rect 0 890 42 898
rect 50 890 550 898
rect 558 890 600 898
rect 0 888 600 890
rect 0 880 50 888
rect 58 880 542 888
rect 550 880 600 888
rect 0 844 600 848
rect 0 836 24 844
rect 42 836 54 844
rect 72 836 84 844
rect 102 836 114 844
rect 132 836 144 844
rect 162 836 174 844
rect 192 836 204 844
rect 222 836 234 844
rect 242 836 264 844
rect 272 836 286 844
rect 294 836 306 844
rect 314 836 328 844
rect 336 836 358 844
rect 366 836 378 844
rect 396 836 408 844
rect 426 836 438 844
rect 456 836 468 844
rect 486 836 498 844
rect 516 836 528 844
rect 546 836 558 844
rect 576 836 600 844
rect 0 828 14 836
rect 22 828 44 836
rect 52 828 74 836
rect 82 828 104 836
rect 112 828 134 836
rect 142 828 164 836
rect 172 828 194 836
rect 202 828 224 836
rect 232 828 244 836
rect 262 828 274 836
rect 282 828 296 836
rect 304 828 318 836
rect 326 828 338 836
rect 356 828 368 836
rect 376 828 398 836
rect 406 828 428 836
rect 436 828 458 836
rect 466 828 488 836
rect 496 828 518 836
rect 526 828 548 836
rect 556 828 578 836
rect 586 828 600 836
rect 0 826 600 828
rect 0 818 4 826
rect 12 818 24 826
rect 32 818 54 826
rect 62 818 84 826
rect 92 818 114 826
rect 122 818 144 826
rect 152 818 174 826
rect 182 818 204 826
rect 212 818 234 826
rect 242 818 264 826
rect 272 818 286 826
rect 294 818 306 826
rect 314 818 328 826
rect 336 818 358 826
rect 366 818 388 826
rect 396 818 418 826
rect 426 818 448 826
rect 456 818 478 826
rect 486 818 508 826
rect 516 818 538 826
rect 546 818 568 826
rect 576 818 588 826
rect 596 818 600 826
rect 0 816 600 818
rect 0 808 14 816
rect 22 808 44 816
rect 52 808 74 816
rect 82 808 104 816
rect 112 808 134 816
rect 142 808 164 816
rect 172 808 194 816
rect 202 808 224 816
rect 232 808 244 816
rect 262 808 276 816
rect 284 808 296 816
rect 304 808 316 816
rect 324 808 338 816
rect 356 808 368 816
rect 376 808 398 816
rect 406 808 428 816
rect 436 808 458 816
rect 466 808 488 816
rect 496 808 518 816
rect 526 808 548 816
rect 556 808 578 816
rect 586 808 600 816
rect 0 806 600 808
rect 0 798 4 806
rect 12 798 24 806
rect 32 798 54 806
rect 62 798 84 806
rect 92 798 114 806
rect 122 798 144 806
rect 152 798 174 806
rect 182 798 204 806
rect 212 798 234 806
rect 242 798 264 806
rect 272 798 286 806
rect 294 798 306 806
rect 314 798 328 806
rect 336 798 358 806
rect 366 798 388 806
rect 396 798 418 806
rect 426 798 448 806
rect 456 798 478 806
rect 486 798 508 806
rect 516 798 538 806
rect 546 798 568 806
rect 576 798 588 806
rect 596 798 600 806
rect 0 796 600 798
rect 0 788 14 796
rect 22 788 44 796
rect 52 788 74 796
rect 82 788 104 796
rect 112 788 134 796
rect 142 788 164 796
rect 172 788 194 796
rect 202 788 224 796
rect 232 788 244 796
rect 262 788 276 796
rect 284 788 296 796
rect 304 788 316 796
rect 324 788 338 796
rect 356 788 368 796
rect 376 788 398 796
rect 406 788 428 796
rect 436 788 458 796
rect 466 788 488 796
rect 496 788 518 796
rect 526 788 548 796
rect 556 788 578 796
rect 586 788 600 796
rect 0 786 600 788
rect 0 778 4 786
rect 12 778 24 786
rect 32 778 54 786
rect 62 778 84 786
rect 92 778 114 786
rect 122 778 144 786
rect 152 778 174 786
rect 182 778 204 786
rect 212 778 234 786
rect 242 778 264 786
rect 272 778 286 786
rect 294 778 306 786
rect 314 778 328 786
rect 336 778 358 786
rect 366 778 388 786
rect 396 778 418 786
rect 426 778 448 786
rect 456 778 478 786
rect 486 778 508 786
rect 516 778 538 786
rect 546 778 568 786
rect 576 778 588 786
rect 596 778 600 786
rect 0 776 100 778
rect 0 768 14 776
rect 22 768 44 776
rect 52 768 74 776
rect 82 768 100 776
rect 500 776 600 778
rect 500 768 518 776
rect 526 768 548 776
rect 556 768 578 776
rect 586 768 600 776
rect 0 766 600 768
rect 0 758 4 766
rect 12 758 24 766
rect 32 758 54 766
rect 62 758 84 766
rect 92 758 114 766
rect 122 758 144 766
rect 152 758 174 766
rect 182 758 204 766
rect 212 758 234 766
rect 242 758 264 766
rect 272 758 286 766
rect 294 758 306 766
rect 314 758 328 766
rect 336 758 358 766
rect 366 758 388 766
rect 396 758 418 766
rect 426 758 448 766
rect 456 758 478 766
rect 486 758 508 766
rect 516 758 538 766
rect 546 758 568 766
rect 576 758 588 766
rect 596 758 600 766
rect 0 756 600 758
rect 0 748 14 756
rect 22 748 44 756
rect 52 748 74 756
rect 82 748 104 756
rect 112 748 134 756
rect 142 748 164 756
rect 172 748 194 756
rect 202 748 224 756
rect 232 748 244 756
rect 262 748 274 756
rect 282 748 296 756
rect 304 748 318 756
rect 326 748 338 756
rect 356 748 368 756
rect 376 748 398 756
rect 406 748 428 756
rect 436 748 458 756
rect 466 748 488 756
rect 496 748 518 756
rect 526 748 548 756
rect 556 748 578 756
rect 586 748 600 756
rect 0 746 600 748
rect 0 738 4 746
rect 12 738 24 746
rect 32 738 54 746
rect 62 738 84 746
rect 92 738 114 746
rect 122 738 144 746
rect 152 738 174 746
rect 182 738 204 746
rect 212 738 234 746
rect 242 738 264 746
rect 272 738 286 746
rect 294 738 306 746
rect 314 738 328 746
rect 336 738 358 746
rect 366 738 388 746
rect 396 738 418 746
rect 426 738 448 746
rect 456 738 478 746
rect 486 738 508 746
rect 516 738 538 746
rect 546 738 568 746
rect 576 738 588 746
rect 596 738 600 746
rect 0 736 600 738
rect 0 728 14 736
rect 22 728 224 736
rect 232 728 244 736
rect 262 728 276 736
rect 284 728 296 736
rect 304 728 316 736
rect 324 728 338 736
rect 356 728 368 736
rect 376 728 578 736
rect 586 728 600 736
rect 0 726 600 728
rect 0 718 4 726
rect 12 718 24 726
rect 32 718 54 726
rect 62 718 84 726
rect 92 718 114 726
rect 122 718 144 726
rect 152 718 174 726
rect 182 718 204 726
rect 212 718 234 726
rect 242 718 264 726
rect 272 718 286 726
rect 294 718 306 726
rect 314 718 328 726
rect 336 718 358 726
rect 366 718 388 726
rect 396 718 418 726
rect 426 718 448 726
rect 456 718 478 726
rect 486 718 508 726
rect 516 718 538 726
rect 546 718 568 726
rect 576 718 588 726
rect 596 718 600 726
rect 0 716 600 718
rect 0 708 14 716
rect 22 708 44 716
rect 52 708 74 716
rect 82 708 104 716
rect 112 708 134 716
rect 142 708 164 716
rect 172 708 194 716
rect 202 708 224 716
rect 232 708 244 716
rect 262 708 276 716
rect 284 708 296 716
rect 304 708 316 716
rect 324 708 338 716
rect 356 708 368 716
rect 376 708 398 716
rect 406 708 428 716
rect 436 708 458 716
rect 466 708 488 716
rect 496 708 518 716
rect 526 708 548 716
rect 556 708 578 716
rect 586 708 600 716
rect 0 706 600 708
rect 0 698 4 706
rect 12 698 24 706
rect 32 698 54 706
rect 62 698 84 706
rect 92 698 114 706
rect 122 698 144 706
rect 152 698 174 706
rect 182 698 204 706
rect 212 698 234 706
rect 242 698 264 706
rect 272 698 286 706
rect 294 698 306 706
rect 314 698 328 706
rect 336 698 358 706
rect 366 698 388 706
rect 396 698 418 706
rect 426 698 448 706
rect 456 698 478 706
rect 486 698 508 706
rect 516 698 538 706
rect 546 698 568 706
rect 576 698 588 706
rect 596 698 600 706
rect 0 697 600 698
rect 0 696 296 697
rect 0 688 14 696
rect 22 688 44 696
rect 52 688 74 696
rect 82 688 104 696
rect 112 688 134 696
rect 142 688 164 696
rect 172 688 194 696
rect 202 688 224 696
rect 232 688 244 696
rect 262 688 274 696
rect 282 689 296 696
rect 304 696 600 697
rect 304 689 318 696
rect 282 688 318 689
rect 326 688 338 696
rect 356 688 368 696
rect 376 688 398 696
rect 406 688 428 696
rect 436 688 458 696
rect 466 688 488 696
rect 496 688 518 696
rect 526 688 548 696
rect 556 688 578 696
rect 586 688 600 696
rect 0 644 14 652
rect 22 644 44 652
rect 52 644 74 652
rect 82 644 104 652
rect 112 644 134 652
rect 142 644 164 652
rect 172 644 290 652
rect 298 644 302 652
rect 310 644 428 652
rect 436 644 458 652
rect 466 644 488 652
rect 496 644 518 652
rect 526 644 548 652
rect 556 644 578 652
rect 586 644 600 652
rect 0 642 600 644
rect 0 634 4 642
rect 12 634 24 642
rect 32 634 54 642
rect 62 634 84 642
rect 92 634 114 642
rect 122 634 144 642
rect 152 634 174 642
rect 182 634 418 642
rect 426 634 448 642
rect 456 634 478 642
rect 486 634 508 642
rect 516 634 538 642
rect 546 634 568 642
rect 576 634 588 642
rect 596 634 600 642
rect 0 632 600 634
rect 0 624 14 632
rect 22 624 44 632
rect 52 624 74 632
rect 82 624 104 632
rect 112 624 134 632
rect 142 624 164 632
rect 172 624 290 632
rect 298 624 302 632
rect 310 624 428 632
rect 436 624 458 632
rect 466 624 488 632
rect 496 624 518 632
rect 526 624 548 632
rect 556 624 578 632
rect 586 624 600 632
rect 0 622 600 624
rect 0 614 4 622
rect 12 614 24 622
rect 32 614 54 622
rect 62 614 84 622
rect 92 614 114 622
rect 122 614 144 622
rect 152 614 174 622
rect 182 614 418 622
rect 426 614 448 622
rect 456 614 478 622
rect 486 614 508 622
rect 516 614 538 622
rect 546 614 568 622
rect 576 614 588 622
rect 596 614 600 622
rect 0 612 600 614
rect 0 604 14 612
rect 22 604 290 612
rect 298 604 302 612
rect 310 604 578 612
rect 586 604 600 612
rect 0 602 600 604
rect 0 594 4 602
rect 12 594 24 602
rect 32 594 54 602
rect 62 594 84 602
rect 92 594 114 602
rect 122 594 144 602
rect 152 594 174 602
rect 182 594 418 602
rect 426 594 448 602
rect 456 594 478 602
rect 486 594 508 602
rect 516 594 538 602
rect 546 594 568 602
rect 576 594 588 602
rect 596 594 600 602
rect 0 592 290 594
rect 0 584 14 592
rect 22 584 44 592
rect 52 584 74 592
rect 82 584 104 592
rect 112 584 134 592
rect 142 584 164 592
rect 172 586 290 592
rect 298 586 302 594
rect 310 592 600 594
rect 310 586 428 592
rect 172 584 428 586
rect 436 584 458 592
rect 466 584 488 592
rect 496 584 518 592
rect 526 584 548 592
rect 556 584 578 592
rect 586 584 600 592
rect 0 582 600 584
rect 0 574 4 582
rect 12 574 24 582
rect 32 574 54 582
rect 62 574 84 582
rect 92 574 100 582
rect 0 572 100 574
rect 500 574 508 582
rect 516 574 538 582
rect 546 574 568 582
rect 576 574 588 582
rect 596 574 600 582
rect 500 572 600 574
rect 0 564 14 572
rect 22 564 44 572
rect 52 564 74 572
rect 82 564 104 572
rect 112 564 134 572
rect 142 564 164 572
rect 172 564 428 572
rect 436 564 458 572
rect 466 564 488 572
rect 496 564 518 572
rect 526 564 548 572
rect 556 564 578 572
rect 586 564 600 572
rect 0 562 290 564
rect 0 554 4 562
rect 12 554 24 562
rect 32 554 54 562
rect 62 554 84 562
rect 92 554 114 562
rect 122 554 144 562
rect 152 554 174 562
rect 182 556 290 562
rect 298 556 302 564
rect 310 562 600 564
rect 310 556 418 562
rect 182 554 418 556
rect 426 554 448 562
rect 456 554 478 562
rect 486 554 508 562
rect 516 554 538 562
rect 546 554 568 562
rect 576 554 588 562
rect 596 554 600 562
rect 0 552 600 554
rect 0 544 14 552
rect 22 544 44 552
rect 52 544 74 552
rect 82 544 104 552
rect 112 544 134 552
rect 142 544 164 552
rect 172 544 428 552
rect 436 544 458 552
rect 466 544 488 552
rect 496 544 518 552
rect 526 544 548 552
rect 556 544 578 552
rect 586 544 600 552
rect 0 542 290 544
rect 0 534 4 542
rect 12 534 24 542
rect 32 534 54 542
rect 62 534 84 542
rect 92 534 114 542
rect 122 534 144 542
rect 152 534 174 542
rect 182 536 290 542
rect 298 536 302 544
rect 310 542 600 544
rect 310 536 418 542
rect 182 534 418 536
rect 426 534 448 542
rect 456 534 478 542
rect 486 534 508 542
rect 516 534 538 542
rect 546 534 568 542
rect 576 534 588 542
rect 596 534 600 542
rect 0 532 600 534
rect 0 524 14 532
rect 22 524 44 532
rect 52 524 74 532
rect 82 524 104 532
rect 112 524 134 532
rect 142 524 164 532
rect 172 524 428 532
rect 436 524 458 532
rect 466 524 488 532
rect 496 524 518 532
rect 526 524 548 532
rect 556 524 578 532
rect 586 524 600 532
rect 0 516 290 524
rect 298 516 302 524
rect 310 516 600 524
rect 0 508 14 516
rect 22 508 34 516
rect 42 508 54 516
rect 62 508 74 516
rect 82 508 94 516
rect 102 508 114 516
rect 122 508 134 516
rect 142 508 154 516
rect 162 508 174 516
rect 182 508 418 516
rect 426 508 438 516
rect 446 508 458 516
rect 466 508 478 516
rect 486 508 498 516
rect 506 508 518 516
rect 526 508 538 516
rect 546 508 558 516
rect 566 508 578 516
rect 586 508 600 516
rect 0 492 600 508
rect 0 459 600 460
rect 0 451 30 459
rect 38 451 50 459
rect 58 451 80 459
rect 88 451 110 459
rect 118 451 140 459
rect 148 451 170 459
rect 178 451 200 459
rect 208 451 230 459
rect 238 451 260 459
rect 268 451 290 459
rect 298 451 320 459
rect 328 451 350 459
rect 358 451 380 459
rect 388 451 410 459
rect 418 451 440 459
rect 448 451 470 459
rect 478 451 500 459
rect 508 451 530 459
rect 538 451 560 459
rect 568 451 600 459
rect 0 449 600 451
rect 0 441 40 449
rect 48 441 70 449
rect 78 441 100 449
rect 108 441 130 449
rect 138 441 160 449
rect 168 441 190 449
rect 198 441 220 449
rect 228 441 250 449
rect 258 441 280 449
rect 288 441 310 449
rect 318 441 340 449
rect 348 441 370 449
rect 378 441 400 449
rect 408 441 430 449
rect 438 441 460 449
rect 468 441 490 449
rect 498 441 520 449
rect 528 441 550 449
rect 558 441 600 449
rect 0 439 600 441
rect 0 431 30 439
rect 38 431 50 439
rect 58 431 80 439
rect 88 431 110 439
rect 118 431 140 439
rect 148 431 170 439
rect 178 431 200 439
rect 208 431 230 439
rect 238 431 260 439
rect 268 431 290 439
rect 298 431 320 439
rect 328 431 350 439
rect 358 431 380 439
rect 388 431 410 439
rect 418 431 440 439
rect 448 431 470 439
rect 478 431 500 439
rect 508 431 530 439
rect 538 431 560 439
rect 568 431 600 439
rect 0 429 600 431
rect 0 421 40 429
rect 48 421 70 429
rect 78 421 100 429
rect 108 421 130 429
rect 138 421 160 429
rect 168 421 190 429
rect 198 421 220 429
rect 228 421 250 429
rect 258 421 280 429
rect 288 421 310 429
rect 318 421 340 429
rect 348 421 370 429
rect 378 421 400 429
rect 408 421 430 429
rect 438 421 460 429
rect 468 421 490 429
rect 498 421 520 429
rect 528 421 550 429
rect 558 421 600 429
rect 0 419 600 421
rect 0 411 30 419
rect 38 411 50 419
rect 58 411 80 419
rect 88 411 110 419
rect 118 411 140 419
rect 148 411 170 419
rect 178 411 200 419
rect 208 411 230 419
rect 238 411 260 419
rect 268 411 290 419
rect 298 411 320 419
rect 328 411 350 419
rect 358 411 380 419
rect 388 411 410 419
rect 418 411 440 419
rect 448 411 470 419
rect 478 411 500 419
rect 508 411 530 419
rect 538 411 560 419
rect 568 411 600 419
rect 0 409 600 411
rect 0 401 40 409
rect 48 401 70 409
rect 78 401 100 409
rect 108 401 130 409
rect 138 401 160 409
rect 168 401 190 409
rect 198 401 220 409
rect 228 401 250 409
rect 258 401 280 409
rect 288 401 310 409
rect 318 401 340 409
rect 348 401 370 409
rect 378 401 400 409
rect 408 401 430 409
rect 438 401 460 409
rect 468 401 490 409
rect 498 401 520 409
rect 528 401 550 409
rect 558 401 600 409
rect 0 399 600 401
rect 0 371 30 399
rect 38 371 50 399
rect 58 371 80 399
rect 88 391 110 399
rect 118 391 140 399
rect 148 391 170 399
rect 178 391 200 399
rect 208 391 230 399
rect 238 391 260 399
rect 268 391 290 399
rect 298 391 320 399
rect 328 391 350 399
rect 358 391 380 399
rect 388 391 410 399
rect 418 391 440 399
rect 448 391 470 399
rect 478 391 500 399
rect 88 379 500 391
rect 88 371 110 379
rect 118 371 140 379
rect 148 371 170 379
rect 178 371 200 379
rect 208 371 230 379
rect 238 371 260 379
rect 268 371 290 379
rect 298 371 320 379
rect 328 371 350 379
rect 358 371 380 379
rect 388 371 410 379
rect 418 371 440 379
rect 448 371 470 379
rect 478 371 500 379
rect 508 391 530 399
rect 538 391 560 399
rect 568 391 600 399
rect 508 389 600 391
rect 508 381 520 389
rect 528 381 550 389
rect 558 381 600 389
rect 508 379 600 381
rect 508 371 530 379
rect 538 371 560 379
rect 568 371 600 379
rect 0 369 600 371
rect 0 361 40 369
rect 48 361 70 369
rect 78 361 100 369
rect 108 361 130 369
rect 138 361 160 369
rect 168 361 190 369
rect 198 361 220 369
rect 228 361 250 369
rect 258 361 280 369
rect 288 361 310 369
rect 318 361 340 369
rect 348 361 370 369
rect 378 361 400 369
rect 408 361 430 369
rect 438 361 460 369
rect 468 361 490 369
rect 498 361 520 369
rect 528 361 550 369
rect 558 361 600 369
rect 0 359 600 361
rect 0 351 30 359
rect 38 351 50 359
rect 58 351 80 359
rect 88 351 110 359
rect 118 351 140 359
rect 148 351 170 359
rect 178 351 200 359
rect 208 351 230 359
rect 238 351 260 359
rect 268 351 290 359
rect 298 351 320 359
rect 328 351 350 359
rect 358 351 380 359
rect 388 351 410 359
rect 418 351 440 359
rect 448 351 470 359
rect 478 351 500 359
rect 508 351 530 359
rect 538 351 560 359
rect 568 351 600 359
rect 0 349 600 351
rect 0 341 40 349
rect 48 341 70 349
rect 78 341 100 349
rect 108 341 130 349
rect 138 341 160 349
rect 168 341 190 349
rect 198 341 220 349
rect 228 341 250 349
rect 258 341 280 349
rect 288 341 310 349
rect 318 341 340 349
rect 348 341 370 349
rect 378 341 400 349
rect 408 341 430 349
rect 438 341 460 349
rect 468 341 490 349
rect 498 341 520 349
rect 528 341 550 349
rect 558 341 600 349
rect 0 339 600 341
rect 0 331 30 339
rect 38 331 50 339
rect 58 331 80 339
rect 88 331 110 339
rect 118 331 140 339
rect 148 331 170 339
rect 178 331 200 339
rect 208 331 230 339
rect 238 331 260 339
rect 268 331 290 339
rect 298 331 320 339
rect 328 331 350 339
rect 358 331 380 339
rect 388 331 410 339
rect 418 331 440 339
rect 448 331 470 339
rect 478 331 500 339
rect 508 331 530 339
rect 538 331 560 339
rect 568 331 600 339
rect 0 329 600 331
rect 0 321 40 329
rect 48 321 70 329
rect 78 321 100 329
rect 108 321 130 329
rect 138 321 160 329
rect 168 321 190 329
rect 198 321 220 329
rect 228 321 250 329
rect 258 321 280 329
rect 288 321 310 329
rect 318 321 340 329
rect 348 321 370 329
rect 378 321 400 329
rect 408 321 430 329
rect 438 321 460 329
rect 468 321 490 329
rect 498 321 520 329
rect 528 321 550 329
rect 558 321 600 329
rect 0 319 600 321
rect 0 311 30 319
rect 38 311 50 319
rect 58 311 80 319
rect 88 311 110 319
rect 118 311 140 319
rect 148 311 170 319
rect 178 311 200 319
rect 208 311 230 319
rect 238 311 260 319
rect 268 311 290 319
rect 298 311 320 319
rect 328 311 350 319
rect 358 311 380 319
rect 388 311 410 319
rect 418 311 440 319
rect 448 311 470 319
rect 478 311 500 319
rect 508 311 530 319
rect 538 311 560 319
rect 568 311 600 319
rect 0 310 600 311
rect 0 309 100 310
rect 0 301 40 309
rect 48 301 70 309
rect 78 301 90 309
rect 98 301 100 309
rect 0 300 100 301
rect 500 309 600 310
rect 500 301 520 309
rect 528 301 550 309
rect 558 301 600 309
rect 500 300 600 301
rect 0 299 600 300
rect 0 291 30 299
rect 38 291 50 299
rect 58 291 80 299
rect 88 291 110 299
rect 118 291 140 299
rect 148 291 170 299
rect 178 291 200 299
rect 208 291 230 299
rect 238 291 260 299
rect 268 291 290 299
rect 298 291 320 299
rect 328 291 350 299
rect 358 291 380 299
rect 388 291 410 299
rect 418 291 440 299
rect 448 291 470 299
rect 478 291 500 299
rect 508 291 530 299
rect 538 291 560 299
rect 568 291 600 299
rect 0 289 600 291
rect 0 281 40 289
rect 48 281 70 289
rect 78 281 100 289
rect 108 281 130 289
rect 138 281 160 289
rect 168 281 190 289
rect 198 281 220 289
rect 228 281 250 289
rect 258 281 280 289
rect 288 281 310 289
rect 318 281 340 289
rect 348 281 370 289
rect 378 281 400 289
rect 408 281 430 289
rect 438 281 460 289
rect 468 281 490 289
rect 498 281 520 289
rect 528 281 550 289
rect 558 281 600 289
rect 0 279 600 281
rect 0 271 30 279
rect 38 271 50 279
rect 58 271 80 279
rect 88 271 110 279
rect 118 271 140 279
rect 148 271 170 279
rect 178 271 200 279
rect 208 271 230 279
rect 238 271 260 279
rect 268 271 290 279
rect 298 271 320 279
rect 328 271 350 279
rect 358 271 380 279
rect 388 271 410 279
rect 418 271 440 279
rect 448 271 470 279
rect 478 271 500 279
rect 508 271 530 279
rect 538 271 560 279
rect 568 271 600 279
rect 0 269 600 271
rect 0 261 40 269
rect 48 261 70 269
rect 78 261 100 269
rect 108 261 130 269
rect 138 261 160 269
rect 168 261 190 269
rect 198 261 220 269
rect 228 261 250 269
rect 258 261 280 269
rect 288 261 310 269
rect 318 261 340 269
rect 348 261 370 269
rect 378 261 400 269
rect 408 261 430 269
rect 438 261 460 269
rect 468 261 490 269
rect 498 261 520 269
rect 528 261 550 269
rect 558 261 600 269
rect 0 259 600 261
rect 0 251 30 259
rect 38 251 50 259
rect 58 251 80 259
rect 88 251 110 259
rect 118 251 140 259
rect 148 251 170 259
rect 178 251 200 259
rect 208 251 230 259
rect 238 251 260 259
rect 268 251 290 259
rect 298 251 320 259
rect 328 251 350 259
rect 358 251 380 259
rect 388 251 410 259
rect 418 251 440 259
rect 448 251 470 259
rect 478 251 500 259
rect 508 251 530 259
rect 538 251 560 259
rect 568 251 600 259
rect 0 249 600 251
rect 0 241 40 249
rect 48 241 70 249
rect 0 239 70 241
rect 0 231 30 239
rect 38 231 50 239
rect 58 231 70 239
rect 0 229 70 231
rect 0 221 40 229
rect 48 221 70 229
rect 78 241 100 249
rect 108 241 130 249
rect 138 241 160 249
rect 168 241 190 249
rect 198 241 220 249
rect 228 241 250 249
rect 258 241 280 249
rect 288 241 310 249
rect 318 241 340 249
rect 348 241 370 249
rect 378 241 400 249
rect 408 241 430 249
rect 438 241 460 249
rect 468 241 490 249
rect 498 241 520 249
rect 528 241 550 249
rect 558 241 600 249
rect 78 239 600 241
rect 78 231 510 239
rect 518 231 530 239
rect 538 231 560 239
rect 568 231 600 239
rect 78 229 600 231
rect 78 221 100 229
rect 108 221 130 229
rect 138 221 160 229
rect 168 221 190 229
rect 198 221 220 229
rect 228 221 250 229
rect 258 221 280 229
rect 288 221 310 229
rect 318 221 340 229
rect 348 221 370 229
rect 378 221 400 229
rect 408 221 430 229
rect 438 221 460 229
rect 468 221 490 229
rect 498 221 520 229
rect 528 221 550 229
rect 558 221 600 229
rect 0 219 600 221
rect 0 211 30 219
rect 38 211 50 219
rect 58 211 80 219
rect 88 211 110 219
rect 118 211 140 219
rect 148 211 170 219
rect 178 211 200 219
rect 208 211 230 219
rect 238 211 260 219
rect 268 211 290 219
rect 298 211 320 219
rect 328 211 350 219
rect 358 211 380 219
rect 388 211 410 219
rect 418 211 440 219
rect 448 211 470 219
rect 478 211 500 219
rect 508 211 530 219
rect 538 211 560 219
rect 568 211 600 219
rect 0 209 600 211
rect 0 201 40 209
rect 48 201 70 209
rect 78 201 100 209
rect 108 201 130 209
rect 138 201 160 209
rect 168 201 190 209
rect 198 201 220 209
rect 228 201 250 209
rect 258 201 280 209
rect 288 201 310 209
rect 318 201 340 209
rect 348 201 370 209
rect 378 201 400 209
rect 408 201 430 209
rect 438 201 460 209
rect 468 201 490 209
rect 498 201 520 209
rect 528 201 550 209
rect 558 201 600 209
rect 0 199 600 201
rect 0 191 30 199
rect 38 191 50 199
rect 58 191 80 199
rect 88 191 110 199
rect 118 191 140 199
rect 148 191 170 199
rect 178 191 200 199
rect 208 191 230 199
rect 238 191 260 199
rect 268 191 290 199
rect 298 191 320 199
rect 328 191 350 199
rect 358 191 380 199
rect 388 191 410 199
rect 418 191 440 199
rect 448 191 470 199
rect 478 191 500 199
rect 508 191 530 199
rect 538 191 560 199
rect 568 191 600 199
rect 0 189 600 191
rect 0 181 40 189
rect 48 181 70 189
rect 78 181 100 189
rect 108 181 130 189
rect 138 181 160 189
rect 168 181 190 189
rect 198 181 220 189
rect 228 181 250 189
rect 258 181 280 189
rect 288 181 310 189
rect 318 181 340 189
rect 348 181 370 189
rect 378 181 400 189
rect 408 181 430 189
rect 438 181 460 189
rect 468 181 490 189
rect 498 181 520 189
rect 528 181 550 189
rect 558 181 600 189
rect 0 179 600 181
rect 0 171 30 179
rect 38 171 50 179
rect 58 171 80 179
rect 88 171 110 179
rect 118 171 140 179
rect 148 171 170 179
rect 178 171 200 179
rect 208 171 230 179
rect 238 171 260 179
rect 268 171 290 179
rect 298 171 320 179
rect 328 171 350 179
rect 358 171 380 179
rect 388 171 410 179
rect 418 171 440 179
rect 448 171 470 179
rect 478 171 500 179
rect 508 171 530 179
rect 538 171 560 179
rect 568 171 600 179
rect 0 169 600 171
rect 0 161 40 169
rect 48 161 70 169
rect 78 161 100 169
rect 108 161 130 169
rect 138 161 160 169
rect 168 161 190 169
rect 198 161 220 169
rect 228 161 250 169
rect 258 161 280 169
rect 288 161 310 169
rect 318 161 340 169
rect 348 161 370 169
rect 378 161 400 169
rect 408 161 430 169
rect 438 161 460 169
rect 468 161 490 169
rect 498 161 520 169
rect 528 161 550 169
rect 558 161 600 169
rect 0 160 600 161
rect 0 159 100 160
rect 0 151 30 159
rect 38 151 50 159
rect 58 151 80 159
rect 88 151 100 159
rect 0 150 100 151
rect 500 159 600 160
rect 500 151 510 159
rect 518 151 530 159
rect 538 151 560 159
rect 568 151 600 159
rect 500 150 600 151
rect 0 149 600 150
rect 0 141 40 149
rect 48 141 70 149
rect 78 141 100 149
rect 108 141 130 149
rect 138 141 160 149
rect 168 141 190 149
rect 198 141 220 149
rect 228 141 250 149
rect 258 141 280 149
rect 288 141 310 149
rect 318 141 340 149
rect 348 141 370 149
rect 378 141 400 149
rect 408 141 430 149
rect 438 141 460 149
rect 468 141 490 149
rect 498 141 520 149
rect 528 141 550 149
rect 558 141 600 149
rect 0 139 600 141
rect 0 131 30 139
rect 38 131 50 139
rect 58 131 80 139
rect 88 131 110 139
rect 118 131 140 139
rect 148 131 170 139
rect 178 131 200 139
rect 208 131 230 139
rect 238 131 260 139
rect 268 131 290 139
rect 298 131 320 139
rect 328 131 350 139
rect 358 131 380 139
rect 388 131 410 139
rect 418 131 440 139
rect 448 131 470 139
rect 478 131 500 139
rect 508 131 530 139
rect 538 131 560 139
rect 568 131 600 139
rect 0 129 600 131
rect 0 121 40 129
rect 48 121 70 129
rect 78 121 100 129
rect 108 121 130 129
rect 138 121 160 129
rect 168 121 190 129
rect 198 121 220 129
rect 228 121 250 129
rect 258 121 280 129
rect 288 121 310 129
rect 318 121 340 129
rect 348 121 370 129
rect 378 121 400 129
rect 408 121 430 129
rect 438 121 460 129
rect 468 121 490 129
rect 498 121 520 129
rect 528 121 550 129
rect 558 121 600 129
rect 0 119 600 121
rect 0 111 30 119
rect 38 111 50 119
rect 58 111 80 119
rect 88 111 110 119
rect 118 111 140 119
rect 148 111 170 119
rect 178 111 200 119
rect 208 111 230 119
rect 238 111 260 119
rect 268 111 290 119
rect 298 111 320 119
rect 328 111 350 119
rect 358 111 380 119
rect 388 111 410 119
rect 418 111 440 119
rect 448 111 470 119
rect 478 111 500 119
rect 508 111 530 119
rect 538 111 560 119
rect 568 111 600 119
rect 0 109 600 111
rect 0 101 40 109
rect 48 101 70 109
rect 78 101 100 109
rect 108 101 130 109
rect 138 101 160 109
rect 168 101 190 109
rect 198 101 220 109
rect 228 101 250 109
rect 258 101 280 109
rect 288 101 310 109
rect 318 101 340 109
rect 348 101 370 109
rect 378 101 400 109
rect 408 101 430 109
rect 438 101 460 109
rect 468 101 490 109
rect 498 101 520 109
rect 528 101 550 109
rect 558 101 600 109
rect 0 99 600 101
rect 0 91 30 99
rect 38 91 50 99
rect 58 91 80 99
rect 88 91 110 99
rect 118 91 140 99
rect 148 91 170 99
rect 178 91 200 99
rect 208 91 230 99
rect 238 91 260 99
rect 268 91 290 99
rect 298 91 320 99
rect 328 91 350 99
rect 358 91 380 99
rect 388 91 410 99
rect 418 91 440 99
rect 448 91 470 99
rect 478 91 500 99
rect 508 91 530 99
rect 538 91 560 99
rect 568 91 600 99
rect 0 89 600 91
rect 0 81 40 89
rect 48 81 70 89
rect 78 81 100 89
rect 108 81 130 89
rect 138 81 160 89
rect 168 81 190 89
rect 198 81 220 89
rect 228 81 250 89
rect 258 81 280 89
rect 288 81 310 89
rect 318 81 340 89
rect 348 81 370 89
rect 378 81 400 89
rect 408 81 430 89
rect 438 81 460 89
rect 468 81 490 89
rect 498 81 520 89
rect 528 81 550 89
rect 558 81 600 89
rect 0 79 600 81
rect 0 71 30 79
rect 38 71 50 79
rect 58 71 80 79
rect 88 71 110 79
rect 118 71 140 79
rect 148 71 170 79
rect 178 71 200 79
rect 208 71 230 79
rect 238 71 260 79
rect 268 71 290 79
rect 298 71 320 79
rect 328 71 350 79
rect 358 71 380 79
rect 388 71 410 79
rect 418 71 440 79
rect 448 71 470 79
rect 478 71 500 79
rect 508 71 530 79
rect 538 71 560 79
rect 568 71 600 79
rect 0 69 600 71
rect 0 61 40 69
rect 48 61 70 69
rect 78 61 100 69
rect 108 61 130 69
rect 138 61 160 69
rect 168 61 190 69
rect 198 61 220 69
rect 228 61 250 69
rect 258 61 280 69
rect 288 61 310 69
rect 318 61 340 69
rect 348 61 370 69
rect 378 61 400 69
rect 408 61 430 69
rect 438 61 460 69
rect 468 61 490 69
rect 498 61 520 69
rect 528 61 550 69
rect 558 61 600 69
rect 0 59 600 61
rect 0 51 30 59
rect 38 51 50 59
rect 58 51 80 59
rect 88 51 110 59
rect 118 51 140 59
rect 148 51 170 59
rect 178 51 200 59
rect 208 51 230 59
rect 238 51 260 59
rect 268 51 290 59
rect 298 51 320 59
rect 328 51 350 59
rect 358 51 380 59
rect 388 51 410 59
rect 418 51 440 59
rect 448 51 470 59
rect 478 51 500 59
rect 508 51 530 59
rect 538 51 560 59
rect 568 51 600 59
rect 0 49 600 51
rect 0 41 40 49
rect 48 41 70 49
rect 78 41 100 49
rect 108 41 130 49
rect 138 41 160 49
rect 168 41 190 49
rect 198 41 220 49
rect 228 41 250 49
rect 258 41 280 49
rect 288 41 310 49
rect 318 41 340 49
rect 348 41 370 49
rect 378 41 400 49
rect 408 41 430 49
rect 438 41 460 49
rect 468 41 490 49
rect 498 41 520 49
rect 528 41 550 49
rect 558 41 600 49
rect 0 39 600 41
rect 0 31 30 39
rect 38 31 50 39
rect 58 31 80 39
rect 88 31 110 39
rect 118 31 140 39
rect 148 31 170 39
rect 178 31 200 39
rect 208 31 230 39
rect 238 31 260 39
rect 268 31 290 39
rect 298 31 320 39
rect 328 31 350 39
rect 358 31 380 39
rect 388 31 410 39
rect 418 31 440 39
rect 448 31 470 39
rect 478 31 500 39
rect 508 31 530 39
rect 538 31 560 39
rect 568 31 600 39
rect 0 12 600 31
rect 0 4 206 12
rect 394 4 600 12
rect 0 0 600 4
use PadBox  PadBox_0
timestamp 1570494029
transform 1 0 40 0 1 1480
box 0 0 520 520
<< labels >>
flabel nwell 600 -6 600 -6 6 FreeSans 16 0 0 0 VddNW
flabel nwell 0 -6 0 -6 4 FreeSans 16 0 0 0 VddNW
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 VddAct
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 VddAct
flabel psubstratepdiff 0 686 0 686 4 FreeSans 16 0 0 0 GndAct
flabel psubstratepdiff 600 686 600 686 6 FreeSans 16 0 0 0 GndAct
flabel metal1 204 0 204 0 4 FreeSans 64 0 0 0 GND
flabel metal2 0 0 0 0 4 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 0 600 0 6 FreeSans 16 0 0 0 GndM2A
flabel metal2 600 688 600 688 6 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 688 0 688 4 FreeSans 16 0 0 0 GndM2B
flabel metal2 0 880 0 880 4 FreeSans 16 0 0 0 VddM2A
flabel metal2 600 880 600 880 6 FreeSans 16 0 0 0 VddM2A
flabel metal2 0 492 0 492 4 FreeSans 16 0 0 0 VddM2B
flabel metal2 600 492 600 492 6 FreeSans 16 0 0 0 VddM2B
<< properties >>
string path 603.000 0.000 747.000 0.000 747.000 54.000 603.000 54.000 603.000 0.000 
<< end >>
